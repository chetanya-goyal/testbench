* NGSPICE file created from diffpair634.ext - technology: sky130A

.subckt diffpair634 minus drain_right drain_left source plus
X0 drain_left.t9 plus.t0 source.t8 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X1 a_n2072_n4888# a_n2072_n4888# a_n2072_n4888# a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.8
X2 drain_right.t9 minus.t0 source.t19 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X3 drain_right.t8 minus.t1 source.t4 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X4 a_n2072_n4888# a_n2072_n4888# a_n2072_n4888# a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X5 a_n2072_n4888# a_n2072_n4888# a_n2072_n4888# a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X6 source.t5 minus.t2 drain_right.t7 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X7 source.t11 plus.t1 drain_left.t8 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X8 drain_right.t6 minus.t3 source.t6 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X9 a_n2072_n4888# a_n2072_n4888# a_n2072_n4888# a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X10 source.t7 minus.t4 drain_right.t5 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X11 source.t10 plus.t2 drain_left.t7 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X12 drain_right.t4 minus.t5 source.t18 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X13 source.t1 minus.t6 drain_right.t3 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X14 source.t0 minus.t7 drain_right.t2 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X15 drain_right.t1 minus.t8 source.t2 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X16 source.t15 plus.t3 drain_left.t6 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X17 drain_left.t5 plus.t4 source.t9 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X18 drain_left.t4 plus.t5 source.t14 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X19 drain_left.t3 plus.t6 source.t12 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X20 drain_left.t2 plus.t7 source.t13 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X21 source.t17 plus.t8 drain_left.t1 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X22 drain_right.t0 minus.t9 source.t3 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X23 drain_left.t0 plus.t9 source.t16 a_n2072_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
R0 plus.n3 plus.t9 674.801
R1 plus.n13 plus.t0 674.801
R2 plus.n8 plus.t7 651.605
R3 plus.n6 plus.t3 651.605
R4 plus.n5 plus.t4 651.605
R5 plus.n4 plus.t8 651.605
R6 plus.n18 plus.t5 651.605
R7 plus.n16 plus.t1 651.605
R8 plus.n15 plus.t6 651.605
R9 plus.n14 plus.t2 651.605
R10 plus.n7 plus.n0 161.3
R11 plus.n9 plus.n8 161.3
R12 plus.n17 plus.n10 161.3
R13 plus.n19 plus.n18 161.3
R14 plus.n5 plus.n2 80.6037
R15 plus.n6 plus.n1 80.6037
R16 plus.n15 plus.n12 80.6037
R17 plus.n16 plus.n11 80.6037
R18 plus.n6 plus.n5 48.2005
R19 plus.n5 plus.n4 48.2005
R20 plus.n16 plus.n15 48.2005
R21 plus.n15 plus.n14 48.2005
R22 plus plus.n19 34.0577
R23 plus.n7 plus.n6 32.1338
R24 plus.n17 plus.n16 32.1338
R25 plus.n3 plus.n2 31.8629
R26 plus.n13 plus.n12 31.8629
R27 plus.n4 plus.n3 16.2333
R28 plus.n14 plus.n13 16.2333
R29 plus.n8 plus.n7 16.0672
R30 plus.n18 plus.n17 16.0672
R31 plus plus.n9 15.3509
R32 plus.n2 plus.n1 0.380177
R33 plus.n12 plus.n11 0.380177
R34 plus.n1 plus.n0 0.285035
R35 plus.n11 plus.n10 0.285035
R36 plus.n9 plus.n0 0.189894
R37 plus.n19 plus.n10 0.189894
R38 source.n0 source.t13 44.1297
R39 source.n5 source.t18 44.1296
R40 source.n19 source.t19 44.1295
R41 source.n14 source.t8 44.1295
R42 source.n2 source.n1 43.1397
R43 source.n4 source.n3 43.1397
R44 source.n7 source.n6 43.1397
R45 source.n9 source.n8 43.1397
R46 source.n18 source.n17 43.1396
R47 source.n16 source.n15 43.1396
R48 source.n13 source.n12 43.1396
R49 source.n11 source.n10 43.1396
R50 source.n11 source.n9 29.2966
R51 source.n20 source.n0 22.5725
R52 source.n20 source.n19 5.7505
R53 source.n17 source.t3 0.9905
R54 source.n17 source.t5 0.9905
R55 source.n15 source.t4 0.9905
R56 source.n15 source.t1 0.9905
R57 source.n12 source.t12 0.9905
R58 source.n12 source.t10 0.9905
R59 source.n10 source.t14 0.9905
R60 source.n10 source.t11 0.9905
R61 source.n1 source.t9 0.9905
R62 source.n1 source.t15 0.9905
R63 source.n3 source.t16 0.9905
R64 source.n3 source.t17 0.9905
R65 source.n6 source.t6 0.9905
R66 source.n6 source.t7 0.9905
R67 source.n8 source.t2 0.9905
R68 source.n8 source.t0 0.9905
R69 source.n9 source.n7 0.974638
R70 source.n7 source.n5 0.974638
R71 source.n4 source.n2 0.974638
R72 source.n2 source.n0 0.974638
R73 source.n13 source.n11 0.974638
R74 source.n14 source.n13 0.974638
R75 source.n18 source.n16 0.974638
R76 source.n19 source.n18 0.974638
R77 source.n5 source.n4 0.957397
R78 source.n16 source.n14 0.957397
R79 source source.n20 0.188
R80 drain_left.n5 drain_left.t0 61.7825
R81 drain_left.n1 drain_left.t4 61.7824
R82 drain_left.n3 drain_left.n2 60.4937
R83 drain_left.n7 drain_left.n6 59.8185
R84 drain_left.n5 drain_left.n4 59.8185
R85 drain_left.n1 drain_left.n0 59.8184
R86 drain_left drain_left.n3 37.5678
R87 drain_left drain_left.n7 6.62735
R88 drain_left.n2 drain_left.t7 0.9905
R89 drain_left.n2 drain_left.t9 0.9905
R90 drain_left.n0 drain_left.t8 0.9905
R91 drain_left.n0 drain_left.t3 0.9905
R92 drain_left.n6 drain_left.t6 0.9905
R93 drain_left.n6 drain_left.t2 0.9905
R94 drain_left.n4 drain_left.t1 0.9905
R95 drain_left.n4 drain_left.t5 0.9905
R96 drain_left.n7 drain_left.n5 0.974638
R97 drain_left.n3 drain_left.n1 0.188688
R98 minus.n3 minus.t5 674.801
R99 minus.n13 minus.t1 674.801
R100 minus.n2 minus.t4 651.605
R101 minus.n1 minus.t3 651.605
R102 minus.n6 minus.t7 651.605
R103 minus.n8 minus.t8 651.605
R104 minus.n12 minus.t6 651.605
R105 minus.n11 minus.t9 651.605
R106 minus.n16 minus.t2 651.605
R107 minus.n18 minus.t0 651.605
R108 minus.n9 minus.n8 161.3
R109 minus.n7 minus.n0 161.3
R110 minus.n19 minus.n18 161.3
R111 minus.n17 minus.n10 161.3
R112 minus.n6 minus.n5 80.6037
R113 minus.n4 minus.n1 80.6037
R114 minus.n16 minus.n15 80.6037
R115 minus.n14 minus.n11 80.6037
R116 minus.n2 minus.n1 48.2005
R117 minus.n6 minus.n1 48.2005
R118 minus.n12 minus.n11 48.2005
R119 minus.n16 minus.n11 48.2005
R120 minus.n20 minus.n9 43.2069
R121 minus.n7 minus.n6 32.1338
R122 minus.n17 minus.n16 32.1338
R123 minus.n4 minus.n3 31.8629
R124 minus.n14 minus.n13 31.8629
R125 minus.n3 minus.n2 16.2333
R126 minus.n13 minus.n12 16.2333
R127 minus.n8 minus.n7 16.0672
R128 minus.n18 minus.n17 16.0672
R129 minus.n20 minus.n19 6.67664
R130 minus.n5 minus.n4 0.380177
R131 minus.n15 minus.n14 0.380177
R132 minus.n5 minus.n0 0.285035
R133 minus.n15 minus.n10 0.285035
R134 minus.n9 minus.n0 0.189894
R135 minus.n19 minus.n10 0.189894
R136 minus minus.n20 0.188
R137 drain_right.n1 drain_right.t8 61.7824
R138 drain_right.n7 drain_right.t1 60.8084
R139 drain_right.n6 drain_right.n4 60.7926
R140 drain_right.n3 drain_right.n2 60.4937
R141 drain_right.n6 drain_right.n5 59.8185
R142 drain_right.n1 drain_right.n0 59.8184
R143 drain_right drain_right.n3 37.0145
R144 drain_right drain_right.n7 6.14028
R145 drain_right.n2 drain_right.t7 0.9905
R146 drain_right.n2 drain_right.t9 0.9905
R147 drain_right.n0 drain_right.t3 0.9905
R148 drain_right.n0 drain_right.t0 0.9905
R149 drain_right.n4 drain_right.t5 0.9905
R150 drain_right.n4 drain_right.t4 0.9905
R151 drain_right.n5 drain_right.t2 0.9905
R152 drain_right.n5 drain_right.t6 0.9905
R153 drain_right.n7 drain_right.n6 0.974638
R154 drain_right.n3 drain_right.n1 0.188688
C0 drain_right source 20.8318f
C1 drain_left plus 11.870599f
C2 drain_right plus 0.36134f
C3 drain_left drain_right 1.03631f
C4 minus source 11.2391f
C5 plus minus 7.205891f
C6 plus source 11.253901f
C7 drain_left minus 0.172418f
C8 drain_right minus 11.6715f
C9 drain_left source 20.8422f
C10 drain_right a_n2072_n4888# 9.211081f
C11 drain_left a_n2072_n4888# 9.521801f
C12 source a_n2072_n4888# 9.589526f
C13 minus a_n2072_n4888# 8.655111f
C14 plus a_n2072_n4888# 10.68226f
C15 drain_right.t8 a_n2072_n4888# 4.39301f
C16 drain_right.t3 a_n2072_n4888# 0.375239f
C17 drain_right.t0 a_n2072_n4888# 0.375239f
C18 drain_right.n0 a_n2072_n4888# 3.43051f
C19 drain_right.n1 a_n2072_n4888# 0.637524f
C20 drain_right.t7 a_n2072_n4888# 0.375239f
C21 drain_right.t9 a_n2072_n4888# 0.375239f
C22 drain_right.n2 a_n2072_n4888# 3.43427f
C23 drain_right.n3 a_n2072_n4888# 1.99504f
C24 drain_right.t5 a_n2072_n4888# 0.375239f
C25 drain_right.t4 a_n2072_n4888# 0.375239f
C26 drain_right.n4 a_n2072_n4888# 3.43626f
C27 drain_right.t2 a_n2072_n4888# 0.375239f
C28 drain_right.t6 a_n2072_n4888# 0.375239f
C29 drain_right.n5 a_n2072_n4888# 3.43051f
C30 drain_right.n6 a_n2072_n4888# 0.702622f
C31 drain_right.t1 a_n2072_n4888# 4.38749f
C32 drain_right.n7 a_n2072_n4888# 0.574019f
C33 minus.n0 a_n2072_n4888# 0.053505f
C34 minus.t3 a_n2072_n4888# 1.81683f
C35 minus.n1 a_n2072_n4888# 0.686136f
C36 minus.t7 a_n2072_n4888# 1.81683f
C37 minus.t5 a_n2072_n4888# 1.84009f
C38 minus.t4 a_n2072_n4888# 1.81683f
C39 minus.n2 a_n2072_n4888# 0.685166f
C40 minus.n3 a_n2072_n4888# 0.658113f
C41 minus.n4 a_n2072_n4888# 0.246065f
C42 minus.n5 a_n2072_n4888# 0.066787f
C43 minus.n6 a_n2072_n4888# 0.683417f
C44 minus.n7 a_n2072_n4888# 0.009099f
C45 minus.t8 a_n2072_n4888# 1.81683f
C46 minus.n8 a_n2072_n4888# 0.671598f
C47 minus.n9 a_n2072_n4888# 1.85559f
C48 minus.n10 a_n2072_n4888# 0.053505f
C49 minus.t9 a_n2072_n4888# 1.81683f
C50 minus.n11 a_n2072_n4888# 0.686136f
C51 minus.t1 a_n2072_n4888# 1.84009f
C52 minus.t6 a_n2072_n4888# 1.81683f
C53 minus.n12 a_n2072_n4888# 0.685166f
C54 minus.n13 a_n2072_n4888# 0.658113f
C55 minus.n14 a_n2072_n4888# 0.246065f
C56 minus.n15 a_n2072_n4888# 0.066787f
C57 minus.t2 a_n2072_n4888# 1.81683f
C58 minus.n16 a_n2072_n4888# 0.683417f
C59 minus.n17 a_n2072_n4888# 0.009099f
C60 minus.t0 a_n2072_n4888# 1.81683f
C61 minus.n18 a_n2072_n4888# 0.671598f
C62 minus.n19 a_n2072_n4888# 0.278696f
C63 minus.n20 a_n2072_n4888# 2.20479f
C64 drain_left.t4 a_n2072_n4888# 4.40744f
C65 drain_left.t8 a_n2072_n4888# 0.376472f
C66 drain_left.t3 a_n2072_n4888# 0.376472f
C67 drain_left.n0 a_n2072_n4888# 3.44179f
C68 drain_left.n1 a_n2072_n4888# 0.639619f
C69 drain_left.t7 a_n2072_n4888# 0.376472f
C70 drain_left.t9 a_n2072_n4888# 0.376472f
C71 drain_left.n2 a_n2072_n4888# 3.44556f
C72 drain_left.n3 a_n2072_n4888# 2.05103f
C73 drain_left.t0 a_n2072_n4888# 4.40746f
C74 drain_left.t1 a_n2072_n4888# 0.376472f
C75 drain_left.t5 a_n2072_n4888# 0.376472f
C76 drain_left.n4 a_n2072_n4888# 3.44178f
C77 drain_left.n5 a_n2072_n4888# 0.696998f
C78 drain_left.t6 a_n2072_n4888# 0.376472f
C79 drain_left.t2 a_n2072_n4888# 0.376472f
C80 drain_left.n6 a_n2072_n4888# 3.44178f
C81 drain_left.n7 a_n2072_n4888# 0.56415f
C82 source.t13 a_n2072_n4888# 4.3924f
C83 source.n0 a_n2072_n4888# 1.92146f
C84 source.t9 a_n2072_n4888# 0.384341f
C85 source.t15 a_n2072_n4888# 0.384341f
C86 source.n1 a_n2072_n4888# 3.43618f
C87 source.n2 a_n2072_n4888# 0.402381f
C88 source.t16 a_n2072_n4888# 0.384341f
C89 source.t17 a_n2072_n4888# 0.384341f
C90 source.n3 a_n2072_n4888# 3.43618f
C91 source.n4 a_n2072_n4888# 0.40103f
C92 source.t18 a_n2072_n4888# 4.39241f
C93 source.n5 a_n2072_n4888# 0.493001f
C94 source.t6 a_n2072_n4888# 0.384341f
C95 source.t7 a_n2072_n4888# 0.384341f
C96 source.n6 a_n2072_n4888# 3.43618f
C97 source.n7 a_n2072_n4888# 0.402381f
C98 source.t2 a_n2072_n4888# 0.384341f
C99 source.t0 a_n2072_n4888# 0.384341f
C100 source.n8 a_n2072_n4888# 3.43618f
C101 source.n9 a_n2072_n4888# 2.3511f
C102 source.t14 a_n2072_n4888# 0.384341f
C103 source.t11 a_n2072_n4888# 0.384341f
C104 source.n10 a_n2072_n4888# 3.43618f
C105 source.n11 a_n2072_n4888# 2.35109f
C106 source.t12 a_n2072_n4888# 0.384341f
C107 source.t10 a_n2072_n4888# 0.384341f
C108 source.n12 a_n2072_n4888# 3.43618f
C109 source.n13 a_n2072_n4888# 0.402374f
C110 source.t8 a_n2072_n4888# 4.39239f
C111 source.n14 a_n2072_n4888# 0.493025f
C112 source.t4 a_n2072_n4888# 0.384341f
C113 source.t1 a_n2072_n4888# 0.384341f
C114 source.n15 a_n2072_n4888# 3.43618f
C115 source.n16 a_n2072_n4888# 0.401023f
C116 source.t3 a_n2072_n4888# 0.384341f
C117 source.t5 a_n2072_n4888# 0.384341f
C118 source.n17 a_n2072_n4888# 3.43618f
C119 source.n18 a_n2072_n4888# 0.402374f
C120 source.t19 a_n2072_n4888# 4.39239f
C121 source.n19 a_n2072_n4888# 0.618753f
C122 source.n20 a_n2072_n4888# 2.21059f
C123 plus.n0 a_n2072_n4888# 0.054184f
C124 plus.t7 a_n2072_n4888# 1.83989f
C125 plus.t3 a_n2072_n4888# 1.83989f
C126 plus.n1 a_n2072_n4888# 0.067635f
C127 plus.t4 a_n2072_n4888# 1.83989f
C128 plus.n2 a_n2072_n4888# 0.249189f
C129 plus.t8 a_n2072_n4888# 1.83989f
C130 plus.t9 a_n2072_n4888# 1.86345f
C131 plus.n3 a_n2072_n4888# 0.666468f
C132 plus.n4 a_n2072_n4888# 0.693864f
C133 plus.n5 a_n2072_n4888# 0.694847f
C134 plus.n6 a_n2072_n4888# 0.692093f
C135 plus.n7 a_n2072_n4888# 0.009214f
C136 plus.n8 a_n2072_n4888# 0.680124f
C137 plus.n9 a_n2072_n4888# 0.633025f
C138 plus.n10 a_n2072_n4888# 0.054184f
C139 plus.t5 a_n2072_n4888# 1.83989f
C140 plus.n11 a_n2072_n4888# 0.067635f
C141 plus.t1 a_n2072_n4888# 1.83989f
C142 plus.n12 a_n2072_n4888# 0.249189f
C143 plus.t6 a_n2072_n4888# 1.83989f
C144 plus.t0 a_n2072_n4888# 1.86345f
C145 plus.n13 a_n2072_n4888# 0.666468f
C146 plus.t2 a_n2072_n4888# 1.83989f
C147 plus.n14 a_n2072_n4888# 0.693864f
C148 plus.n15 a_n2072_n4888# 0.694847f
C149 plus.n16 a_n2072_n4888# 0.692093f
C150 plus.n17 a_n2072_n4888# 0.009214f
C151 plus.n18 a_n2072_n4888# 0.680124f
C152 plus.n19 a_n2072_n4888# 1.49447f
.ends

