* NGSPICE file created from diffpair387.ext - technology: sky130A

.subckt diffpair387 minus drain_right drain_left source plus
X0 source.t31 plus.t0 drain_left.t14 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X1 source.t30 plus.t1 drain_left.t13 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X2 source.t8 minus.t0 drain_right.t15 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X3 source.t29 plus.t2 drain_left.t1 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X4 source.t28 plus.t3 drain_left.t15 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X5 a_n2570_n2688# a_n2570_n2688# a_n2570_n2688# a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.7
X6 a_n2570_n2688# a_n2570_n2688# a_n2570_n2688# a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X7 source.t27 plus.t4 drain_left.t3 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X8 drain_left.t4 plus.t5 source.t26 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X9 drain_right.t14 minus.t1 source.t12 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X10 drain_right.t13 minus.t2 source.t6 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X11 drain_right.t12 minus.t3 source.t7 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X12 drain_left.t6 plus.t6 source.t25 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X13 drain_left.t2 plus.t7 source.t24 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X14 drain_right.t11 minus.t4 source.t11 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X15 drain_left.t7 plus.t8 source.t23 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X16 drain_left.t9 plus.t9 source.t22 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X17 drain_right.t10 minus.t5 source.t0 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X18 drain_right.t9 minus.t6 source.t10 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X19 source.t14 minus.t7 drain_right.t8 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X20 drain_left.t11 plus.t10 source.t21 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X21 source.t20 plus.t11 drain_left.t0 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X22 drain_left.t10 plus.t12 source.t19 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X23 source.t1 minus.t8 drain_right.t7 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X24 source.t18 plus.t13 drain_left.t5 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X25 drain_right.t6 minus.t9 source.t2 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X26 source.t3 minus.t10 drain_right.t5 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X27 a_n2570_n2688# a_n2570_n2688# a_n2570_n2688# a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X28 source.t9 minus.t11 drain_right.t4 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X29 a_n2570_n2688# a_n2570_n2688# a_n2570_n2688# a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X30 source.t17 plus.t14 drain_left.t12 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X31 drain_left.t8 plus.t15 source.t16 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X32 source.t13 minus.t12 drain_right.t3 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X33 source.t4 minus.t13 drain_right.t2 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X34 drain_right.t1 minus.t14 source.t5 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X35 source.t15 minus.t15 drain_right.t0 a_n2570_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
R0 plus.n7 plus.t3 390.351
R1 plus.n33 plus.t12 390.351
R2 plus.n24 plus.t6 365.976
R3 plus.n22 plus.t0 365.976
R4 plus.n2 plus.t9 365.976
R5 plus.n16 plus.t2 365.976
R6 plus.n4 plus.t8 365.976
R7 plus.n10 plus.t1 365.976
R8 plus.n6 plus.t10 365.976
R9 plus.n50 plus.t11 365.976
R10 plus.n48 plus.t15 365.976
R11 plus.n28 plus.t14 365.976
R12 plus.n42 plus.t5 365.976
R13 plus.n30 plus.t4 365.976
R14 plus.n36 plus.t7 365.976
R15 plus.n32 plus.t13 365.976
R16 plus.n9 plus.n8 161.3
R17 plus.n10 plus.n5 161.3
R18 plus.n12 plus.n11 161.3
R19 plus.n13 plus.n4 161.3
R20 plus.n15 plus.n14 161.3
R21 plus.n16 plus.n3 161.3
R22 plus.n18 plus.n17 161.3
R23 plus.n19 plus.n2 161.3
R24 plus.n21 plus.n20 161.3
R25 plus.n22 plus.n1 161.3
R26 plus.n23 plus.n0 161.3
R27 plus.n25 plus.n24 161.3
R28 plus.n35 plus.n34 161.3
R29 plus.n36 plus.n31 161.3
R30 plus.n38 plus.n37 161.3
R31 plus.n39 plus.n30 161.3
R32 plus.n41 plus.n40 161.3
R33 plus.n42 plus.n29 161.3
R34 plus.n44 plus.n43 161.3
R35 plus.n45 plus.n28 161.3
R36 plus.n47 plus.n46 161.3
R37 plus.n48 plus.n27 161.3
R38 plus.n49 plus.n26 161.3
R39 plus.n51 plus.n50 161.3
R40 plus.n8 plus.n7 44.9377
R41 plus.n34 plus.n33 44.9377
R42 plus.n24 plus.n23 37.246
R43 plus.n50 plus.n49 37.246
R44 plus.n22 plus.n21 32.8641
R45 plus.n9 plus.n6 32.8641
R46 plus.n48 plus.n47 32.8641
R47 plus.n35 plus.n32 32.8641
R48 plus plus.n51 31.7566
R49 plus.n17 plus.n2 28.4823
R50 plus.n11 plus.n10 28.4823
R51 plus.n43 plus.n28 28.4823
R52 plus.n37 plus.n36 28.4823
R53 plus.n15 plus.n4 24.1005
R54 plus.n16 plus.n15 24.1005
R55 plus.n42 plus.n41 24.1005
R56 plus.n41 plus.n30 24.1005
R57 plus.n17 plus.n16 19.7187
R58 plus.n11 plus.n4 19.7187
R59 plus.n43 plus.n42 19.7187
R60 plus.n37 plus.n30 19.7187
R61 plus.n7 plus.n6 17.0522
R62 plus.n33 plus.n32 17.0522
R63 plus.n21 plus.n2 15.3369
R64 plus.n10 plus.n9 15.3369
R65 plus.n47 plus.n28 15.3369
R66 plus.n36 plus.n35 15.3369
R67 plus plus.n25 11.1634
R68 plus.n23 plus.n22 10.955
R69 plus.n49 plus.n48 10.955
R70 plus.n8 plus.n5 0.189894
R71 plus.n12 plus.n5 0.189894
R72 plus.n13 plus.n12 0.189894
R73 plus.n14 plus.n13 0.189894
R74 plus.n14 plus.n3 0.189894
R75 plus.n18 plus.n3 0.189894
R76 plus.n19 plus.n18 0.189894
R77 plus.n20 plus.n19 0.189894
R78 plus.n20 plus.n1 0.189894
R79 plus.n1 plus.n0 0.189894
R80 plus.n25 plus.n0 0.189894
R81 plus.n51 plus.n26 0.189894
R82 plus.n27 plus.n26 0.189894
R83 plus.n46 plus.n27 0.189894
R84 plus.n46 plus.n45 0.189894
R85 plus.n45 plus.n44 0.189894
R86 plus.n44 plus.n29 0.189894
R87 plus.n40 plus.n29 0.189894
R88 plus.n40 plus.n39 0.189894
R89 plus.n39 plus.n38 0.189894
R90 plus.n38 plus.n31 0.189894
R91 plus.n34 plus.n31 0.189894
R92 drain_left.n9 drain_left.n7 66.4255
R93 drain_left.n5 drain_left.n3 66.4253
R94 drain_left.n2 drain_left.n0 66.4253
R95 drain_left.n11 drain_left.n10 65.5376
R96 drain_left.n9 drain_left.n8 65.5376
R97 drain_left.n13 drain_left.n12 65.5374
R98 drain_left.n5 drain_left.n4 65.5373
R99 drain_left.n2 drain_left.n1 65.5373
R100 drain_left drain_left.n6 30.8659
R101 drain_left drain_left.n13 6.54115
R102 drain_left.n3 drain_left.t5 2.2005
R103 drain_left.n3 drain_left.t10 2.2005
R104 drain_left.n4 drain_left.t3 2.2005
R105 drain_left.n4 drain_left.t2 2.2005
R106 drain_left.n1 drain_left.t12 2.2005
R107 drain_left.n1 drain_left.t4 2.2005
R108 drain_left.n0 drain_left.t0 2.2005
R109 drain_left.n0 drain_left.t8 2.2005
R110 drain_left.n12 drain_left.t14 2.2005
R111 drain_left.n12 drain_left.t6 2.2005
R112 drain_left.n10 drain_left.t1 2.2005
R113 drain_left.n10 drain_left.t9 2.2005
R114 drain_left.n8 drain_left.t13 2.2005
R115 drain_left.n8 drain_left.t7 2.2005
R116 drain_left.n7 drain_left.t15 2.2005
R117 drain_left.n7 drain_left.t11 2.2005
R118 drain_left.n11 drain_left.n9 0.888431
R119 drain_left.n13 drain_left.n11 0.888431
R120 drain_left.n6 drain_left.n5 0.389119
R121 drain_left.n6 drain_left.n2 0.389119
R122 source.n7 source.t28 51.0588
R123 source.n8 source.t10 51.0588
R124 source.n15 source.t3 51.0588
R125 source.n31 source.t6 51.0586
R126 source.n24 source.t15 51.0586
R127 source.n23 source.t19 51.0586
R128 source.n16 source.t20 51.0586
R129 source.n0 source.t25 51.0586
R130 source.n2 source.n1 48.8588
R131 source.n4 source.n3 48.8588
R132 source.n6 source.n5 48.8588
R133 source.n10 source.n9 48.8588
R134 source.n12 source.n11 48.8588
R135 source.n14 source.n13 48.8588
R136 source.n30 source.n29 48.8586
R137 source.n28 source.n27 48.8586
R138 source.n26 source.n25 48.8586
R139 source.n22 source.n21 48.8586
R140 source.n20 source.n19 48.8586
R141 source.n18 source.n17 48.8586
R142 source.n16 source.n15 19.9029
R143 source.n32 source.n0 14.196
R144 source.n32 source.n31 5.7074
R145 source.n29 source.t0 2.2005
R146 source.n29 source.t14 2.2005
R147 source.n27 source.t2 2.2005
R148 source.n27 source.t9 2.2005
R149 source.n25 source.t5 2.2005
R150 source.n25 source.t1 2.2005
R151 source.n21 source.t24 2.2005
R152 source.n21 source.t18 2.2005
R153 source.n19 source.t26 2.2005
R154 source.n19 source.t27 2.2005
R155 source.n17 source.t16 2.2005
R156 source.n17 source.t17 2.2005
R157 source.n1 source.t22 2.2005
R158 source.n1 source.t31 2.2005
R159 source.n3 source.t23 2.2005
R160 source.n3 source.t29 2.2005
R161 source.n5 source.t21 2.2005
R162 source.n5 source.t30 2.2005
R163 source.n9 source.t11 2.2005
R164 source.n9 source.t8 2.2005
R165 source.n11 source.t7 2.2005
R166 source.n11 source.t13 2.2005
R167 source.n13 source.t12 2.2005
R168 source.n13 source.t4 2.2005
R169 source.n15 source.n14 0.888431
R170 source.n14 source.n12 0.888431
R171 source.n12 source.n10 0.888431
R172 source.n10 source.n8 0.888431
R173 source.n7 source.n6 0.888431
R174 source.n6 source.n4 0.888431
R175 source.n4 source.n2 0.888431
R176 source.n2 source.n0 0.888431
R177 source.n18 source.n16 0.888431
R178 source.n20 source.n18 0.888431
R179 source.n22 source.n20 0.888431
R180 source.n23 source.n22 0.888431
R181 source.n26 source.n24 0.888431
R182 source.n28 source.n26 0.888431
R183 source.n30 source.n28 0.888431
R184 source.n31 source.n30 0.888431
R185 source.n8 source.n7 0.470328
R186 source.n24 source.n23 0.470328
R187 source source.n32 0.188
R188 minus.n7 minus.t6 390.351
R189 minus.n33 minus.t15 390.351
R190 minus.n6 minus.t0 365.976
R191 minus.n10 minus.t4 365.976
R192 minus.n12 minus.t12 365.976
R193 minus.n16 minus.t3 365.976
R194 minus.n18 minus.t13 365.976
R195 minus.n22 minus.t1 365.976
R196 minus.n24 minus.t10 365.976
R197 minus.n32 minus.t14 365.976
R198 minus.n36 minus.t8 365.976
R199 minus.n38 minus.t9 365.976
R200 minus.n42 minus.t11 365.976
R201 minus.n44 minus.t5 365.976
R202 minus.n48 minus.t7 365.976
R203 minus.n50 minus.t2 365.976
R204 minus.n25 minus.n24 161.3
R205 minus.n23 minus.n0 161.3
R206 minus.n22 minus.n21 161.3
R207 minus.n20 minus.n1 161.3
R208 minus.n19 minus.n18 161.3
R209 minus.n17 minus.n2 161.3
R210 minus.n16 minus.n15 161.3
R211 minus.n14 minus.n3 161.3
R212 minus.n13 minus.n12 161.3
R213 minus.n11 minus.n4 161.3
R214 minus.n10 minus.n9 161.3
R215 minus.n8 minus.n5 161.3
R216 minus.n51 minus.n50 161.3
R217 minus.n49 minus.n26 161.3
R218 minus.n48 minus.n47 161.3
R219 minus.n46 minus.n27 161.3
R220 minus.n45 minus.n44 161.3
R221 minus.n43 minus.n28 161.3
R222 minus.n42 minus.n41 161.3
R223 minus.n40 minus.n29 161.3
R224 minus.n39 minus.n38 161.3
R225 minus.n37 minus.n30 161.3
R226 minus.n36 minus.n35 161.3
R227 minus.n34 minus.n31 161.3
R228 minus.n8 minus.n7 44.9377
R229 minus.n34 minus.n33 44.9377
R230 minus.n24 minus.n23 37.246
R231 minus.n50 minus.n49 37.246
R232 minus.n52 minus.n25 36.7391
R233 minus.n6 minus.n5 32.8641
R234 minus.n22 minus.n1 32.8641
R235 minus.n32 minus.n31 32.8641
R236 minus.n48 minus.n27 32.8641
R237 minus.n11 minus.n10 28.4823
R238 minus.n18 minus.n17 28.4823
R239 minus.n37 minus.n36 28.4823
R240 minus.n44 minus.n43 28.4823
R241 minus.n16 minus.n3 24.1005
R242 minus.n12 minus.n3 24.1005
R243 minus.n38 minus.n29 24.1005
R244 minus.n42 minus.n29 24.1005
R245 minus.n12 minus.n11 19.7187
R246 minus.n17 minus.n16 19.7187
R247 minus.n38 minus.n37 19.7187
R248 minus.n43 minus.n42 19.7187
R249 minus.n7 minus.n6 17.0522
R250 minus.n33 minus.n32 17.0522
R251 minus.n10 minus.n5 15.3369
R252 minus.n18 minus.n1 15.3369
R253 minus.n36 minus.n31 15.3369
R254 minus.n44 minus.n27 15.3369
R255 minus.n23 minus.n22 10.955
R256 minus.n49 minus.n48 10.955
R257 minus.n52 minus.n51 6.6558
R258 minus.n25 minus.n0 0.189894
R259 minus.n21 minus.n0 0.189894
R260 minus.n21 minus.n20 0.189894
R261 minus.n20 minus.n19 0.189894
R262 minus.n19 minus.n2 0.189894
R263 minus.n15 minus.n2 0.189894
R264 minus.n15 minus.n14 0.189894
R265 minus.n14 minus.n13 0.189894
R266 minus.n13 minus.n4 0.189894
R267 minus.n9 minus.n4 0.189894
R268 minus.n9 minus.n8 0.189894
R269 minus.n35 minus.n34 0.189894
R270 minus.n35 minus.n30 0.189894
R271 minus.n39 minus.n30 0.189894
R272 minus.n40 minus.n39 0.189894
R273 minus.n41 minus.n40 0.189894
R274 minus.n41 minus.n28 0.189894
R275 minus.n45 minus.n28 0.189894
R276 minus.n46 minus.n45 0.189894
R277 minus.n47 minus.n46 0.189894
R278 minus.n47 minus.n26 0.189894
R279 minus.n51 minus.n26 0.189894
R280 minus minus.n52 0.188
R281 drain_right.n9 drain_right.n7 66.4254
R282 drain_right.n5 drain_right.n3 66.4253
R283 drain_right.n2 drain_right.n0 66.4253
R284 drain_right.n9 drain_right.n8 65.5376
R285 drain_right.n11 drain_right.n10 65.5376
R286 drain_right.n13 drain_right.n12 65.5376
R287 drain_right.n5 drain_right.n4 65.5373
R288 drain_right.n2 drain_right.n1 65.5373
R289 drain_right drain_right.n6 30.3127
R290 drain_right drain_right.n13 6.54115
R291 drain_right.n3 drain_right.t8 2.2005
R292 drain_right.n3 drain_right.t13 2.2005
R293 drain_right.n4 drain_right.t4 2.2005
R294 drain_right.n4 drain_right.t10 2.2005
R295 drain_right.n1 drain_right.t7 2.2005
R296 drain_right.n1 drain_right.t6 2.2005
R297 drain_right.n0 drain_right.t0 2.2005
R298 drain_right.n0 drain_right.t1 2.2005
R299 drain_right.n7 drain_right.t15 2.2005
R300 drain_right.n7 drain_right.t9 2.2005
R301 drain_right.n8 drain_right.t3 2.2005
R302 drain_right.n8 drain_right.t11 2.2005
R303 drain_right.n10 drain_right.t2 2.2005
R304 drain_right.n10 drain_right.t12 2.2005
R305 drain_right.n12 drain_right.t5 2.2005
R306 drain_right.n12 drain_right.t14 2.2005
R307 drain_right.n13 drain_right.n11 0.888431
R308 drain_right.n11 drain_right.n9 0.888431
R309 drain_right.n6 drain_right.n5 0.389119
R310 drain_right.n6 drain_right.n2 0.389119
C0 minus drain_right 7.82625f
C1 drain_left drain_right 1.34352f
C2 source plus 7.98327f
C3 minus plus 5.79461f
C4 minus source 7.96923f
C5 plus drain_left 8.08089f
C6 plus drain_right 0.410755f
C7 source drain_left 15.712001f
C8 source drain_right 15.714201f
C9 minus drain_left 0.172697f
C10 drain_right a_n2570_n2688# 6.21433f
C11 drain_left a_n2570_n2688# 6.58649f
C12 source a_n2570_n2688# 7.57809f
C13 minus a_n2570_n2688# 10.05377f
C14 plus a_n2570_n2688# 11.66627f
C15 drain_right.t0 a_n2570_n2688# 0.19227f
C16 drain_right.t1 a_n2570_n2688# 0.19227f
C17 drain_right.n0 a_n2570_n2688# 1.68683f
C18 drain_right.t7 a_n2570_n2688# 0.19227f
C19 drain_right.t6 a_n2570_n2688# 0.19227f
C20 drain_right.n1 a_n2570_n2688# 1.68172f
C21 drain_right.n2 a_n2570_n2688# 0.706387f
C22 drain_right.t8 a_n2570_n2688# 0.19227f
C23 drain_right.t13 a_n2570_n2688# 0.19227f
C24 drain_right.n3 a_n2570_n2688# 1.68683f
C25 drain_right.t4 a_n2570_n2688# 0.19227f
C26 drain_right.t10 a_n2570_n2688# 0.19227f
C27 drain_right.n4 a_n2570_n2688# 1.68172f
C28 drain_right.n5 a_n2570_n2688# 0.706387f
C29 drain_right.n6 a_n2570_n2688# 1.31376f
C30 drain_right.t15 a_n2570_n2688# 0.19227f
C31 drain_right.t9 a_n2570_n2688# 0.19227f
C32 drain_right.n7 a_n2570_n2688# 1.68683f
C33 drain_right.t3 a_n2570_n2688# 0.19227f
C34 drain_right.t11 a_n2570_n2688# 0.19227f
C35 drain_right.n8 a_n2570_n2688# 1.68173f
C36 drain_right.n9 a_n2570_n2688# 0.74827f
C37 drain_right.t2 a_n2570_n2688# 0.19227f
C38 drain_right.t12 a_n2570_n2688# 0.19227f
C39 drain_right.n10 a_n2570_n2688# 1.68173f
C40 drain_right.n11 a_n2570_n2688# 0.371241f
C41 drain_right.t5 a_n2570_n2688# 0.19227f
C42 drain_right.t14 a_n2570_n2688# 0.19227f
C43 drain_right.n12 a_n2570_n2688# 1.68173f
C44 drain_right.n13 a_n2570_n2688# 0.610362f
C45 minus.n0 a_n2570_n2688# 0.040766f
C46 minus.n1 a_n2570_n2688# 0.009251f
C47 minus.t1 a_n2570_n2688# 0.736537f
C48 minus.n2 a_n2570_n2688# 0.040766f
C49 minus.n3 a_n2570_n2688# 0.009251f
C50 minus.t3 a_n2570_n2688# 0.736537f
C51 minus.n4 a_n2570_n2688# 0.040766f
C52 minus.n5 a_n2570_n2688# 0.009251f
C53 minus.t4 a_n2570_n2688# 0.736537f
C54 minus.t6 a_n2570_n2688# 0.75587f
C55 minus.t0 a_n2570_n2688# 0.736537f
C56 minus.n6 a_n2570_n2688# 0.31504f
C57 minus.n7 a_n2570_n2688# 0.293514f
C58 minus.n8 a_n2570_n2688# 0.172511f
C59 minus.n9 a_n2570_n2688# 0.040766f
C60 minus.n10 a_n2570_n2688# 0.309456f
C61 minus.n11 a_n2570_n2688# 0.009251f
C62 minus.t12 a_n2570_n2688# 0.736537f
C63 minus.n12 a_n2570_n2688# 0.309456f
C64 minus.n13 a_n2570_n2688# 0.040766f
C65 minus.n14 a_n2570_n2688# 0.040766f
C66 minus.n15 a_n2570_n2688# 0.040766f
C67 minus.n16 a_n2570_n2688# 0.309456f
C68 minus.n17 a_n2570_n2688# 0.009251f
C69 minus.t13 a_n2570_n2688# 0.736537f
C70 minus.n18 a_n2570_n2688# 0.309456f
C71 minus.n19 a_n2570_n2688# 0.040766f
C72 minus.n20 a_n2570_n2688# 0.040766f
C73 minus.n21 a_n2570_n2688# 0.040766f
C74 minus.n22 a_n2570_n2688# 0.309456f
C75 minus.n23 a_n2570_n2688# 0.009251f
C76 minus.t10 a_n2570_n2688# 0.736537f
C77 minus.n24 a_n2570_n2688# 0.308325f
C78 minus.n25 a_n2570_n2688# 1.47951f
C79 minus.n26 a_n2570_n2688# 0.040766f
C80 minus.n27 a_n2570_n2688# 0.009251f
C81 minus.n28 a_n2570_n2688# 0.040766f
C82 minus.n29 a_n2570_n2688# 0.009251f
C83 minus.n30 a_n2570_n2688# 0.040766f
C84 minus.n31 a_n2570_n2688# 0.009251f
C85 minus.t15 a_n2570_n2688# 0.75587f
C86 minus.t14 a_n2570_n2688# 0.736537f
C87 minus.n32 a_n2570_n2688# 0.31504f
C88 minus.n33 a_n2570_n2688# 0.293514f
C89 minus.n34 a_n2570_n2688# 0.172511f
C90 minus.n35 a_n2570_n2688# 0.040766f
C91 minus.t8 a_n2570_n2688# 0.736537f
C92 minus.n36 a_n2570_n2688# 0.309456f
C93 minus.n37 a_n2570_n2688# 0.009251f
C94 minus.t9 a_n2570_n2688# 0.736537f
C95 minus.n38 a_n2570_n2688# 0.309456f
C96 minus.n39 a_n2570_n2688# 0.040766f
C97 minus.n40 a_n2570_n2688# 0.040766f
C98 minus.n41 a_n2570_n2688# 0.040766f
C99 minus.t11 a_n2570_n2688# 0.736537f
C100 minus.n42 a_n2570_n2688# 0.309456f
C101 minus.n43 a_n2570_n2688# 0.009251f
C102 minus.t5 a_n2570_n2688# 0.736537f
C103 minus.n44 a_n2570_n2688# 0.309456f
C104 minus.n45 a_n2570_n2688# 0.040766f
C105 minus.n46 a_n2570_n2688# 0.040766f
C106 minus.n47 a_n2570_n2688# 0.040766f
C107 minus.t7 a_n2570_n2688# 0.736537f
C108 minus.n48 a_n2570_n2688# 0.309456f
C109 minus.n49 a_n2570_n2688# 0.009251f
C110 minus.t2 a_n2570_n2688# 0.736537f
C111 minus.n50 a_n2570_n2688# 0.308325f
C112 minus.n51 a_n2570_n2688# 0.281371f
C113 minus.n52 a_n2570_n2688# 1.78944f
C114 source.t25 a_n2570_n2688# 1.81247f
C115 source.n0 a_n2570_n2688# 1.08662f
C116 source.t22 a_n2570_n2688# 0.16997f
C117 source.t31 a_n2570_n2688# 0.16997f
C118 source.n1 a_n2570_n2688# 1.42288f
C119 source.n2 a_n2570_n2688# 0.359495f
C120 source.t23 a_n2570_n2688# 0.16997f
C121 source.t29 a_n2570_n2688# 0.16997f
C122 source.n3 a_n2570_n2688# 1.42288f
C123 source.n4 a_n2570_n2688# 0.359495f
C124 source.t21 a_n2570_n2688# 0.16997f
C125 source.t30 a_n2570_n2688# 0.16997f
C126 source.n5 a_n2570_n2688# 1.42288f
C127 source.n6 a_n2570_n2688# 0.359495f
C128 source.t28 a_n2570_n2688# 1.81247f
C129 source.n7 a_n2570_n2688# 0.401256f
C130 source.t10 a_n2570_n2688# 1.81247f
C131 source.n8 a_n2570_n2688# 0.401256f
C132 source.t11 a_n2570_n2688# 0.16997f
C133 source.t8 a_n2570_n2688# 0.16997f
C134 source.n9 a_n2570_n2688# 1.42288f
C135 source.n10 a_n2570_n2688# 0.359495f
C136 source.t7 a_n2570_n2688# 0.16997f
C137 source.t13 a_n2570_n2688# 0.16997f
C138 source.n11 a_n2570_n2688# 1.42288f
C139 source.n12 a_n2570_n2688# 0.359495f
C140 source.t12 a_n2570_n2688# 0.16997f
C141 source.t4 a_n2570_n2688# 0.16997f
C142 source.n13 a_n2570_n2688# 1.42288f
C143 source.n14 a_n2570_n2688# 0.359495f
C144 source.t3 a_n2570_n2688# 1.81247f
C145 source.n15 a_n2570_n2688# 1.44257f
C146 source.t20 a_n2570_n2688# 1.81247f
C147 source.n16 a_n2570_n2688# 1.44257f
C148 source.t16 a_n2570_n2688# 0.16997f
C149 source.t17 a_n2570_n2688# 0.16997f
C150 source.n17 a_n2570_n2688# 1.42287f
C151 source.n18 a_n2570_n2688# 0.359499f
C152 source.t26 a_n2570_n2688# 0.16997f
C153 source.t27 a_n2570_n2688# 0.16997f
C154 source.n19 a_n2570_n2688# 1.42287f
C155 source.n20 a_n2570_n2688# 0.359499f
C156 source.t24 a_n2570_n2688# 0.16997f
C157 source.t18 a_n2570_n2688# 0.16997f
C158 source.n21 a_n2570_n2688# 1.42287f
C159 source.n22 a_n2570_n2688# 0.359499f
C160 source.t19 a_n2570_n2688# 1.81247f
C161 source.n23 a_n2570_n2688# 0.401261f
C162 source.t15 a_n2570_n2688# 1.81247f
C163 source.n24 a_n2570_n2688# 0.401261f
C164 source.t5 a_n2570_n2688# 0.16997f
C165 source.t1 a_n2570_n2688# 0.16997f
C166 source.n25 a_n2570_n2688# 1.42287f
C167 source.n26 a_n2570_n2688# 0.359499f
C168 source.t2 a_n2570_n2688# 0.16997f
C169 source.t9 a_n2570_n2688# 0.16997f
C170 source.n27 a_n2570_n2688# 1.42287f
C171 source.n28 a_n2570_n2688# 0.359499f
C172 source.t0 a_n2570_n2688# 0.16997f
C173 source.t14 a_n2570_n2688# 0.16997f
C174 source.n29 a_n2570_n2688# 1.42287f
C175 source.n30 a_n2570_n2688# 0.359499f
C176 source.t6 a_n2570_n2688# 1.81247f
C177 source.n31 a_n2570_n2688# 0.557153f
C178 source.n32 a_n2570_n2688# 1.25838f
C179 drain_left.t0 a_n2570_n2688# 0.193852f
C180 drain_left.t8 a_n2570_n2688# 0.193852f
C181 drain_left.n0 a_n2570_n2688# 1.70071f
C182 drain_left.t12 a_n2570_n2688# 0.193852f
C183 drain_left.t4 a_n2570_n2688# 0.193852f
C184 drain_left.n1 a_n2570_n2688# 1.69556f
C185 drain_left.n2 a_n2570_n2688# 0.7122f
C186 drain_left.t5 a_n2570_n2688# 0.193852f
C187 drain_left.t10 a_n2570_n2688# 0.193852f
C188 drain_left.n3 a_n2570_n2688# 1.70071f
C189 drain_left.t3 a_n2570_n2688# 0.193852f
C190 drain_left.t2 a_n2570_n2688# 0.193852f
C191 drain_left.n4 a_n2570_n2688# 1.69556f
C192 drain_left.n5 a_n2570_n2688# 0.7122f
C193 drain_left.n6 a_n2570_n2688# 1.38001f
C194 drain_left.t15 a_n2570_n2688# 0.193852f
C195 drain_left.t11 a_n2570_n2688# 0.193852f
C196 drain_left.n7 a_n2570_n2688# 1.70071f
C197 drain_left.t13 a_n2570_n2688# 0.193852f
C198 drain_left.t7 a_n2570_n2688# 0.193852f
C199 drain_left.n8 a_n2570_n2688# 1.69556f
C200 drain_left.n9 a_n2570_n2688# 0.754421f
C201 drain_left.t1 a_n2570_n2688# 0.193852f
C202 drain_left.t9 a_n2570_n2688# 0.193852f
C203 drain_left.n10 a_n2570_n2688# 1.69556f
C204 drain_left.n11 a_n2570_n2688# 0.374296f
C205 drain_left.t14 a_n2570_n2688# 0.193852f
C206 drain_left.t6 a_n2570_n2688# 0.193852f
C207 drain_left.n12 a_n2570_n2688# 1.69556f
C208 drain_left.n13 a_n2570_n2688# 0.615391f
C209 plus.n0 a_n2570_n2688# 0.04149f
C210 plus.t6 a_n2570_n2688# 0.749627f
C211 plus.t0 a_n2570_n2688# 0.749627f
C212 plus.n1 a_n2570_n2688# 0.04149f
C213 plus.t9 a_n2570_n2688# 0.749627f
C214 plus.n2 a_n2570_n2688# 0.314956f
C215 plus.n3 a_n2570_n2688# 0.04149f
C216 plus.t2 a_n2570_n2688# 0.749627f
C217 plus.t8 a_n2570_n2688# 0.749627f
C218 plus.n4 a_n2570_n2688# 0.314956f
C219 plus.n5 a_n2570_n2688# 0.04149f
C220 plus.t1 a_n2570_n2688# 0.749627f
C221 plus.t10 a_n2570_n2688# 0.749627f
C222 plus.n6 a_n2570_n2688# 0.320639f
C223 plus.t3 a_n2570_n2688# 0.769305f
C224 plus.n7 a_n2570_n2688# 0.298731f
C225 plus.n8 a_n2570_n2688# 0.175577f
C226 plus.n9 a_n2570_n2688# 0.009415f
C227 plus.n10 a_n2570_n2688# 0.314956f
C228 plus.n11 a_n2570_n2688# 0.009415f
C229 plus.n12 a_n2570_n2688# 0.04149f
C230 plus.n13 a_n2570_n2688# 0.04149f
C231 plus.n14 a_n2570_n2688# 0.04149f
C232 plus.n15 a_n2570_n2688# 0.009415f
C233 plus.n16 a_n2570_n2688# 0.314956f
C234 plus.n17 a_n2570_n2688# 0.009415f
C235 plus.n18 a_n2570_n2688# 0.04149f
C236 plus.n19 a_n2570_n2688# 0.04149f
C237 plus.n20 a_n2570_n2688# 0.04149f
C238 plus.n21 a_n2570_n2688# 0.009415f
C239 plus.n22 a_n2570_n2688# 0.314956f
C240 plus.n23 a_n2570_n2688# 0.009415f
C241 plus.n24 a_n2570_n2688# 0.313805f
C242 plus.n25 a_n2570_n2688# 0.423168f
C243 plus.n26 a_n2570_n2688# 0.04149f
C244 plus.t11 a_n2570_n2688# 0.749627f
C245 plus.n27 a_n2570_n2688# 0.04149f
C246 plus.t15 a_n2570_n2688# 0.749627f
C247 plus.t14 a_n2570_n2688# 0.749627f
C248 plus.n28 a_n2570_n2688# 0.314956f
C249 plus.n29 a_n2570_n2688# 0.04149f
C250 plus.t5 a_n2570_n2688# 0.749627f
C251 plus.t4 a_n2570_n2688# 0.749627f
C252 plus.n30 a_n2570_n2688# 0.314956f
C253 plus.n31 a_n2570_n2688# 0.04149f
C254 plus.t7 a_n2570_n2688# 0.749627f
C255 plus.t13 a_n2570_n2688# 0.749627f
C256 plus.n32 a_n2570_n2688# 0.320639f
C257 plus.t12 a_n2570_n2688# 0.769305f
C258 plus.n33 a_n2570_n2688# 0.298731f
C259 plus.n34 a_n2570_n2688# 0.175577f
C260 plus.n35 a_n2570_n2688# 0.009415f
C261 plus.n36 a_n2570_n2688# 0.314956f
C262 plus.n37 a_n2570_n2688# 0.009415f
C263 plus.n38 a_n2570_n2688# 0.04149f
C264 plus.n39 a_n2570_n2688# 0.04149f
C265 plus.n40 a_n2570_n2688# 0.04149f
C266 plus.n41 a_n2570_n2688# 0.009415f
C267 plus.n42 a_n2570_n2688# 0.314956f
C268 plus.n43 a_n2570_n2688# 0.009415f
C269 plus.n44 a_n2570_n2688# 0.04149f
C270 plus.n45 a_n2570_n2688# 0.04149f
C271 plus.n46 a_n2570_n2688# 0.04149f
C272 plus.n47 a_n2570_n2688# 0.009415f
C273 plus.n48 a_n2570_n2688# 0.314956f
C274 plus.n49 a_n2570_n2688# 0.009415f
C275 plus.n50 a_n2570_n2688# 0.313805f
C276 plus.n51 a_n2570_n2688# 1.32069f
.ends

