* NGSPICE file created from diffpair243.ext - technology: sky130A

.subckt diffpair243 minus drain_right drain_left source plus
X0 source.t12 plus.t0 drain_left.t0 a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X1 a_n1366_n2088# a_n1366_n2088# a_n1366_n2088# a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=22.8 ps=103.6 w=6 l=0.15
X2 a_n1366_n2088# a_n1366_n2088# a_n1366_n2088# a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X3 drain_left.t1 plus.t1 source.t11 a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X4 a_n1366_n2088# a_n1366_n2088# a_n1366_n2088# a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X5 drain_right.t7 minus.t0 source.t1 a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X6 source.t10 plus.t2 drain_left.t2 a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X7 source.t0 minus.t1 drain_right.t6 a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X8 a_n1366_n2088# a_n1366_n2088# a_n1366_n2088# a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X9 source.t13 minus.t2 drain_right.t5 a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X10 drain_right.t4 minus.t3 source.t14 a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X11 drain_right.t3 minus.t4 source.t15 a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X12 source.t3 minus.t5 drain_right.t2 a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X13 source.t9 plus.t3 drain_left.t3 a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X14 drain_right.t1 minus.t6 source.t2 a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X15 source.t4 minus.t7 drain_right.t0 a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X16 drain_left.t4 plus.t4 source.t8 a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X17 source.t7 plus.t5 drain_left.t5 a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X18 drain_left.t6 plus.t6 source.t6 a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X19 drain_left.t7 plus.t7 source.t5 a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
R0 plus.n1 plus.t3 1242.25
R1 plus.n5 plus.t4 1242.25
R2 plus.n8 plus.t1 1242.25
R3 plus.n12 plus.t0 1242.25
R4 plus.n2 plus.t7 1172.87
R5 plus.n4 plus.t5 1172.87
R6 plus.n9 plus.t2 1172.87
R7 plus.n11 plus.t6 1172.87
R8 plus.n1 plus.n0 161.489
R9 plus.n8 plus.n7 161.489
R10 plus.n3 plus.n0 161.3
R11 plus.n6 plus.n5 161.3
R12 plus.n10 plus.n7 161.3
R13 plus.n13 plus.n12 161.3
R14 plus.n3 plus.n2 47.4702
R15 plus.n4 plus.n3 47.4702
R16 plus.n11 plus.n10 47.4702
R17 plus.n10 plus.n9 47.4702
R18 plus plus.n13 25.9839
R19 plus.n2 plus.n1 25.5611
R20 plus.n5 plus.n4 25.5611
R21 plus.n12 plus.n11 25.5611
R22 plus.n9 plus.n8 25.5611
R23 plus plus.n6 9.95126
R24 plus.n6 plus.n0 0.189894
R25 plus.n13 plus.n7 0.189894
R26 drain_left.n5 drain_left.n3 67.7512
R27 drain_left.n2 drain_left.n1 67.4155
R28 drain_left.n2 drain_left.n0 67.4155
R29 drain_left.n5 drain_left.n4 67.1907
R30 drain_left drain_left.n2 24.7828
R31 drain_left drain_left.n5 6.21356
R32 drain_left.n1 drain_left.t2 5.0005
R33 drain_left.n1 drain_left.t1 5.0005
R34 drain_left.n0 drain_left.t0 5.0005
R35 drain_left.n0 drain_left.t6 5.0005
R36 drain_left.n4 drain_left.t5 5.0005
R37 drain_left.n4 drain_left.t4 5.0005
R38 drain_left.n3 drain_left.t3 5.0005
R39 drain_left.n3 drain_left.t7 5.0005
R40 source.n3 source.t9 55.512
R41 source.n4 source.t14 55.512
R42 source.n7 source.t3 55.512
R43 source.n0 source.t8 55.5119
R44 source.n15 source.t15 55.5119
R45 source.n12 source.t4 55.5119
R46 source.n11 source.t11 55.5119
R47 source.n8 source.t12 55.5119
R48 source.n2 source.n1 50.512
R49 source.n6 source.n5 50.512
R50 source.n14 source.n13 50.5119
R51 source.n10 source.n9 50.5119
R52 source.n8 source.n7 17.3026
R53 source.n16 source.n0 11.7595
R54 source.n16 source.n15 5.5436
R55 source.n13 source.t1 5.0005
R56 source.n13 source.t0 5.0005
R57 source.n9 source.t6 5.0005
R58 source.n9 source.t10 5.0005
R59 source.n1 source.t5 5.0005
R60 source.n1 source.t7 5.0005
R61 source.n5 source.t2 5.0005
R62 source.n5 source.t13 5.0005
R63 source.n7 source.n6 0.560845
R64 source.n6 source.n4 0.560845
R65 source.n3 source.n2 0.560845
R66 source.n2 source.n0 0.560845
R67 source.n10 source.n8 0.560845
R68 source.n11 source.n10 0.560845
R69 source.n14 source.n12 0.560845
R70 source.n15 source.n14 0.560845
R71 source.n4 source.n3 0.470328
R72 source.n12 source.n11 0.470328
R73 source source.n16 0.188
R74 minus.n5 minus.t5 1242.25
R75 minus.n1 minus.t3 1242.25
R76 minus.n12 minus.t4 1242.25
R77 minus.n8 minus.t7 1242.25
R78 minus.n4 minus.t6 1172.87
R79 minus.n2 minus.t2 1172.87
R80 minus.n11 minus.t1 1172.87
R81 minus.n9 minus.t0 1172.87
R82 minus.n1 minus.n0 161.489
R83 minus.n8 minus.n7 161.489
R84 minus.n6 minus.n5 161.3
R85 minus.n3 minus.n0 161.3
R86 minus.n13 minus.n12 161.3
R87 minus.n10 minus.n7 161.3
R88 minus.n4 minus.n3 47.4702
R89 minus.n3 minus.n2 47.4702
R90 minus.n10 minus.n9 47.4702
R91 minus.n11 minus.n10 47.4702
R92 minus.n14 minus.n6 29.83
R93 minus.n5 minus.n4 25.5611
R94 minus.n2 minus.n1 25.5611
R95 minus.n9 minus.n8 25.5611
R96 minus.n12 minus.n11 25.5611
R97 minus.n14 minus.n13 6.58005
R98 minus.n6 minus.n0 0.189894
R99 minus.n13 minus.n7 0.189894
R100 minus minus.n14 0.188
R101 drain_right.n5 drain_right.n3 67.751
R102 drain_right.n2 drain_right.n1 67.4155
R103 drain_right.n2 drain_right.n0 67.4155
R104 drain_right.n5 drain_right.n4 67.1908
R105 drain_right drain_right.n2 24.2296
R106 drain_right drain_right.n5 6.21356
R107 drain_right.n1 drain_right.t6 5.0005
R108 drain_right.n1 drain_right.t3 5.0005
R109 drain_right.n0 drain_right.t0 5.0005
R110 drain_right.n0 drain_right.t7 5.0005
R111 drain_right.n3 drain_right.t5 5.0005
R112 drain_right.n3 drain_right.t4 5.0005
R113 drain_right.n4 drain_right.t2 5.0005
R114 drain_right.n4 drain_right.t1 5.0005
C0 drain_right source 9.38169f
C1 drain_right plus 0.282599f
C2 drain_right minus 1.26502f
C3 source drain_left 9.38236f
C4 drain_left plus 1.39442f
C5 drain_left minus 0.170499f
C6 source plus 1.05199f
C7 source minus 1.03797f
C8 minus plus 3.72396f
C9 drain_right drain_left 0.640281f
C10 drain_right a_n1366_n2088# 3.91311f
C11 drain_left a_n1366_n2088# 4.08544f
C12 source a_n1366_n2088# 5.174729f
C13 minus a_n1366_n2088# 4.517116f
C14 plus a_n1366_n2088# 5.47999f
C15 drain_right.t0 a_n1366_n2088# 0.175183f
C16 drain_right.t7 a_n1366_n2088# 0.175183f
C17 drain_right.n0 a_n1366_n2088# 1.08431f
C18 drain_right.t6 a_n1366_n2088# 0.175183f
C19 drain_right.t3 a_n1366_n2088# 0.175183f
C20 drain_right.n1 a_n1366_n2088# 1.08431f
C21 drain_right.n2 a_n1366_n2088# 1.2507f
C22 drain_right.t5 a_n1366_n2088# 0.175183f
C23 drain_right.t4 a_n1366_n2088# 0.175183f
C24 drain_right.n3 a_n1366_n2088# 1.08585f
C25 drain_right.t2 a_n1366_n2088# 0.175183f
C26 drain_right.t1 a_n1366_n2088# 0.175183f
C27 drain_right.n4 a_n1366_n2088# 1.08341f
C28 drain_right.n5 a_n1366_n2088# 0.782975f
C29 minus.n0 a_n1366_n2088# 0.084448f
C30 minus.t5 a_n1366_n2088# 0.094239f
C31 minus.t6 a_n1366_n2088# 0.091434f
C32 minus.t2 a_n1366_n2088# 0.091434f
C33 minus.t3 a_n1366_n2088# 0.094239f
C34 minus.n1 a_n1366_n2088# 0.062593f
C35 minus.n2 a_n1366_n2088# 0.047466f
C36 minus.n3 a_n1366_n2088# 0.015126f
C37 minus.n4 a_n1366_n2088# 0.047466f
C38 minus.n5 a_n1366_n2088# 0.062536f
C39 minus.n6 a_n1366_n2088# 0.921295f
C40 minus.n7 a_n1366_n2088# 0.084448f
C41 minus.t1 a_n1366_n2088# 0.091434f
C42 minus.t0 a_n1366_n2088# 0.091434f
C43 minus.t7 a_n1366_n2088# 0.094239f
C44 minus.n8 a_n1366_n2088# 0.062593f
C45 minus.n9 a_n1366_n2088# 0.047466f
C46 minus.n10 a_n1366_n2088# 0.015126f
C47 minus.n11 a_n1366_n2088# 0.047466f
C48 minus.t4 a_n1366_n2088# 0.094239f
C49 minus.n12 a_n1366_n2088# 0.062536f
C50 minus.n13 a_n1366_n2088# 0.239816f
C51 minus.n14 a_n1366_n2088# 1.13351f
C52 source.t8 a_n1366_n2088# 0.99784f
C53 source.n0 a_n1366_n2088# 0.734087f
C54 source.t5 a_n1366_n2088# 0.142065f
C55 source.t7 a_n1366_n2088# 0.142065f
C56 source.n1 a_n1366_n2088# 0.826838f
C57 source.n2 a_n1366_n2088# 0.256787f
C58 source.t9 a_n1366_n2088# 0.997845f
C59 source.n3 a_n1366_n2088# 0.335731f
C60 source.t14 a_n1366_n2088# 0.997845f
C61 source.n4 a_n1366_n2088# 0.335731f
C62 source.t2 a_n1366_n2088# 0.142065f
C63 source.t13 a_n1366_n2088# 0.142065f
C64 source.n5 a_n1366_n2088# 0.826838f
C65 source.n6 a_n1366_n2088# 0.256787f
C66 source.t3 a_n1366_n2088# 0.997845f
C67 source.n7 a_n1366_n2088# 0.988984f
C68 source.t12 a_n1366_n2088# 0.99784f
C69 source.n8 a_n1366_n2088# 0.988989f
C70 source.t6 a_n1366_n2088# 0.142065f
C71 source.t10 a_n1366_n2088# 0.142065f
C72 source.n9 a_n1366_n2088# 0.826833f
C73 source.n10 a_n1366_n2088# 0.256792f
C74 source.t11 a_n1366_n2088# 0.99784f
C75 source.n11 a_n1366_n2088# 0.335736f
C76 source.t4 a_n1366_n2088# 0.99784f
C77 source.n12 a_n1366_n2088# 0.335736f
C78 source.t1 a_n1366_n2088# 0.142065f
C79 source.t0 a_n1366_n2088# 0.142065f
C80 source.n13 a_n1366_n2088# 0.826833f
C81 source.n14 a_n1366_n2088# 0.256792f
C82 source.t15 a_n1366_n2088# 0.99784f
C83 source.n15 a_n1366_n2088# 0.448246f
C84 source.n16 a_n1366_n2088# 0.809712f
C85 drain_left.t0 a_n1366_n2088# 0.173423f
C86 drain_left.t6 a_n1366_n2088# 0.173423f
C87 drain_left.n0 a_n1366_n2088# 1.07342f
C88 drain_left.t2 a_n1366_n2088# 0.173423f
C89 drain_left.t1 a_n1366_n2088# 0.173423f
C90 drain_left.n1 a_n1366_n2088# 1.07342f
C91 drain_left.n2 a_n1366_n2088# 1.28754f
C92 drain_left.t3 a_n1366_n2088# 0.173423f
C93 drain_left.t7 a_n1366_n2088# 0.173423f
C94 drain_left.n3 a_n1366_n2088# 1.07495f
C95 drain_left.t5 a_n1366_n2088# 0.173423f
C96 drain_left.t4 a_n1366_n2088# 0.173423f
C97 drain_left.n4 a_n1366_n2088# 1.07252f
C98 drain_left.n5 a_n1366_n2088# 0.775109f
C99 plus.n0 a_n1366_n2088# 0.086126f
C100 plus.t5 a_n1366_n2088# 0.093251f
C101 plus.t7 a_n1366_n2088# 0.093251f
C102 plus.t3 a_n1366_n2088# 0.096112f
C103 plus.n1 a_n1366_n2088# 0.063837f
C104 plus.n2 a_n1366_n2088# 0.048409f
C105 plus.n3 a_n1366_n2088# 0.015427f
C106 plus.n4 a_n1366_n2088# 0.048409f
C107 plus.t4 a_n1366_n2088# 0.096112f
C108 plus.n5 a_n1366_n2088# 0.063779f
C109 plus.n6 a_n1366_n2088# 0.318751f
C110 plus.n7 a_n1366_n2088# 0.086126f
C111 plus.t0 a_n1366_n2088# 0.096112f
C112 plus.t6 a_n1366_n2088# 0.093251f
C113 plus.t2 a_n1366_n2088# 0.093251f
C114 plus.t1 a_n1366_n2088# 0.096112f
C115 plus.n8 a_n1366_n2088# 0.063837f
C116 plus.n9 a_n1366_n2088# 0.048409f
C117 plus.n10 a_n1366_n2088# 0.015427f
C118 plus.n11 a_n1366_n2088# 0.048409f
C119 plus.n12 a_n1366_n2088# 0.063779f
C120 plus.n13 a_n1366_n2088# 0.850239f
.ends

