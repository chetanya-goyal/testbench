* NGSPICE file created from diffpair99.ext - technology: sky130A

.subckt diffpair99 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t46 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X1 source.t20 minus.t0 drain_right.t23 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X2 drain_right.t22 minus.t1 source.t19 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X3 source.t47 plus.t1 drain_left.t22 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X4 source.t33 plus.t2 drain_left.t21 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X5 drain_right.t21 minus.t2 source.t18 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X6 drain_right.t20 minus.t3 source.t17 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X7 source.t44 plus.t3 drain_left.t20 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X8 source.t45 plus.t4 drain_left.t19 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X9 a_n2094_n1288# a_n2094_n1288# a_n2094_n1288# a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.2
X10 source.t14 minus.t4 drain_right.t19 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X11 drain_right.t18 minus.t5 source.t21 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X12 source.t43 plus.t5 drain_left.t18 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X13 drain_left.t17 plus.t6 source.t27 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X14 drain_left.t16 plus.t7 source.t38 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X15 source.t5 minus.t6 drain_right.t17 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X16 source.t7 minus.t7 drain_right.t16 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X17 drain_left.t15 plus.t8 source.t41 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X18 drain_left.t14 plus.t9 source.t42 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X19 source.t10 minus.t8 drain_right.t15 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X20 drain_right.t14 minus.t9 source.t16 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X21 source.t0 minus.t10 drain_right.t13 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X22 drain_left.t13 plus.t10 source.t37 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X23 source.t35 plus.t11 drain_left.t12 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X24 a_n2094_n1288# a_n2094_n1288# a_n2094_n1288# a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X25 source.t15 minus.t11 drain_right.t12 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X26 drain_right.t11 minus.t12 source.t22 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X27 source.t26 plus.t12 drain_left.t11 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X28 a_n2094_n1288# a_n2094_n1288# a_n2094_n1288# a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X29 source.t2 minus.t13 drain_right.t10 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X30 drain_right.t9 minus.t14 source.t12 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X31 a_n2094_n1288# a_n2094_n1288# a_n2094_n1288# a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X32 drain_left.t10 plus.t13 source.t36 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X33 drain_right.t8 minus.t15 source.t3 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X34 drain_right.t7 minus.t16 source.t4 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X35 source.t34 plus.t14 drain_left.t9 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X36 source.t30 plus.t15 drain_left.t8 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X37 drain_right.t6 minus.t17 source.t6 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X38 source.t8 minus.t18 drain_right.t5 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X39 source.t25 plus.t16 drain_left.t7 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X40 drain_left.t6 plus.t17 source.t24 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X41 drain_right.t4 minus.t19 source.t11 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X42 source.t28 plus.t18 drain_left.t5 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X43 source.t1 minus.t20 drain_right.t3 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X44 source.t23 minus.t21 drain_right.t2 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X45 source.t9 minus.t22 drain_right.t1 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X46 drain_left.t4 plus.t19 source.t31 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X47 drain_left.t3 plus.t20 source.t29 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X48 drain_left.t2 plus.t21 source.t32 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X49 source.t39 plus.t22 drain_left.t1 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X50 drain_right.t0 minus.t23 source.t13 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X51 drain_left.t0 plus.t23 source.t40 a_n2094_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
R0 plus.n6 plus.t11 458.265
R1 plus.n29 plus.t19 458.265
R2 plus.n37 plus.t20 458.265
R3 plus.n60 plus.t14 458.265
R4 plus.n7 plus.t6 397.651
R5 plus.n5 plus.t22 397.651
R6 plus.n12 plus.t17 397.651
R7 plus.n14 plus.t16 397.651
R8 plus.n3 plus.t10 397.651
R9 plus.n19 plus.t5 397.651
R10 plus.n21 plus.t21 397.651
R11 plus.n1 plus.t15 397.651
R12 plus.n26 plus.t8 397.651
R13 plus.n28 plus.t2 397.651
R14 plus.n38 plus.t3 397.651
R15 plus.n36 plus.t13 397.651
R16 plus.n43 plus.t1 397.651
R17 plus.n45 plus.t7 397.651
R18 plus.n34 plus.t18 397.651
R19 plus.n50 plus.t0 397.651
R20 plus.n52 plus.t12 397.651
R21 plus.n32 plus.t23 397.651
R22 plus.n57 plus.t4 397.651
R23 plus.n59 plus.t9 397.651
R24 plus.n9 plus.n6 161.489
R25 plus.n40 plus.n37 161.489
R26 plus.n9 plus.n8 161.3
R27 plus.n11 plus.n10 161.3
R28 plus.n13 plus.n4 161.3
R29 plus.n16 plus.n15 161.3
R30 plus.n18 plus.n17 161.3
R31 plus.n20 plus.n2 161.3
R32 plus.n23 plus.n22 161.3
R33 plus.n25 plus.n24 161.3
R34 plus.n27 plus.n0 161.3
R35 plus.n30 plus.n29 161.3
R36 plus.n40 plus.n39 161.3
R37 plus.n42 plus.n41 161.3
R38 plus.n44 plus.n35 161.3
R39 plus.n47 plus.n46 161.3
R40 plus.n49 plus.n48 161.3
R41 plus.n51 plus.n33 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n56 plus.n55 161.3
R44 plus.n58 plus.n31 161.3
R45 plus.n61 plus.n60 161.3
R46 plus.n8 plus.n7 56.2338
R47 plus.n28 plus.n27 56.2338
R48 plus.n59 plus.n58 56.2338
R49 plus.n39 plus.n38 56.2338
R50 plus.n11 plus.n5 51.852
R51 plus.n26 plus.n25 51.852
R52 plus.n57 plus.n56 51.852
R53 plus.n42 plus.n36 51.852
R54 plus.n13 plus.n12 47.4702
R55 plus.n22 plus.n1 47.4702
R56 plus.n53 plus.n32 47.4702
R57 plus.n44 plus.n43 47.4702
R58 plus.n15 plus.n14 43.0884
R59 plus.n21 plus.n20 43.0884
R60 plus.n52 plus.n51 43.0884
R61 plus.n46 plus.n45 43.0884
R62 plus.n18 plus.n3 38.7066
R63 plus.n19 plus.n18 38.7066
R64 plus.n50 plus.n49 38.7066
R65 plus.n49 plus.n34 38.7066
R66 plus.n15 plus.n3 34.3247
R67 plus.n20 plus.n19 34.3247
R68 plus.n51 plus.n50 34.3247
R69 plus.n46 plus.n34 34.3247
R70 plus.n14 plus.n13 29.9429
R71 plus.n22 plus.n21 29.9429
R72 plus.n53 plus.n52 29.9429
R73 plus.n45 plus.n44 29.9429
R74 plus plus.n61 27.1354
R75 plus.n12 plus.n11 25.5611
R76 plus.n25 plus.n1 25.5611
R77 plus.n56 plus.n32 25.5611
R78 plus.n43 plus.n42 25.5611
R79 plus.n8 plus.n5 21.1793
R80 plus.n27 plus.n26 21.1793
R81 plus.n58 plus.n57 21.1793
R82 plus.n39 plus.n36 21.1793
R83 plus.n7 plus.n6 16.7975
R84 plus.n29 plus.n28 16.7975
R85 plus.n60 plus.n59 16.7975
R86 plus.n38 plus.n37 16.7975
R87 plus plus.n30 8.3452
R88 plus.n10 plus.n9 0.189894
R89 plus.n10 plus.n4 0.189894
R90 plus.n16 plus.n4 0.189894
R91 plus.n17 plus.n16 0.189894
R92 plus.n17 plus.n2 0.189894
R93 plus.n23 plus.n2 0.189894
R94 plus.n24 plus.n23 0.189894
R95 plus.n24 plus.n0 0.189894
R96 plus.n30 plus.n0 0.189894
R97 plus.n61 plus.n31 0.189894
R98 plus.n55 plus.n31 0.189894
R99 plus.n55 plus.n54 0.189894
R100 plus.n54 plus.n33 0.189894
R101 plus.n48 plus.n33 0.189894
R102 plus.n48 plus.n47 0.189894
R103 plus.n47 plus.n35 0.189894
R104 plus.n41 plus.n35 0.189894
R105 plus.n41 plus.n40 0.189894
R106 source.n98 source.n96 289.615
R107 source.n80 source.n78 289.615
R108 source.n72 source.n70 289.615
R109 source.n54 source.n52 289.615
R110 source.n2 source.n0 289.615
R111 source.n20 source.n18 289.615
R112 source.n28 source.n26 289.615
R113 source.n46 source.n44 289.615
R114 source.n99 source.n98 185
R115 source.n81 source.n80 185
R116 source.n73 source.n72 185
R117 source.n55 source.n54 185
R118 source.n3 source.n2 185
R119 source.n21 source.n20 185
R120 source.n29 source.n28 185
R121 source.n47 source.n46 185
R122 source.t6 source.n97 167.117
R123 source.t9 source.n79 167.117
R124 source.t29 source.n71 167.117
R125 source.t34 source.n53 167.117
R126 source.t31 source.n1 167.117
R127 source.t35 source.n19 167.117
R128 source.t3 source.n27 167.117
R129 source.t14 source.n45 167.117
R130 source.n9 source.n8 84.1169
R131 source.n11 source.n10 84.1169
R132 source.n13 source.n12 84.1169
R133 source.n15 source.n14 84.1169
R134 source.n17 source.n16 84.1169
R135 source.n35 source.n34 84.1169
R136 source.n37 source.n36 84.1169
R137 source.n39 source.n38 84.1169
R138 source.n41 source.n40 84.1169
R139 source.n43 source.n42 84.1169
R140 source.n95 source.n94 84.1168
R141 source.n93 source.n92 84.1168
R142 source.n91 source.n90 84.1168
R143 source.n89 source.n88 84.1168
R144 source.n87 source.n86 84.1168
R145 source.n69 source.n68 84.1168
R146 source.n67 source.n66 84.1168
R147 source.n65 source.n64 84.1168
R148 source.n63 source.n62 84.1168
R149 source.n61 source.n60 84.1168
R150 source.n98 source.t6 52.3082
R151 source.n80 source.t9 52.3082
R152 source.n72 source.t29 52.3082
R153 source.n54 source.t34 52.3082
R154 source.n2 source.t31 52.3082
R155 source.n20 source.t35 52.3082
R156 source.n28 source.t3 52.3082
R157 source.n46 source.t14 52.3082
R158 source.n103 source.n102 31.4096
R159 source.n85 source.n84 31.4096
R160 source.n77 source.n76 31.4096
R161 source.n59 source.n58 31.4096
R162 source.n7 source.n6 31.4096
R163 source.n25 source.n24 31.4096
R164 source.n33 source.n32 31.4096
R165 source.n51 source.n50 31.4096
R166 source.n59 source.n51 14.1689
R167 source.n94 source.t13 9.9005
R168 source.n94 source.t0 9.9005
R169 source.n92 source.t21 9.9005
R170 source.n92 source.t15 9.9005
R171 source.n90 source.t22 9.9005
R172 source.n90 source.t8 9.9005
R173 source.n88 source.t11 9.9005
R174 source.n88 source.t20 9.9005
R175 source.n86 source.t19 9.9005
R176 source.n86 source.t2 9.9005
R177 source.n68 source.t36 9.9005
R178 source.n68 source.t44 9.9005
R179 source.n66 source.t38 9.9005
R180 source.n66 source.t47 9.9005
R181 source.n64 source.t46 9.9005
R182 source.n64 source.t28 9.9005
R183 source.n62 source.t40 9.9005
R184 source.n62 source.t26 9.9005
R185 source.n60 source.t42 9.9005
R186 source.n60 source.t45 9.9005
R187 source.n8 source.t41 9.9005
R188 source.n8 source.t33 9.9005
R189 source.n10 source.t32 9.9005
R190 source.n10 source.t30 9.9005
R191 source.n12 source.t37 9.9005
R192 source.n12 source.t43 9.9005
R193 source.n14 source.t24 9.9005
R194 source.n14 source.t25 9.9005
R195 source.n16 source.t27 9.9005
R196 source.n16 source.t39 9.9005
R197 source.n34 source.t18 9.9005
R198 source.n34 source.t7 9.9005
R199 source.n36 source.t4 9.9005
R200 source.n36 source.t1 9.9005
R201 source.n38 source.t17 9.9005
R202 source.n38 source.t5 9.9005
R203 source.n40 source.t12 9.9005
R204 source.n40 source.t23 9.9005
R205 source.n42 source.t16 9.9005
R206 source.n42 source.t10 9.9005
R207 source.n99 source.n97 9.71174
R208 source.n81 source.n79 9.71174
R209 source.n73 source.n71 9.71174
R210 source.n55 source.n53 9.71174
R211 source.n3 source.n1 9.71174
R212 source.n21 source.n19 9.71174
R213 source.n29 source.n27 9.71174
R214 source.n47 source.n45 9.71174
R215 source.n102 source.n101 9.45567
R216 source.n84 source.n83 9.45567
R217 source.n76 source.n75 9.45567
R218 source.n58 source.n57 9.45567
R219 source.n6 source.n5 9.45567
R220 source.n24 source.n23 9.45567
R221 source.n32 source.n31 9.45567
R222 source.n50 source.n49 9.45567
R223 source.n101 source.n100 9.3005
R224 source.n83 source.n82 9.3005
R225 source.n75 source.n74 9.3005
R226 source.n57 source.n56 9.3005
R227 source.n5 source.n4 9.3005
R228 source.n23 source.n22 9.3005
R229 source.n31 source.n30 9.3005
R230 source.n49 source.n48 9.3005
R231 source.n104 source.n7 8.67749
R232 source.n102 source.n96 8.14595
R233 source.n84 source.n78 8.14595
R234 source.n76 source.n70 8.14595
R235 source.n58 source.n52 8.14595
R236 source.n6 source.n0 8.14595
R237 source.n24 source.n18 8.14595
R238 source.n32 source.n26 8.14595
R239 source.n50 source.n44 8.14595
R240 source.n100 source.n99 7.3702
R241 source.n82 source.n81 7.3702
R242 source.n74 source.n73 7.3702
R243 source.n56 source.n55 7.3702
R244 source.n4 source.n3 7.3702
R245 source.n22 source.n21 7.3702
R246 source.n30 source.n29 7.3702
R247 source.n48 source.n47 7.3702
R248 source.n100 source.n96 5.81868
R249 source.n82 source.n78 5.81868
R250 source.n74 source.n70 5.81868
R251 source.n56 source.n52 5.81868
R252 source.n4 source.n0 5.81868
R253 source.n22 source.n18 5.81868
R254 source.n30 source.n26 5.81868
R255 source.n48 source.n44 5.81868
R256 source.n104 source.n103 5.49188
R257 source.n101 source.n97 3.44771
R258 source.n83 source.n79 3.44771
R259 source.n75 source.n71 3.44771
R260 source.n57 source.n53 3.44771
R261 source.n5 source.n1 3.44771
R262 source.n23 source.n19 3.44771
R263 source.n31 source.n27 3.44771
R264 source.n49 source.n45 3.44771
R265 source.n33 source.n25 0.470328
R266 source.n85 source.n77 0.470328
R267 source.n51 source.n43 0.457397
R268 source.n43 source.n41 0.457397
R269 source.n41 source.n39 0.457397
R270 source.n39 source.n37 0.457397
R271 source.n37 source.n35 0.457397
R272 source.n35 source.n33 0.457397
R273 source.n25 source.n17 0.457397
R274 source.n17 source.n15 0.457397
R275 source.n15 source.n13 0.457397
R276 source.n13 source.n11 0.457397
R277 source.n11 source.n9 0.457397
R278 source.n9 source.n7 0.457397
R279 source.n61 source.n59 0.457397
R280 source.n63 source.n61 0.457397
R281 source.n65 source.n63 0.457397
R282 source.n67 source.n65 0.457397
R283 source.n69 source.n67 0.457397
R284 source.n77 source.n69 0.457397
R285 source.n87 source.n85 0.457397
R286 source.n89 source.n87 0.457397
R287 source.n91 source.n89 0.457397
R288 source.n93 source.n91 0.457397
R289 source.n95 source.n93 0.457397
R290 source.n103 source.n95 0.457397
R291 source source.n104 0.188
R292 drain_left.n13 drain_left.n11 101.252
R293 drain_left.n7 drain_left.n5 101.252
R294 drain_left.n2 drain_left.n0 101.252
R295 drain_left.n21 drain_left.n20 100.796
R296 drain_left.n19 drain_left.n18 100.796
R297 drain_left.n17 drain_left.n16 100.796
R298 drain_left.n15 drain_left.n14 100.796
R299 drain_left.n13 drain_left.n12 100.796
R300 drain_left.n7 drain_left.n6 100.796
R301 drain_left.n9 drain_left.n8 100.796
R302 drain_left.n4 drain_left.n3 100.796
R303 drain_left.n2 drain_left.n1 100.796
R304 drain_left drain_left.n10 24.1318
R305 drain_left.n5 drain_left.t20 9.9005
R306 drain_left.n5 drain_left.t3 9.9005
R307 drain_left.n6 drain_left.t22 9.9005
R308 drain_left.n6 drain_left.t10 9.9005
R309 drain_left.n8 drain_left.t5 9.9005
R310 drain_left.n8 drain_left.t16 9.9005
R311 drain_left.n3 drain_left.t11 9.9005
R312 drain_left.n3 drain_left.t23 9.9005
R313 drain_left.n1 drain_left.t19 9.9005
R314 drain_left.n1 drain_left.t0 9.9005
R315 drain_left.n0 drain_left.t9 9.9005
R316 drain_left.n0 drain_left.t14 9.9005
R317 drain_left.n20 drain_left.t21 9.9005
R318 drain_left.n20 drain_left.t4 9.9005
R319 drain_left.n18 drain_left.t8 9.9005
R320 drain_left.n18 drain_left.t15 9.9005
R321 drain_left.n16 drain_left.t18 9.9005
R322 drain_left.n16 drain_left.t2 9.9005
R323 drain_left.n14 drain_left.t7 9.9005
R324 drain_left.n14 drain_left.t13 9.9005
R325 drain_left.n12 drain_left.t1 9.9005
R326 drain_left.n12 drain_left.t6 9.9005
R327 drain_left.n11 drain_left.t12 9.9005
R328 drain_left.n11 drain_left.t17 9.9005
R329 drain_left drain_left.n21 6.11011
R330 drain_left.n9 drain_left.n7 0.457397
R331 drain_left.n4 drain_left.n2 0.457397
R332 drain_left.n15 drain_left.n13 0.457397
R333 drain_left.n17 drain_left.n15 0.457397
R334 drain_left.n19 drain_left.n17 0.457397
R335 drain_left.n21 drain_left.n19 0.457397
R336 drain_left.n10 drain_left.n9 0.173602
R337 drain_left.n10 drain_left.n4 0.173602
R338 minus.n29 minus.t4 458.265
R339 minus.n6 minus.t15 458.265
R340 minus.n60 minus.t17 458.265
R341 minus.n37 minus.t22 458.265
R342 minus.n28 minus.t9 397.651
R343 minus.n26 minus.t8 397.651
R344 minus.n1 minus.t14 397.651
R345 minus.n21 minus.t21 397.651
R346 minus.n19 minus.t3 397.651
R347 minus.n3 minus.t6 397.651
R348 minus.n14 minus.t16 397.651
R349 minus.n12 minus.t20 397.651
R350 minus.n5 minus.t2 397.651
R351 minus.n7 minus.t7 397.651
R352 minus.n59 minus.t10 397.651
R353 minus.n57 minus.t23 397.651
R354 minus.n32 minus.t11 397.651
R355 minus.n52 minus.t5 397.651
R356 minus.n50 minus.t18 397.651
R357 minus.n34 minus.t12 397.651
R358 minus.n45 minus.t0 397.651
R359 minus.n43 minus.t19 397.651
R360 minus.n36 minus.t13 397.651
R361 minus.n38 minus.t1 397.651
R362 minus.n9 minus.n6 161.489
R363 minus.n40 minus.n37 161.489
R364 minus.n30 minus.n29 161.3
R365 minus.n27 minus.n0 161.3
R366 minus.n25 minus.n24 161.3
R367 minus.n23 minus.n22 161.3
R368 minus.n20 minus.n2 161.3
R369 minus.n18 minus.n17 161.3
R370 minus.n16 minus.n15 161.3
R371 minus.n13 minus.n4 161.3
R372 minus.n11 minus.n10 161.3
R373 minus.n9 minus.n8 161.3
R374 minus.n61 minus.n60 161.3
R375 minus.n58 minus.n31 161.3
R376 minus.n56 minus.n55 161.3
R377 minus.n54 minus.n53 161.3
R378 minus.n51 minus.n33 161.3
R379 minus.n49 minus.n48 161.3
R380 minus.n47 minus.n46 161.3
R381 minus.n44 minus.n35 161.3
R382 minus.n42 minus.n41 161.3
R383 minus.n40 minus.n39 161.3
R384 minus.n28 minus.n27 56.2338
R385 minus.n8 minus.n7 56.2338
R386 minus.n39 minus.n38 56.2338
R387 minus.n59 minus.n58 56.2338
R388 minus.n26 minus.n25 51.852
R389 minus.n11 minus.n5 51.852
R390 minus.n42 minus.n36 51.852
R391 minus.n57 minus.n56 51.852
R392 minus.n22 minus.n1 47.4702
R393 minus.n13 minus.n12 47.4702
R394 minus.n44 minus.n43 47.4702
R395 minus.n53 minus.n32 47.4702
R396 minus.n21 minus.n20 43.0884
R397 minus.n15 minus.n14 43.0884
R398 minus.n46 minus.n45 43.0884
R399 minus.n52 minus.n51 43.0884
R400 minus.n19 minus.n18 38.7066
R401 minus.n18 minus.n3 38.7066
R402 minus.n49 minus.n34 38.7066
R403 minus.n50 minus.n49 38.7066
R404 minus.n20 minus.n19 34.3247
R405 minus.n15 minus.n3 34.3247
R406 minus.n46 minus.n34 34.3247
R407 minus.n51 minus.n50 34.3247
R408 minus.n22 minus.n21 29.9429
R409 minus.n14 minus.n13 29.9429
R410 minus.n45 minus.n44 29.9429
R411 minus.n53 minus.n52 29.9429
R412 minus.n62 minus.n30 29.4664
R413 minus.n25 minus.n1 25.5611
R414 minus.n12 minus.n11 25.5611
R415 minus.n43 minus.n42 25.5611
R416 minus.n56 minus.n32 25.5611
R417 minus.n27 minus.n26 21.1793
R418 minus.n8 minus.n5 21.1793
R419 minus.n39 minus.n36 21.1793
R420 minus.n58 minus.n57 21.1793
R421 minus.n29 minus.n28 16.7975
R422 minus.n7 minus.n6 16.7975
R423 minus.n38 minus.n37 16.7975
R424 minus.n60 minus.n59 16.7975
R425 minus.n62 minus.n61 6.48914
R426 minus.n30 minus.n0 0.189894
R427 minus.n24 minus.n0 0.189894
R428 minus.n24 minus.n23 0.189894
R429 minus.n23 minus.n2 0.189894
R430 minus.n17 minus.n2 0.189894
R431 minus.n17 minus.n16 0.189894
R432 minus.n16 minus.n4 0.189894
R433 minus.n10 minus.n4 0.189894
R434 minus.n10 minus.n9 0.189894
R435 minus.n41 minus.n40 0.189894
R436 minus.n41 minus.n35 0.189894
R437 minus.n47 minus.n35 0.189894
R438 minus.n48 minus.n47 0.189894
R439 minus.n48 minus.n33 0.189894
R440 minus.n54 minus.n33 0.189894
R441 minus.n55 minus.n54 0.189894
R442 minus.n55 minus.n31 0.189894
R443 minus.n61 minus.n31 0.189894
R444 minus minus.n62 0.188
R445 drain_right.n13 drain_right.n11 101.252
R446 drain_right.n7 drain_right.n5 101.252
R447 drain_right.n2 drain_right.n0 101.252
R448 drain_right.n13 drain_right.n12 100.796
R449 drain_right.n15 drain_right.n14 100.796
R450 drain_right.n17 drain_right.n16 100.796
R451 drain_right.n19 drain_right.n18 100.796
R452 drain_right.n21 drain_right.n20 100.796
R453 drain_right.n7 drain_right.n6 100.796
R454 drain_right.n9 drain_right.n8 100.796
R455 drain_right.n4 drain_right.n3 100.796
R456 drain_right.n2 drain_right.n1 100.796
R457 drain_right drain_right.n10 23.5786
R458 drain_right.n5 drain_right.t13 9.9005
R459 drain_right.n5 drain_right.t6 9.9005
R460 drain_right.n6 drain_right.t12 9.9005
R461 drain_right.n6 drain_right.t0 9.9005
R462 drain_right.n8 drain_right.t5 9.9005
R463 drain_right.n8 drain_right.t18 9.9005
R464 drain_right.n3 drain_right.t23 9.9005
R465 drain_right.n3 drain_right.t11 9.9005
R466 drain_right.n1 drain_right.t10 9.9005
R467 drain_right.n1 drain_right.t4 9.9005
R468 drain_right.n0 drain_right.t1 9.9005
R469 drain_right.n0 drain_right.t22 9.9005
R470 drain_right.n11 drain_right.t16 9.9005
R471 drain_right.n11 drain_right.t8 9.9005
R472 drain_right.n12 drain_right.t3 9.9005
R473 drain_right.n12 drain_right.t21 9.9005
R474 drain_right.n14 drain_right.t17 9.9005
R475 drain_right.n14 drain_right.t7 9.9005
R476 drain_right.n16 drain_right.t2 9.9005
R477 drain_right.n16 drain_right.t20 9.9005
R478 drain_right.n18 drain_right.t15 9.9005
R479 drain_right.n18 drain_right.t9 9.9005
R480 drain_right.n20 drain_right.t19 9.9005
R481 drain_right.n20 drain_right.t14 9.9005
R482 drain_right drain_right.n21 6.11011
R483 drain_right.n9 drain_right.n7 0.457397
R484 drain_right.n4 drain_right.n2 0.457397
R485 drain_right.n21 drain_right.n19 0.457397
R486 drain_right.n19 drain_right.n17 0.457397
R487 drain_right.n17 drain_right.n15 0.457397
R488 drain_right.n15 drain_right.n13 0.457397
R489 drain_right.n10 drain_right.n9 0.173602
R490 drain_right.n10 drain_right.n4 0.173602
C0 drain_left drain_right 1.11966f
C1 minus plus 3.92245f
C2 source drain_right 12.0035f
C3 minus drain_right 1.57508f
C4 source drain_left 12.003201f
C5 drain_right plus 0.366634f
C6 minus drain_left 0.177815f
C7 drain_left plus 1.78022f
C8 source minus 1.79046f
C9 source plus 1.80442f
C10 drain_right a_n2094_n1288# 4.64399f
C11 drain_left a_n2094_n1288# 4.94032f
C12 source a_n2094_n1288# 3.253778f
C13 minus a_n2094_n1288# 7.340168f
C14 plus a_n2094_n1288# 7.981494f
C15 drain_right.t1 a_n2094_n1288# 0.050259f
C16 drain_right.t22 a_n2094_n1288# 0.050259f
C17 drain_right.n0 a_n2094_n1288# 0.317324f
C18 drain_right.t10 a_n2094_n1288# 0.050259f
C19 drain_right.t4 a_n2094_n1288# 0.050259f
C20 drain_right.n1 a_n2094_n1288# 0.315745f
C21 drain_right.n2 a_n2094_n1288# 0.685296f
C22 drain_right.t23 a_n2094_n1288# 0.050259f
C23 drain_right.t11 a_n2094_n1288# 0.050259f
C24 drain_right.n3 a_n2094_n1288# 0.315745f
C25 drain_right.n4 a_n2094_n1288# 0.312212f
C26 drain_right.t13 a_n2094_n1288# 0.050259f
C27 drain_right.t6 a_n2094_n1288# 0.050259f
C28 drain_right.n5 a_n2094_n1288# 0.317324f
C29 drain_right.t12 a_n2094_n1288# 0.050259f
C30 drain_right.t0 a_n2094_n1288# 0.050259f
C31 drain_right.n6 a_n2094_n1288# 0.315745f
C32 drain_right.n7 a_n2094_n1288# 0.685296f
C33 drain_right.t5 a_n2094_n1288# 0.050259f
C34 drain_right.t18 a_n2094_n1288# 0.050259f
C35 drain_right.n8 a_n2094_n1288# 0.315745f
C36 drain_right.n9 a_n2094_n1288# 0.312212f
C37 drain_right.n10 a_n2094_n1288# 0.914422f
C38 drain_right.t16 a_n2094_n1288# 0.050259f
C39 drain_right.t8 a_n2094_n1288# 0.050259f
C40 drain_right.n11 a_n2094_n1288# 0.317325f
C41 drain_right.t3 a_n2094_n1288# 0.050259f
C42 drain_right.t21 a_n2094_n1288# 0.050259f
C43 drain_right.n12 a_n2094_n1288# 0.315747f
C44 drain_right.n13 a_n2094_n1288# 0.685294f
C45 drain_right.t17 a_n2094_n1288# 0.050259f
C46 drain_right.t7 a_n2094_n1288# 0.050259f
C47 drain_right.n14 a_n2094_n1288# 0.315747f
C48 drain_right.n15 a_n2094_n1288# 0.337032f
C49 drain_right.t2 a_n2094_n1288# 0.050259f
C50 drain_right.t20 a_n2094_n1288# 0.050259f
C51 drain_right.n16 a_n2094_n1288# 0.315747f
C52 drain_right.n17 a_n2094_n1288# 0.337032f
C53 drain_right.t15 a_n2094_n1288# 0.050259f
C54 drain_right.t9 a_n2094_n1288# 0.050259f
C55 drain_right.n18 a_n2094_n1288# 0.315747f
C56 drain_right.n19 a_n2094_n1288# 0.337032f
C57 drain_right.t19 a_n2094_n1288# 0.050259f
C58 drain_right.t14 a_n2094_n1288# 0.050259f
C59 drain_right.n20 a_n2094_n1288# 0.315747f
C60 drain_right.n21 a_n2094_n1288# 0.597289f
C61 minus.n0 a_n2094_n1288# 0.027346f
C62 minus.t4 a_n2094_n1288# 0.035789f
C63 minus.t9 a_n2094_n1288# 0.032187f
C64 minus.t8 a_n2094_n1288# 0.032187f
C65 minus.t14 a_n2094_n1288# 0.032187f
C66 minus.n1 a_n2094_n1288# 0.02529f
C67 minus.n2 a_n2094_n1288# 0.027346f
C68 minus.t21 a_n2094_n1288# 0.032187f
C69 minus.t3 a_n2094_n1288# 0.032187f
C70 minus.t6 a_n2094_n1288# 0.032187f
C71 minus.n3 a_n2094_n1288# 0.02529f
C72 minus.n4 a_n2094_n1288# 0.027346f
C73 minus.t16 a_n2094_n1288# 0.032187f
C74 minus.t20 a_n2094_n1288# 0.032187f
C75 minus.t2 a_n2094_n1288# 0.032187f
C76 minus.n5 a_n2094_n1288# 0.02529f
C77 minus.t15 a_n2094_n1288# 0.035789f
C78 minus.n6 a_n2094_n1288# 0.033247f
C79 minus.t7 a_n2094_n1288# 0.032187f
C80 minus.n7 a_n2094_n1288# 0.02529f
C81 minus.n8 a_n2094_n1288# 0.009577f
C82 minus.n9 a_n2094_n1288# 0.063586f
C83 minus.n10 a_n2094_n1288# 0.027346f
C84 minus.n11 a_n2094_n1288# 0.009577f
C85 minus.n12 a_n2094_n1288# 0.02529f
C86 minus.n13 a_n2094_n1288# 0.009577f
C87 minus.n14 a_n2094_n1288# 0.02529f
C88 minus.n15 a_n2094_n1288# 0.009577f
C89 minus.n16 a_n2094_n1288# 0.027346f
C90 minus.n17 a_n2094_n1288# 0.027346f
C91 minus.n18 a_n2094_n1288# 0.009577f
C92 minus.n19 a_n2094_n1288# 0.02529f
C93 minus.n20 a_n2094_n1288# 0.009577f
C94 minus.n21 a_n2094_n1288# 0.02529f
C95 minus.n22 a_n2094_n1288# 0.009577f
C96 minus.n23 a_n2094_n1288# 0.027346f
C97 minus.n24 a_n2094_n1288# 0.027346f
C98 minus.n25 a_n2094_n1288# 0.009577f
C99 minus.n26 a_n2094_n1288# 0.02529f
C100 minus.n27 a_n2094_n1288# 0.009577f
C101 minus.n28 a_n2094_n1288# 0.02529f
C102 minus.n29 a_n2094_n1288# 0.033205f
C103 minus.n30 a_n2094_n1288# 0.68954f
C104 minus.n31 a_n2094_n1288# 0.027346f
C105 minus.t10 a_n2094_n1288# 0.032187f
C106 minus.t23 a_n2094_n1288# 0.032187f
C107 minus.t11 a_n2094_n1288# 0.032187f
C108 minus.n32 a_n2094_n1288# 0.02529f
C109 minus.n33 a_n2094_n1288# 0.027346f
C110 minus.t5 a_n2094_n1288# 0.032187f
C111 minus.t18 a_n2094_n1288# 0.032187f
C112 minus.t12 a_n2094_n1288# 0.032187f
C113 minus.n34 a_n2094_n1288# 0.02529f
C114 minus.n35 a_n2094_n1288# 0.027346f
C115 minus.t0 a_n2094_n1288# 0.032187f
C116 minus.t19 a_n2094_n1288# 0.032187f
C117 minus.t13 a_n2094_n1288# 0.032187f
C118 minus.n36 a_n2094_n1288# 0.02529f
C119 minus.t22 a_n2094_n1288# 0.035789f
C120 minus.n37 a_n2094_n1288# 0.033247f
C121 minus.t1 a_n2094_n1288# 0.032187f
C122 minus.n38 a_n2094_n1288# 0.02529f
C123 minus.n39 a_n2094_n1288# 0.009577f
C124 minus.n40 a_n2094_n1288# 0.063586f
C125 minus.n41 a_n2094_n1288# 0.027346f
C126 minus.n42 a_n2094_n1288# 0.009577f
C127 minus.n43 a_n2094_n1288# 0.02529f
C128 minus.n44 a_n2094_n1288# 0.009577f
C129 minus.n45 a_n2094_n1288# 0.02529f
C130 minus.n46 a_n2094_n1288# 0.009577f
C131 minus.n47 a_n2094_n1288# 0.027346f
C132 minus.n48 a_n2094_n1288# 0.027346f
C133 minus.n49 a_n2094_n1288# 0.009577f
C134 minus.n50 a_n2094_n1288# 0.02529f
C135 minus.n51 a_n2094_n1288# 0.009577f
C136 minus.n52 a_n2094_n1288# 0.02529f
C137 minus.n53 a_n2094_n1288# 0.009577f
C138 minus.n54 a_n2094_n1288# 0.027346f
C139 minus.n55 a_n2094_n1288# 0.027346f
C140 minus.n56 a_n2094_n1288# 0.009577f
C141 minus.n57 a_n2094_n1288# 0.02529f
C142 minus.n58 a_n2094_n1288# 0.009577f
C143 minus.n59 a_n2094_n1288# 0.02529f
C144 minus.t17 a_n2094_n1288# 0.035789f
C145 minus.n60 a_n2094_n1288# 0.033205f
C146 minus.n61 a_n2094_n1288# 0.178082f
C147 minus.n62 a_n2094_n1288# 0.851707f
C148 drain_left.t9 a_n2094_n1288# 0.049744f
C149 drain_left.t14 a_n2094_n1288# 0.049744f
C150 drain_left.n0 a_n2094_n1288# 0.314068f
C151 drain_left.t19 a_n2094_n1288# 0.049744f
C152 drain_left.t0 a_n2094_n1288# 0.049744f
C153 drain_left.n1 a_n2094_n1288# 0.312506f
C154 drain_left.n2 a_n2094_n1288# 0.678265f
C155 drain_left.t11 a_n2094_n1288# 0.049744f
C156 drain_left.t23 a_n2094_n1288# 0.049744f
C157 drain_left.n3 a_n2094_n1288# 0.312506f
C158 drain_left.n4 a_n2094_n1288# 0.309009f
C159 drain_left.t20 a_n2094_n1288# 0.049744f
C160 drain_left.t3 a_n2094_n1288# 0.049744f
C161 drain_left.n5 a_n2094_n1288# 0.314068f
C162 drain_left.t22 a_n2094_n1288# 0.049744f
C163 drain_left.t10 a_n2094_n1288# 0.049744f
C164 drain_left.n6 a_n2094_n1288# 0.312506f
C165 drain_left.n7 a_n2094_n1288# 0.678265f
C166 drain_left.t5 a_n2094_n1288# 0.049744f
C167 drain_left.t16 a_n2094_n1288# 0.049744f
C168 drain_left.n8 a_n2094_n1288# 0.312506f
C169 drain_left.n9 a_n2094_n1288# 0.309009f
C170 drain_left.n10 a_n2094_n1288# 0.966539f
C171 drain_left.t12 a_n2094_n1288# 0.049744f
C172 drain_left.t17 a_n2094_n1288# 0.049744f
C173 drain_left.n11 a_n2094_n1288# 0.314069f
C174 drain_left.t1 a_n2094_n1288# 0.049744f
C175 drain_left.t6 a_n2094_n1288# 0.049744f
C176 drain_left.n12 a_n2094_n1288# 0.312507f
C177 drain_left.n13 a_n2094_n1288# 0.678262f
C178 drain_left.t7 a_n2094_n1288# 0.049744f
C179 drain_left.t13 a_n2094_n1288# 0.049744f
C180 drain_left.n14 a_n2094_n1288# 0.312507f
C181 drain_left.n15 a_n2094_n1288# 0.333574f
C182 drain_left.t18 a_n2094_n1288# 0.049744f
C183 drain_left.t2 a_n2094_n1288# 0.049744f
C184 drain_left.n16 a_n2094_n1288# 0.312507f
C185 drain_left.n17 a_n2094_n1288# 0.333574f
C186 drain_left.t8 a_n2094_n1288# 0.049744f
C187 drain_left.t15 a_n2094_n1288# 0.049744f
C188 drain_left.n18 a_n2094_n1288# 0.312507f
C189 drain_left.n19 a_n2094_n1288# 0.333574f
C190 drain_left.t21 a_n2094_n1288# 0.049744f
C191 drain_left.t4 a_n2094_n1288# 0.049744f
C192 drain_left.n20 a_n2094_n1288# 0.312507f
C193 drain_left.n21 a_n2094_n1288# 0.59116f
C194 source.n0 a_n2094_n1288# 0.048831f
C195 source.n1 a_n2094_n1288# 0.108045f
C196 source.t31 a_n2094_n1288# 0.081082f
C197 source.n2 a_n2094_n1288# 0.08456f
C198 source.n3 a_n2094_n1288# 0.027259f
C199 source.n4 a_n2094_n1288# 0.017978f
C200 source.n5 a_n2094_n1288# 0.238157f
C201 source.n6 a_n2094_n1288# 0.05353f
C202 source.n7 a_n2094_n1288# 0.488602f
C203 source.t41 a_n2094_n1288# 0.052876f
C204 source.t33 a_n2094_n1288# 0.052876f
C205 source.n8 a_n2094_n1288# 0.282672f
C206 source.n9 a_n2094_n1288# 0.358614f
C207 source.t32 a_n2094_n1288# 0.052876f
C208 source.t30 a_n2094_n1288# 0.052876f
C209 source.n10 a_n2094_n1288# 0.282672f
C210 source.n11 a_n2094_n1288# 0.358614f
C211 source.t37 a_n2094_n1288# 0.052876f
C212 source.t43 a_n2094_n1288# 0.052876f
C213 source.n12 a_n2094_n1288# 0.282672f
C214 source.n13 a_n2094_n1288# 0.358614f
C215 source.t24 a_n2094_n1288# 0.052876f
C216 source.t25 a_n2094_n1288# 0.052876f
C217 source.n14 a_n2094_n1288# 0.282672f
C218 source.n15 a_n2094_n1288# 0.358614f
C219 source.t27 a_n2094_n1288# 0.052876f
C220 source.t39 a_n2094_n1288# 0.052876f
C221 source.n16 a_n2094_n1288# 0.282672f
C222 source.n17 a_n2094_n1288# 0.358614f
C223 source.n18 a_n2094_n1288# 0.048831f
C224 source.n19 a_n2094_n1288# 0.108045f
C225 source.t35 a_n2094_n1288# 0.081082f
C226 source.n20 a_n2094_n1288# 0.08456f
C227 source.n21 a_n2094_n1288# 0.027259f
C228 source.n22 a_n2094_n1288# 0.017978f
C229 source.n23 a_n2094_n1288# 0.238157f
C230 source.n24 a_n2094_n1288# 0.05353f
C231 source.n25 a_n2094_n1288# 0.127446f
C232 source.n26 a_n2094_n1288# 0.048831f
C233 source.n27 a_n2094_n1288# 0.108045f
C234 source.t3 a_n2094_n1288# 0.081082f
C235 source.n28 a_n2094_n1288# 0.08456f
C236 source.n29 a_n2094_n1288# 0.027259f
C237 source.n30 a_n2094_n1288# 0.017978f
C238 source.n31 a_n2094_n1288# 0.238157f
C239 source.n32 a_n2094_n1288# 0.05353f
C240 source.n33 a_n2094_n1288# 0.127446f
C241 source.t18 a_n2094_n1288# 0.052876f
C242 source.t7 a_n2094_n1288# 0.052876f
C243 source.n34 a_n2094_n1288# 0.282672f
C244 source.n35 a_n2094_n1288# 0.358614f
C245 source.t4 a_n2094_n1288# 0.052876f
C246 source.t1 a_n2094_n1288# 0.052876f
C247 source.n36 a_n2094_n1288# 0.282672f
C248 source.n37 a_n2094_n1288# 0.358614f
C249 source.t17 a_n2094_n1288# 0.052876f
C250 source.t5 a_n2094_n1288# 0.052876f
C251 source.n38 a_n2094_n1288# 0.282672f
C252 source.n39 a_n2094_n1288# 0.358614f
C253 source.t12 a_n2094_n1288# 0.052876f
C254 source.t23 a_n2094_n1288# 0.052876f
C255 source.n40 a_n2094_n1288# 0.282672f
C256 source.n41 a_n2094_n1288# 0.358614f
C257 source.t16 a_n2094_n1288# 0.052876f
C258 source.t10 a_n2094_n1288# 0.052876f
C259 source.n42 a_n2094_n1288# 0.282672f
C260 source.n43 a_n2094_n1288# 0.358614f
C261 source.n44 a_n2094_n1288# 0.048831f
C262 source.n45 a_n2094_n1288# 0.108045f
C263 source.t14 a_n2094_n1288# 0.081082f
C264 source.n46 a_n2094_n1288# 0.08456f
C265 source.n47 a_n2094_n1288# 0.027259f
C266 source.n48 a_n2094_n1288# 0.017978f
C267 source.n49 a_n2094_n1288# 0.238157f
C268 source.n50 a_n2094_n1288# 0.05353f
C269 source.n51 a_n2094_n1288# 0.798454f
C270 source.n52 a_n2094_n1288# 0.048831f
C271 source.n53 a_n2094_n1288# 0.108045f
C272 source.t34 a_n2094_n1288# 0.081082f
C273 source.n54 a_n2094_n1288# 0.08456f
C274 source.n55 a_n2094_n1288# 0.027259f
C275 source.n56 a_n2094_n1288# 0.017978f
C276 source.n57 a_n2094_n1288# 0.238157f
C277 source.n58 a_n2094_n1288# 0.05353f
C278 source.n59 a_n2094_n1288# 0.798454f
C279 source.t42 a_n2094_n1288# 0.052876f
C280 source.t45 a_n2094_n1288# 0.052876f
C281 source.n60 a_n2094_n1288# 0.282671f
C282 source.n61 a_n2094_n1288# 0.358615f
C283 source.t40 a_n2094_n1288# 0.052876f
C284 source.t26 a_n2094_n1288# 0.052876f
C285 source.n62 a_n2094_n1288# 0.282671f
C286 source.n63 a_n2094_n1288# 0.358615f
C287 source.t46 a_n2094_n1288# 0.052876f
C288 source.t28 a_n2094_n1288# 0.052876f
C289 source.n64 a_n2094_n1288# 0.282671f
C290 source.n65 a_n2094_n1288# 0.358615f
C291 source.t38 a_n2094_n1288# 0.052876f
C292 source.t47 a_n2094_n1288# 0.052876f
C293 source.n66 a_n2094_n1288# 0.282671f
C294 source.n67 a_n2094_n1288# 0.358615f
C295 source.t36 a_n2094_n1288# 0.052876f
C296 source.t44 a_n2094_n1288# 0.052876f
C297 source.n68 a_n2094_n1288# 0.282671f
C298 source.n69 a_n2094_n1288# 0.358615f
C299 source.n70 a_n2094_n1288# 0.048831f
C300 source.n71 a_n2094_n1288# 0.108045f
C301 source.t29 a_n2094_n1288# 0.081082f
C302 source.n72 a_n2094_n1288# 0.08456f
C303 source.n73 a_n2094_n1288# 0.027259f
C304 source.n74 a_n2094_n1288# 0.017978f
C305 source.n75 a_n2094_n1288# 0.238157f
C306 source.n76 a_n2094_n1288# 0.05353f
C307 source.n77 a_n2094_n1288# 0.127446f
C308 source.n78 a_n2094_n1288# 0.048831f
C309 source.n79 a_n2094_n1288# 0.108045f
C310 source.t9 a_n2094_n1288# 0.081082f
C311 source.n80 a_n2094_n1288# 0.08456f
C312 source.n81 a_n2094_n1288# 0.027259f
C313 source.n82 a_n2094_n1288# 0.017978f
C314 source.n83 a_n2094_n1288# 0.238157f
C315 source.n84 a_n2094_n1288# 0.05353f
C316 source.n85 a_n2094_n1288# 0.127446f
C317 source.t19 a_n2094_n1288# 0.052876f
C318 source.t2 a_n2094_n1288# 0.052876f
C319 source.n86 a_n2094_n1288# 0.282671f
C320 source.n87 a_n2094_n1288# 0.358615f
C321 source.t11 a_n2094_n1288# 0.052876f
C322 source.t20 a_n2094_n1288# 0.052876f
C323 source.n88 a_n2094_n1288# 0.282671f
C324 source.n89 a_n2094_n1288# 0.358615f
C325 source.t22 a_n2094_n1288# 0.052876f
C326 source.t8 a_n2094_n1288# 0.052876f
C327 source.n90 a_n2094_n1288# 0.282671f
C328 source.n91 a_n2094_n1288# 0.358615f
C329 source.t21 a_n2094_n1288# 0.052876f
C330 source.t15 a_n2094_n1288# 0.052876f
C331 source.n92 a_n2094_n1288# 0.282671f
C332 source.n93 a_n2094_n1288# 0.358615f
C333 source.t13 a_n2094_n1288# 0.052876f
C334 source.t0 a_n2094_n1288# 0.052876f
C335 source.n94 a_n2094_n1288# 0.282671f
C336 source.n95 a_n2094_n1288# 0.358615f
C337 source.n96 a_n2094_n1288# 0.048831f
C338 source.n97 a_n2094_n1288# 0.108045f
C339 source.t6 a_n2094_n1288# 0.081082f
C340 source.n98 a_n2094_n1288# 0.08456f
C341 source.n99 a_n2094_n1288# 0.027259f
C342 source.n100 a_n2094_n1288# 0.017978f
C343 source.n101 a_n2094_n1288# 0.238157f
C344 source.n102 a_n2094_n1288# 0.05353f
C345 source.n103 a_n2094_n1288# 0.308854f
C346 source.n104 a_n2094_n1288# 0.823249f
C347 plus.n0 a_n2094_n1288# 0.02774f
C348 plus.t2 a_n2094_n1288# 0.03265f
C349 plus.t8 a_n2094_n1288# 0.03265f
C350 plus.t15 a_n2094_n1288# 0.03265f
C351 plus.n1 a_n2094_n1288# 0.025654f
C352 plus.n2 a_n2094_n1288# 0.02774f
C353 plus.t21 a_n2094_n1288# 0.03265f
C354 plus.t5 a_n2094_n1288# 0.03265f
C355 plus.t10 a_n2094_n1288# 0.03265f
C356 plus.n3 a_n2094_n1288# 0.025654f
C357 plus.n4 a_n2094_n1288# 0.02774f
C358 plus.t16 a_n2094_n1288# 0.03265f
C359 plus.t17 a_n2094_n1288# 0.03265f
C360 plus.t22 a_n2094_n1288# 0.03265f
C361 plus.n5 a_n2094_n1288# 0.025654f
C362 plus.t11 a_n2094_n1288# 0.036304f
C363 plus.n6 a_n2094_n1288# 0.033726f
C364 plus.t6 a_n2094_n1288# 0.03265f
C365 plus.n7 a_n2094_n1288# 0.025654f
C366 plus.n8 a_n2094_n1288# 0.009715f
C367 plus.n9 a_n2094_n1288# 0.0645f
C368 plus.n10 a_n2094_n1288# 0.02774f
C369 plus.n11 a_n2094_n1288# 0.009715f
C370 plus.n12 a_n2094_n1288# 0.025654f
C371 plus.n13 a_n2094_n1288# 0.009715f
C372 plus.n14 a_n2094_n1288# 0.025654f
C373 plus.n15 a_n2094_n1288# 0.009715f
C374 plus.n16 a_n2094_n1288# 0.02774f
C375 plus.n17 a_n2094_n1288# 0.02774f
C376 plus.n18 a_n2094_n1288# 0.009715f
C377 plus.n19 a_n2094_n1288# 0.025654f
C378 plus.n20 a_n2094_n1288# 0.009715f
C379 plus.n21 a_n2094_n1288# 0.025654f
C380 plus.n22 a_n2094_n1288# 0.009715f
C381 plus.n23 a_n2094_n1288# 0.02774f
C382 plus.n24 a_n2094_n1288# 0.02774f
C383 plus.n25 a_n2094_n1288# 0.009715f
C384 plus.n26 a_n2094_n1288# 0.025654f
C385 plus.n27 a_n2094_n1288# 0.009715f
C386 plus.n28 a_n2094_n1288# 0.025654f
C387 plus.t19 a_n2094_n1288# 0.036304f
C388 plus.n29 a_n2094_n1288# 0.033682f
C389 plus.n30 a_n2094_n1288# 0.197558f
C390 plus.n31 a_n2094_n1288# 0.02774f
C391 plus.t14 a_n2094_n1288# 0.036304f
C392 plus.t9 a_n2094_n1288# 0.03265f
C393 plus.t4 a_n2094_n1288# 0.03265f
C394 plus.t23 a_n2094_n1288# 0.03265f
C395 plus.n32 a_n2094_n1288# 0.025654f
C396 plus.n33 a_n2094_n1288# 0.02774f
C397 plus.t12 a_n2094_n1288# 0.03265f
C398 plus.t0 a_n2094_n1288# 0.03265f
C399 plus.t18 a_n2094_n1288# 0.03265f
C400 plus.n34 a_n2094_n1288# 0.025654f
C401 plus.n35 a_n2094_n1288# 0.02774f
C402 plus.t7 a_n2094_n1288# 0.03265f
C403 plus.t1 a_n2094_n1288# 0.03265f
C404 plus.t13 a_n2094_n1288# 0.03265f
C405 plus.n36 a_n2094_n1288# 0.025654f
C406 plus.t20 a_n2094_n1288# 0.036304f
C407 plus.n37 a_n2094_n1288# 0.033726f
C408 plus.t3 a_n2094_n1288# 0.03265f
C409 plus.n38 a_n2094_n1288# 0.025654f
C410 plus.n39 a_n2094_n1288# 0.009715f
C411 plus.n40 a_n2094_n1288# 0.0645f
C412 plus.n41 a_n2094_n1288# 0.02774f
C413 plus.n42 a_n2094_n1288# 0.009715f
C414 plus.n43 a_n2094_n1288# 0.025654f
C415 plus.n44 a_n2094_n1288# 0.009715f
C416 plus.n45 a_n2094_n1288# 0.025654f
C417 plus.n46 a_n2094_n1288# 0.009715f
C418 plus.n47 a_n2094_n1288# 0.02774f
C419 plus.n48 a_n2094_n1288# 0.02774f
C420 plus.n49 a_n2094_n1288# 0.009715f
C421 plus.n50 a_n2094_n1288# 0.025654f
C422 plus.n51 a_n2094_n1288# 0.009715f
C423 plus.n52 a_n2094_n1288# 0.025654f
C424 plus.n53 a_n2094_n1288# 0.009715f
C425 plus.n54 a_n2094_n1288# 0.02774f
C426 plus.n55 a_n2094_n1288# 0.02774f
C427 plus.n56 a_n2094_n1288# 0.009715f
C428 plus.n57 a_n2094_n1288# 0.025654f
C429 plus.n58 a_n2094_n1288# 0.009715f
C430 plus.n59 a_n2094_n1288# 0.025654f
C431 plus.n60 a_n2094_n1288# 0.033682f
C432 plus.n61 a_n2094_n1288# 0.666546f
.ends

