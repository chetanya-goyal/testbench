* NGSPICE file created from diffpair181.ext - technology: sky130A

.subckt diffpair181 minus drain_right drain_left source plus
X0 drain_right.t3 minus.t0 source.t5 a_n1064_n1492# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X1 drain_right.t2 minus.t1 source.t4 a_n1064_n1492# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X2 a_n1064_n1492# a_n1064_n1492# a_n1064_n1492# a_n1064_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.25
X3 a_n1064_n1492# a_n1064_n1492# a_n1064_n1492# a_n1064_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X4 drain_left.t3 plus.t0 source.t3 a_n1064_n1492# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X5 source.t6 minus.t2 drain_right.t1 a_n1064_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X6 a_n1064_n1492# a_n1064_n1492# a_n1064_n1492# a_n1064_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X7 a_n1064_n1492# a_n1064_n1492# a_n1064_n1492# a_n1064_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X8 source.t0 plus.t1 drain_left.t2 a_n1064_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X9 source.t1 plus.t2 drain_left.t1 a_n1064_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X10 drain_left.t0 plus.t3 source.t2 a_n1064_n1492# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X11 source.t7 minus.t3 drain_right.t0 a_n1064_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
R0 minus.n0 minus.t2 456.878
R1 minus.n0 minus.t0 456.878
R2 minus.n1 minus.t1 456.878
R3 minus.n1 minus.t3 456.878
R4 minus.n2 minus.n0 187.619
R5 minus.n2 minus.n1 167.77
R6 minus minus.n2 0.188
R7 source.n0 source.t3 69.6943
R8 source.n1 source.t0 69.6943
R9 source.n2 source.t5 69.6943
R10 source.n3 source.t6 69.6943
R11 source.n7 source.t4 69.6942
R12 source.n6 source.t7 69.6942
R13 source.n5 source.t2 69.6942
R14 source.n4 source.t1 69.6942
R15 source.n4 source.n3 14.9847
R16 source.n8 source.n0 9.47176
R17 source.n8 source.n7 5.51343
R18 source.n3 source.n2 0.5005
R19 source.n1 source.n0 0.5005
R20 source.n5 source.n4 0.5005
R21 source.n7 source.n6 0.5005
R22 source.n2 source.n1 0.470328
R23 source.n6 source.n5 0.470328
R24 source source.n8 0.188
R25 drain_right drain_right.n0 100.784
R26 drain_right drain_right.n1 85.9258
R27 drain_right.n0 drain_right.t0 6.6005
R28 drain_right.n0 drain_right.t2 6.6005
R29 drain_right.n1 drain_right.t1 6.6005
R30 drain_right.n1 drain_right.t3 6.6005
R31 plus.n0 plus.t1 456.878
R32 plus.n0 plus.t0 456.878
R33 plus.n1 plus.t3 456.878
R34 plus.n1 plus.t2 456.878
R35 plus plus.n1 184.909
R36 plus plus.n0 170.006
R37 drain_left drain_left.n0 101.337
R38 drain_left drain_left.n1 85.9258
R39 drain_left.n0 drain_left.t1 6.6005
R40 drain_left.n0 drain_left.t0 6.6005
R41 drain_left.n1 drain_left.t2 6.6005
R42 drain_left.n1 drain_left.t3 6.6005
C0 minus drain_right 0.684987f
C1 source minus 0.604552f
C2 plus drain_left 0.782838f
C3 plus drain_right 0.257181f
C4 plus source 0.618551f
C5 plus minus 2.81396f
C6 drain_left drain_right 0.467167f
C7 drain_left source 3.54359f
C8 drain_left minus 0.176155f
C9 source drain_right 3.54184f
C10 drain_right a_n1064_n1492# 3.90363f
C11 drain_left a_n1064_n1492# 4.03087f
C12 source a_n1064_n1492# 3.186625f
C13 minus a_n1064_n1492# 3.357801f
C14 plus a_n1064_n1492# 5.24388f
C15 drain_left.t1 a_n1064_n1492# 0.058215f
C16 drain_left.t0 a_n1064_n1492# 0.058215f
C17 drain_left.n0 a_n1064_n1492# 0.561277f
C18 drain_left.t2 a_n1064_n1492# 0.058215f
C19 drain_left.t3 a_n1064_n1492# 0.058215f
C20 drain_left.n1 a_n1064_n1492# 0.454808f
C21 plus.t1 a_n1064_n1492# 0.096809f
C22 plus.t0 a_n1064_n1492# 0.096809f
C23 plus.n0 a_n1064_n1492# 0.134785f
C24 plus.t2 a_n1064_n1492# 0.096809f
C25 plus.t3 a_n1064_n1492# 0.096809f
C26 plus.n1 a_n1064_n1492# 0.224765f
C27 drain_right.t0 a_n1064_n1492# 0.059858f
C28 drain_right.t2 a_n1064_n1492# 0.059858f
C29 drain_right.n0 a_n1064_n1492# 0.563623f
C30 drain_right.t1 a_n1064_n1492# 0.059858f
C31 drain_right.t3 a_n1064_n1492# 0.059858f
C32 drain_right.n1 a_n1064_n1492# 0.467643f
C33 source.t3 a_n1064_n1492# 0.379888f
C34 source.n0 a_n1064_n1492# 0.514404f
C35 source.t0 a_n1064_n1492# 0.379888f
C36 source.n1 a_n1064_n1492# 0.263365f
C37 source.t5 a_n1064_n1492# 0.379888f
C38 source.n2 a_n1064_n1492# 0.263365f
C39 source.t6 a_n1064_n1492# 0.379888f
C40 source.n3 a_n1064_n1492# 0.715306f
C41 source.t1 a_n1064_n1492# 0.379886f
C42 source.n4 a_n1064_n1492# 0.715308f
C43 source.t2 a_n1064_n1492# 0.379886f
C44 source.n5 a_n1064_n1492# 0.263367f
C45 source.t7 a_n1064_n1492# 0.379886f
C46 source.n6 a_n1064_n1492# 0.263367f
C47 source.t4 a_n1064_n1492# 0.379886f
C48 source.n7 a_n1064_n1492# 0.370156f
C49 source.n8 a_n1064_n1492# 0.55978f
C50 minus.t2 a_n1064_n1492# 0.093947f
C51 minus.t0 a_n1064_n1492# 0.093947f
C52 minus.n0 a_n1064_n1492# 0.234289f
C53 minus.t3 a_n1064_n1492# 0.093947f
C54 minus.t1 a_n1064_n1492# 0.093947f
C55 minus.n1 a_n1064_n1492# 0.125406f
C56 minus.n2 a_n1064_n1492# 2.03764f
.ends

