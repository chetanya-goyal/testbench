* NGSPICE file created from diffpair119.ext - technology: sky130A

.subckt diffpair119 minus drain_right drain_left source plus
X0 drain_right.t23 minus.t0 source.t27 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X1 source.t12 plus.t0 drain_left.t23 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X2 source.t40 minus.t1 drain_right.t22 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X3 source.t5 plus.t1 drain_left.t22 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X4 drain_left.t21 plus.t2 source.t14 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X5 source.t38 minus.t2 drain_right.t21 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X6 a_n2354_n1288# a_n2354_n1288# a_n2354_n1288# a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.3
X7 drain_right.t20 minus.t3 source.t44 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X8 drain_right.t19 minus.t4 source.t45 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X9 source.t46 minus.t5 drain_right.t18 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X10 drain_right.t17 minus.t6 source.t37 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X11 drain_left.t20 plus.t3 source.t6 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X12 source.t19 plus.t4 drain_left.t19 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X13 drain_right.t16 minus.t7 source.t47 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X14 drain_left.t18 plus.t5 source.t23 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X15 source.t35 minus.t8 drain_right.t15 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X16 source.t13 plus.t6 drain_left.t17 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X17 a_n2354_n1288# a_n2354_n1288# a_n2354_n1288# a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X18 drain_right.t14 minus.t9 source.t43 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X19 source.t25 minus.t10 drain_right.t13 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X20 source.t31 minus.t11 drain_right.t12 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X21 drain_left.t16 plus.t7 source.t0 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X22 source.t4 plus.t8 drain_left.t15 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X23 drain_left.t14 plus.t9 source.t9 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X24 drain_right.t11 minus.t12 source.t26 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X25 source.t39 minus.t13 drain_right.t10 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X26 source.t16 plus.t10 drain_left.t13 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X27 source.t21 plus.t11 drain_left.t12 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X28 source.t30 minus.t14 drain_right.t9 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X29 source.t1 plus.t12 drain_left.t11 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X30 source.t8 plus.t13 drain_left.t10 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X31 source.t41 minus.t15 drain_right.t8 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X32 drain_right.t7 minus.t16 source.t42 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X33 drain_left.t9 plus.t14 source.t10 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X34 drain_right.t6 minus.t17 source.t28 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X35 drain_right.t5 minus.t18 source.t33 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X36 drain_left.t8 plus.t15 source.t15 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X37 drain_left.t7 plus.t16 source.t20 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X38 source.t11 plus.t17 drain_left.t6 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X39 source.t34 minus.t19 drain_right.t4 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X40 source.t18 plus.t18 drain_left.t5 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X41 drain_left.t4 plus.t19 source.t17 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X42 drain_right.t3 minus.t20 source.t29 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X43 drain_right.t2 minus.t21 source.t32 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X44 a_n2354_n1288# a_n2354_n1288# a_n2354_n1288# a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X45 a_n2354_n1288# a_n2354_n1288# a_n2354_n1288# a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X46 source.t36 minus.t22 drain_right.t1 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X47 source.t24 minus.t23 drain_right.t0 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X48 drain_left.t3 plus.t20 source.t22 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X49 drain_left.t2 plus.t21 source.t3 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X50 source.t7 plus.t22 drain_left.t1 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X51 drain_left.t0 plus.t23 source.t2 a_n2354_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
R0 minus.n35 minus.t5 296.503
R1 minus.n9 minus.t16 296.503
R2 minus.n72 minus.t0 296.503
R3 minus.n46 minus.t1 296.503
R4 minus.n34 minus.t21 265.101
R5 minus.n1 minus.t10 265.101
R6 minus.n28 minus.t4 265.101
R7 minus.n26 minus.t23 265.101
R8 minus.n3 minus.t9 265.101
R9 minus.n20 minus.t2 265.101
R10 minus.n5 minus.t20 265.101
R11 minus.n15 minus.t14 265.101
R12 minus.n13 minus.t3 265.101
R13 minus.n8 minus.t22 265.101
R14 minus.n71 minus.t11 265.101
R15 minus.n38 minus.t12 265.101
R16 minus.n65 minus.t15 265.101
R17 minus.n63 minus.t7 265.101
R18 minus.n40 minus.t8 265.101
R19 minus.n57 minus.t17 265.101
R20 minus.n42 minus.t19 265.101
R21 minus.n52 minus.t6 265.101
R22 minus.n50 minus.t13 265.101
R23 minus.n45 minus.t18 265.101
R24 minus.n10 minus.n9 161.489
R25 minus.n47 minus.n46 161.489
R26 minus.n36 minus.n35 161.3
R27 minus.n33 minus.n0 161.3
R28 minus.n32 minus.n31 161.3
R29 minus.n30 minus.n29 161.3
R30 minus.n27 minus.n2 161.3
R31 minus.n25 minus.n24 161.3
R32 minus.n23 minus.n22 161.3
R33 minus.n21 minus.n4 161.3
R34 minus.n19 minus.n18 161.3
R35 minus.n17 minus.n16 161.3
R36 minus.n14 minus.n6 161.3
R37 minus.n12 minus.n11 161.3
R38 minus.n10 minus.n7 161.3
R39 minus.n73 minus.n72 161.3
R40 minus.n70 minus.n37 161.3
R41 minus.n69 minus.n68 161.3
R42 minus.n67 minus.n66 161.3
R43 minus.n64 minus.n39 161.3
R44 minus.n62 minus.n61 161.3
R45 minus.n60 minus.n59 161.3
R46 minus.n58 minus.n41 161.3
R47 minus.n56 minus.n55 161.3
R48 minus.n54 minus.n53 161.3
R49 minus.n51 minus.n43 161.3
R50 minus.n49 minus.n48 161.3
R51 minus.n47 minus.n44 161.3
R52 minus.n33 minus.n32 73.0308
R53 minus.n22 minus.n21 73.0308
R54 minus.n12 minus.n7 73.0308
R55 minus.n49 minus.n44 73.0308
R56 minus.n59 minus.n58 73.0308
R57 minus.n70 minus.n69 73.0308
R58 minus.n29 minus.n1 66.4581
R59 minus.n14 minus.n13 66.4581
R60 minus.n51 minus.n50 66.4581
R61 minus.n66 minus.n38 66.4581
R62 minus.n25 minus.n3 63.5369
R63 minus.n20 minus.n19 63.5369
R64 minus.n57 minus.n56 63.5369
R65 minus.n62 minus.n40 63.5369
R66 minus.n35 minus.n34 60.6157
R67 minus.n9 minus.n8 60.6157
R68 minus.n46 minus.n45 60.6157
R69 minus.n72 minus.n71 60.6157
R70 minus.n28 minus.n27 47.4702
R71 minus.n16 minus.n15 47.4702
R72 minus.n53 minus.n52 47.4702
R73 minus.n65 minus.n64 47.4702
R74 minus.n27 minus.n26 44.549
R75 minus.n16 minus.n5 44.549
R76 minus.n53 minus.n42 44.549
R77 minus.n64 minus.n63 44.549
R78 minus.n74 minus.n36 30.4323
R79 minus.n26 minus.n25 28.4823
R80 minus.n19 minus.n5 28.4823
R81 minus.n56 minus.n42 28.4823
R82 minus.n63 minus.n62 28.4823
R83 minus.n29 minus.n28 25.5611
R84 minus.n15 minus.n14 25.5611
R85 minus.n52 minus.n51 25.5611
R86 minus.n66 minus.n65 25.5611
R87 minus.n34 minus.n33 12.4157
R88 minus.n8 minus.n7 12.4157
R89 minus.n45 minus.n44 12.4157
R90 minus.n71 minus.n70 12.4157
R91 minus.n22 minus.n3 9.49444
R92 minus.n21 minus.n20 9.49444
R93 minus.n58 minus.n57 9.49444
R94 minus.n59 minus.n40 9.49444
R95 minus.n32 minus.n1 6.57323
R96 minus.n13 minus.n12 6.57323
R97 minus.n50 minus.n49 6.57323
R98 minus.n69 minus.n38 6.57323
R99 minus.n74 minus.n73 6.4702
R100 minus.n36 minus.n0 0.189894
R101 minus.n31 minus.n0 0.189894
R102 minus.n31 minus.n30 0.189894
R103 minus.n30 minus.n2 0.189894
R104 minus.n24 minus.n2 0.189894
R105 minus.n24 minus.n23 0.189894
R106 minus.n23 minus.n4 0.189894
R107 minus.n18 minus.n4 0.189894
R108 minus.n18 minus.n17 0.189894
R109 minus.n17 minus.n6 0.189894
R110 minus.n11 minus.n6 0.189894
R111 minus.n11 minus.n10 0.189894
R112 minus.n48 minus.n47 0.189894
R113 minus.n48 minus.n43 0.189894
R114 minus.n54 minus.n43 0.189894
R115 minus.n55 minus.n54 0.189894
R116 minus.n55 minus.n41 0.189894
R117 minus.n60 minus.n41 0.189894
R118 minus.n61 minus.n60 0.189894
R119 minus.n61 minus.n39 0.189894
R120 minus.n67 minus.n39 0.189894
R121 minus.n68 minus.n67 0.189894
R122 minus.n68 minus.n37 0.189894
R123 minus.n73 minus.n37 0.189894
R124 minus minus.n74 0.188
R125 source.n98 source.n96 289.615
R126 source.n80 source.n78 289.615
R127 source.n72 source.n70 289.615
R128 source.n54 source.n52 289.615
R129 source.n2 source.n0 289.615
R130 source.n20 source.n18 289.615
R131 source.n28 source.n26 289.615
R132 source.n46 source.n44 289.615
R133 source.n99 source.n98 185
R134 source.n81 source.n80 185
R135 source.n73 source.n72 185
R136 source.n55 source.n54 185
R137 source.n3 source.n2 185
R138 source.n21 source.n20 185
R139 source.n29 source.n28 185
R140 source.n47 source.n46 185
R141 source.t27 source.n97 167.117
R142 source.t40 source.n79 167.117
R143 source.t22 source.n71 167.117
R144 source.t21 source.n53 167.117
R145 source.t23 source.n1 167.117
R146 source.t19 source.n19 167.117
R147 source.t42 source.n27 167.117
R148 source.t46 source.n45 167.117
R149 source.n9 source.n8 84.1169
R150 source.n11 source.n10 84.1169
R151 source.n13 source.n12 84.1169
R152 source.n15 source.n14 84.1169
R153 source.n17 source.n16 84.1169
R154 source.n35 source.n34 84.1169
R155 source.n37 source.n36 84.1169
R156 source.n39 source.n38 84.1169
R157 source.n41 source.n40 84.1169
R158 source.n43 source.n42 84.1169
R159 source.n95 source.n94 84.1168
R160 source.n93 source.n92 84.1168
R161 source.n91 source.n90 84.1168
R162 source.n89 source.n88 84.1168
R163 source.n87 source.n86 84.1168
R164 source.n69 source.n68 84.1168
R165 source.n67 source.n66 84.1168
R166 source.n65 source.n64 84.1168
R167 source.n63 source.n62 84.1168
R168 source.n61 source.n60 84.1168
R169 source.n98 source.t27 52.3082
R170 source.n80 source.t40 52.3082
R171 source.n72 source.t22 52.3082
R172 source.n54 source.t21 52.3082
R173 source.n2 source.t23 52.3082
R174 source.n20 source.t19 52.3082
R175 source.n28 source.t42 52.3082
R176 source.n46 source.t46 52.3082
R177 source.n103 source.n102 31.4096
R178 source.n85 source.n84 31.4096
R179 source.n77 source.n76 31.4096
R180 source.n59 source.n58 31.4096
R181 source.n7 source.n6 31.4096
R182 source.n25 source.n24 31.4096
R183 source.n33 source.n32 31.4096
R184 source.n51 source.n50 31.4096
R185 source.n59 source.n51 14.2551
R186 source.n94 source.t26 9.9005
R187 source.n94 source.t31 9.9005
R188 source.n92 source.t47 9.9005
R189 source.n92 source.t41 9.9005
R190 source.n90 source.t28 9.9005
R191 source.n90 source.t35 9.9005
R192 source.n88 source.t37 9.9005
R193 source.n88 source.t34 9.9005
R194 source.n86 source.t33 9.9005
R195 source.n86 source.t39 9.9005
R196 source.n68 source.t0 9.9005
R197 source.n68 source.t16 9.9005
R198 source.n66 source.t15 9.9005
R199 source.n66 source.t5 9.9005
R200 source.n64 source.t6 9.9005
R201 source.n64 source.t1 9.9005
R202 source.n62 source.t20 9.9005
R203 source.n62 source.t18 9.9005
R204 source.n60 source.t3 9.9005
R205 source.n60 source.t13 9.9005
R206 source.n8 source.t17 9.9005
R207 source.n8 source.t12 9.9005
R208 source.n10 source.t14 9.9005
R209 source.n10 source.t8 9.9005
R210 source.n12 source.t10 9.9005
R211 source.n12 source.t7 9.9005
R212 source.n14 source.t2 9.9005
R213 source.n14 source.t4 9.9005
R214 source.n16 source.t9 9.9005
R215 source.n16 source.t11 9.9005
R216 source.n34 source.t44 9.9005
R217 source.n34 source.t36 9.9005
R218 source.n36 source.t29 9.9005
R219 source.n36 source.t30 9.9005
R220 source.n38 source.t43 9.9005
R221 source.n38 source.t38 9.9005
R222 source.n40 source.t45 9.9005
R223 source.n40 source.t24 9.9005
R224 source.n42 source.t32 9.9005
R225 source.n42 source.t25 9.9005
R226 source.n99 source.n97 9.71174
R227 source.n81 source.n79 9.71174
R228 source.n73 source.n71 9.71174
R229 source.n55 source.n53 9.71174
R230 source.n3 source.n1 9.71174
R231 source.n21 source.n19 9.71174
R232 source.n29 source.n27 9.71174
R233 source.n47 source.n45 9.71174
R234 source.n102 source.n101 9.45567
R235 source.n84 source.n83 9.45567
R236 source.n76 source.n75 9.45567
R237 source.n58 source.n57 9.45567
R238 source.n6 source.n5 9.45567
R239 source.n24 source.n23 9.45567
R240 source.n32 source.n31 9.45567
R241 source.n50 source.n49 9.45567
R242 source.n101 source.n100 9.3005
R243 source.n83 source.n82 9.3005
R244 source.n75 source.n74 9.3005
R245 source.n57 source.n56 9.3005
R246 source.n5 source.n4 9.3005
R247 source.n23 source.n22 9.3005
R248 source.n31 source.n30 9.3005
R249 source.n49 source.n48 9.3005
R250 source.n104 source.n7 8.72059
R251 source.n102 source.n96 8.14595
R252 source.n84 source.n78 8.14595
R253 source.n76 source.n70 8.14595
R254 source.n58 source.n52 8.14595
R255 source.n6 source.n0 8.14595
R256 source.n24 source.n18 8.14595
R257 source.n32 source.n26 8.14595
R258 source.n50 source.n44 8.14595
R259 source.n100 source.n99 7.3702
R260 source.n82 source.n81 7.3702
R261 source.n74 source.n73 7.3702
R262 source.n56 source.n55 7.3702
R263 source.n4 source.n3 7.3702
R264 source.n22 source.n21 7.3702
R265 source.n30 source.n29 7.3702
R266 source.n48 source.n47 7.3702
R267 source.n100 source.n96 5.81868
R268 source.n82 source.n78 5.81868
R269 source.n74 source.n70 5.81868
R270 source.n56 source.n52 5.81868
R271 source.n4 source.n0 5.81868
R272 source.n22 source.n18 5.81868
R273 source.n30 source.n26 5.81868
R274 source.n48 source.n44 5.81868
R275 source.n104 source.n103 5.53498
R276 source.n101 source.n97 3.44771
R277 source.n83 source.n79 3.44771
R278 source.n75 source.n71 3.44771
R279 source.n57 source.n53 3.44771
R280 source.n5 source.n1 3.44771
R281 source.n23 source.n19 3.44771
R282 source.n31 source.n27 3.44771
R283 source.n49 source.n45 3.44771
R284 source.n51 source.n43 0.543603
R285 source.n43 source.n41 0.543603
R286 source.n41 source.n39 0.543603
R287 source.n39 source.n37 0.543603
R288 source.n37 source.n35 0.543603
R289 source.n35 source.n33 0.543603
R290 source.n25 source.n17 0.543603
R291 source.n17 source.n15 0.543603
R292 source.n15 source.n13 0.543603
R293 source.n13 source.n11 0.543603
R294 source.n11 source.n9 0.543603
R295 source.n9 source.n7 0.543603
R296 source.n61 source.n59 0.543603
R297 source.n63 source.n61 0.543603
R298 source.n65 source.n63 0.543603
R299 source.n67 source.n65 0.543603
R300 source.n69 source.n67 0.543603
R301 source.n77 source.n69 0.543603
R302 source.n87 source.n85 0.543603
R303 source.n89 source.n87 0.543603
R304 source.n91 source.n89 0.543603
R305 source.n93 source.n91 0.543603
R306 source.n95 source.n93 0.543603
R307 source.n103 source.n95 0.543603
R308 source.n33 source.n25 0.470328
R309 source.n85 source.n77 0.470328
R310 source source.n104 0.188
R311 drain_right.n13 drain_right.n11 101.338
R312 drain_right.n7 drain_right.n5 101.338
R313 drain_right.n2 drain_right.n0 101.338
R314 drain_right.n13 drain_right.n12 100.796
R315 drain_right.n15 drain_right.n14 100.796
R316 drain_right.n17 drain_right.n16 100.796
R317 drain_right.n19 drain_right.n18 100.796
R318 drain_right.n21 drain_right.n20 100.796
R319 drain_right.n7 drain_right.n6 100.796
R320 drain_right.n9 drain_right.n8 100.796
R321 drain_right.n4 drain_right.n3 100.796
R322 drain_right.n2 drain_right.n1 100.796
R323 drain_right drain_right.n10 24.3976
R324 drain_right.n5 drain_right.t12 9.9005
R325 drain_right.n5 drain_right.t23 9.9005
R326 drain_right.n6 drain_right.t8 9.9005
R327 drain_right.n6 drain_right.t11 9.9005
R328 drain_right.n8 drain_right.t15 9.9005
R329 drain_right.n8 drain_right.t16 9.9005
R330 drain_right.n3 drain_right.t4 9.9005
R331 drain_right.n3 drain_right.t6 9.9005
R332 drain_right.n1 drain_right.t10 9.9005
R333 drain_right.n1 drain_right.t17 9.9005
R334 drain_right.n0 drain_right.t22 9.9005
R335 drain_right.n0 drain_right.t5 9.9005
R336 drain_right.n11 drain_right.t1 9.9005
R337 drain_right.n11 drain_right.t7 9.9005
R338 drain_right.n12 drain_right.t9 9.9005
R339 drain_right.n12 drain_right.t20 9.9005
R340 drain_right.n14 drain_right.t21 9.9005
R341 drain_right.n14 drain_right.t3 9.9005
R342 drain_right.n16 drain_right.t0 9.9005
R343 drain_right.n16 drain_right.t14 9.9005
R344 drain_right.n18 drain_right.t13 9.9005
R345 drain_right.n18 drain_right.t19 9.9005
R346 drain_right.n20 drain_right.t18 9.9005
R347 drain_right.n20 drain_right.t2 9.9005
R348 drain_right drain_right.n21 6.19632
R349 drain_right.n9 drain_right.n7 0.543603
R350 drain_right.n4 drain_right.n2 0.543603
R351 drain_right.n21 drain_right.n19 0.543603
R352 drain_right.n19 drain_right.n17 0.543603
R353 drain_right.n17 drain_right.n15 0.543603
R354 drain_right.n15 drain_right.n13 0.543603
R355 drain_right.n10 drain_right.n9 0.216706
R356 drain_right.n10 drain_right.n4 0.216706
R357 plus.n9 plus.t4 296.503
R358 plus.n35 plus.t5 296.503
R359 plus.n46 plus.t20 296.503
R360 plus.n72 plus.t11 296.503
R361 plus.n8 plus.t9 265.101
R362 plus.n13 plus.t17 265.101
R363 plus.n15 plus.t23 265.101
R364 plus.n5 plus.t8 265.101
R365 plus.n20 plus.t14 265.101
R366 plus.n3 plus.t22 265.101
R367 plus.n26 plus.t2 265.101
R368 plus.n28 plus.t13 265.101
R369 plus.n1 plus.t19 265.101
R370 plus.n34 plus.t0 265.101
R371 plus.n45 plus.t10 265.101
R372 plus.n50 plus.t7 265.101
R373 plus.n52 plus.t1 265.101
R374 plus.n42 plus.t15 265.101
R375 plus.n57 plus.t12 265.101
R376 plus.n40 plus.t3 265.101
R377 plus.n63 plus.t18 265.101
R378 plus.n65 plus.t16 265.101
R379 plus.n38 plus.t6 265.101
R380 plus.n71 plus.t21 265.101
R381 plus.n10 plus.n9 161.489
R382 plus.n47 plus.n46 161.489
R383 plus.n10 plus.n7 161.3
R384 plus.n12 plus.n11 161.3
R385 plus.n14 plus.n6 161.3
R386 plus.n17 plus.n16 161.3
R387 plus.n19 plus.n18 161.3
R388 plus.n21 plus.n4 161.3
R389 plus.n23 plus.n22 161.3
R390 plus.n25 plus.n24 161.3
R391 plus.n27 plus.n2 161.3
R392 plus.n30 plus.n29 161.3
R393 plus.n32 plus.n31 161.3
R394 plus.n33 plus.n0 161.3
R395 plus.n36 plus.n35 161.3
R396 plus.n47 plus.n44 161.3
R397 plus.n49 plus.n48 161.3
R398 plus.n51 plus.n43 161.3
R399 plus.n54 plus.n53 161.3
R400 plus.n56 plus.n55 161.3
R401 plus.n58 plus.n41 161.3
R402 plus.n60 plus.n59 161.3
R403 plus.n62 plus.n61 161.3
R404 plus.n64 plus.n39 161.3
R405 plus.n67 plus.n66 161.3
R406 plus.n69 plus.n68 161.3
R407 plus.n70 plus.n37 161.3
R408 plus.n73 plus.n72 161.3
R409 plus.n12 plus.n7 73.0308
R410 plus.n22 plus.n21 73.0308
R411 plus.n33 plus.n32 73.0308
R412 plus.n70 plus.n69 73.0308
R413 plus.n59 plus.n58 73.0308
R414 plus.n49 plus.n44 73.0308
R415 plus.n14 plus.n13 66.4581
R416 plus.n29 plus.n1 66.4581
R417 plus.n66 plus.n38 66.4581
R418 plus.n51 plus.n50 66.4581
R419 plus.n20 plus.n19 63.5369
R420 plus.n25 plus.n3 63.5369
R421 plus.n62 plus.n40 63.5369
R422 plus.n57 plus.n56 63.5369
R423 plus.n9 plus.n8 60.6157
R424 plus.n35 plus.n34 60.6157
R425 plus.n72 plus.n71 60.6157
R426 plus.n46 plus.n45 60.6157
R427 plus.n16 plus.n15 47.4702
R428 plus.n28 plus.n27 47.4702
R429 plus.n65 plus.n64 47.4702
R430 plus.n53 plus.n52 47.4702
R431 plus.n16 plus.n5 44.549
R432 plus.n27 plus.n26 44.549
R433 plus.n64 plus.n63 44.549
R434 plus.n53 plus.n42 44.549
R435 plus.n19 plus.n5 28.4823
R436 plus.n26 plus.n25 28.4823
R437 plus.n63 plus.n62 28.4823
R438 plus.n56 plus.n42 28.4823
R439 plus plus.n73 28.1013
R440 plus.n15 plus.n14 25.5611
R441 plus.n29 plus.n28 25.5611
R442 plus.n66 plus.n65 25.5611
R443 plus.n52 plus.n51 25.5611
R444 plus.n8 plus.n7 12.4157
R445 plus.n34 plus.n33 12.4157
R446 plus.n71 plus.n70 12.4157
R447 plus.n45 plus.n44 12.4157
R448 plus.n21 plus.n20 9.49444
R449 plus.n22 plus.n3 9.49444
R450 plus.n59 plus.n40 9.49444
R451 plus.n58 plus.n57 9.49444
R452 plus plus.n36 8.32626
R453 plus.n13 plus.n12 6.57323
R454 plus.n32 plus.n1 6.57323
R455 plus.n69 plus.n38 6.57323
R456 plus.n50 plus.n49 6.57323
R457 plus.n11 plus.n10 0.189894
R458 plus.n11 plus.n6 0.189894
R459 plus.n17 plus.n6 0.189894
R460 plus.n18 plus.n17 0.189894
R461 plus.n18 plus.n4 0.189894
R462 plus.n23 plus.n4 0.189894
R463 plus.n24 plus.n23 0.189894
R464 plus.n24 plus.n2 0.189894
R465 plus.n30 plus.n2 0.189894
R466 plus.n31 plus.n30 0.189894
R467 plus.n31 plus.n0 0.189894
R468 plus.n36 plus.n0 0.189894
R469 plus.n73 plus.n37 0.189894
R470 plus.n68 plus.n37 0.189894
R471 plus.n68 plus.n67 0.189894
R472 plus.n67 plus.n39 0.189894
R473 plus.n61 plus.n39 0.189894
R474 plus.n61 plus.n60 0.189894
R475 plus.n60 plus.n41 0.189894
R476 plus.n55 plus.n41 0.189894
R477 plus.n55 plus.n54 0.189894
R478 plus.n54 plus.n43 0.189894
R479 plus.n48 plus.n43 0.189894
R480 plus.n48 plus.n47 0.189894
R481 drain_left.n13 drain_left.n11 101.338
R482 drain_left.n7 drain_left.n5 101.338
R483 drain_left.n2 drain_left.n0 101.338
R484 drain_left.n21 drain_left.n20 100.796
R485 drain_left.n19 drain_left.n18 100.796
R486 drain_left.n17 drain_left.n16 100.796
R487 drain_left.n15 drain_left.n14 100.796
R488 drain_left.n13 drain_left.n12 100.796
R489 drain_left.n7 drain_left.n6 100.796
R490 drain_left.n9 drain_left.n8 100.796
R491 drain_left.n4 drain_left.n3 100.796
R492 drain_left.n2 drain_left.n1 100.796
R493 drain_left drain_left.n10 24.9508
R494 drain_left.n5 drain_left.t13 9.9005
R495 drain_left.n5 drain_left.t3 9.9005
R496 drain_left.n6 drain_left.t22 9.9005
R497 drain_left.n6 drain_left.t16 9.9005
R498 drain_left.n8 drain_left.t11 9.9005
R499 drain_left.n8 drain_left.t8 9.9005
R500 drain_left.n3 drain_left.t5 9.9005
R501 drain_left.n3 drain_left.t20 9.9005
R502 drain_left.n1 drain_left.t17 9.9005
R503 drain_left.n1 drain_left.t7 9.9005
R504 drain_left.n0 drain_left.t12 9.9005
R505 drain_left.n0 drain_left.t2 9.9005
R506 drain_left.n20 drain_left.t23 9.9005
R507 drain_left.n20 drain_left.t18 9.9005
R508 drain_left.n18 drain_left.t10 9.9005
R509 drain_left.n18 drain_left.t4 9.9005
R510 drain_left.n16 drain_left.t1 9.9005
R511 drain_left.n16 drain_left.t21 9.9005
R512 drain_left.n14 drain_left.t15 9.9005
R513 drain_left.n14 drain_left.t9 9.9005
R514 drain_left.n12 drain_left.t6 9.9005
R515 drain_left.n12 drain_left.t0 9.9005
R516 drain_left.n11 drain_left.t19 9.9005
R517 drain_left.n11 drain_left.t14 9.9005
R518 drain_left drain_left.n21 6.19632
R519 drain_left.n9 drain_left.n7 0.543603
R520 drain_left.n4 drain_left.n2 0.543603
R521 drain_left.n15 drain_left.n13 0.543603
R522 drain_left.n17 drain_left.n15 0.543603
R523 drain_left.n19 drain_left.n17 0.543603
R524 drain_left.n21 drain_left.n19 0.543603
R525 drain_left.n10 drain_left.n9 0.216706
R526 drain_left.n10 drain_left.n4 0.216706
C0 drain_right plus 0.39483f
C1 drain_right drain_left 1.26597f
C2 drain_right minus 1.96915f
C3 plus source 2.33714f
C4 drain_left source 10.5827f
C5 minus source 2.32317f
C6 drain_right source 10.5833f
C7 drain_left plus 2.20128f
C8 minus plus 4.25035f
C9 drain_left minus 0.178685f
C10 drain_right a_n2354_n1288# 4.72436f
C11 drain_left a_n2354_n1288# 5.38749f
C12 source a_n2354_n1288# 3.354887f
C13 minus a_n2354_n1288# 8.469373f
C14 plus a_n2354_n1288# 9.881619f
C15 drain_left.t12 a_n2354_n1288# 0.051412f
C16 drain_left.t2 a_n2354_n1288# 0.051412f
C17 drain_left.n0 a_n2354_n1288# 0.325f
C18 drain_left.t17 a_n2354_n1288# 0.051412f
C19 drain_left.t7 a_n2354_n1288# 0.051412f
C20 drain_left.n1 a_n2354_n1288# 0.322985f
C21 drain_left.n2 a_n2354_n1288# 0.736754f
C22 drain_left.t5 a_n2354_n1288# 0.051412f
C23 drain_left.t20 a_n2354_n1288# 0.051412f
C24 drain_left.n3 a_n2354_n1288# 0.322985f
C25 drain_left.n4 a_n2354_n1288# 0.332057f
C26 drain_left.t13 a_n2354_n1288# 0.051412f
C27 drain_left.t3 a_n2354_n1288# 0.051412f
C28 drain_left.n5 a_n2354_n1288# 0.325f
C29 drain_left.t22 a_n2354_n1288# 0.051412f
C30 drain_left.t16 a_n2354_n1288# 0.051412f
C31 drain_left.n6 a_n2354_n1288# 0.322985f
C32 drain_left.n7 a_n2354_n1288# 0.736755f
C33 drain_left.t11 a_n2354_n1288# 0.051412f
C34 drain_left.t8 a_n2354_n1288# 0.051412f
C35 drain_left.n8 a_n2354_n1288# 0.322985f
C36 drain_left.n9 a_n2354_n1288# 0.332057f
C37 drain_left.n10 a_n2354_n1288# 1.0912f
C38 drain_left.t19 a_n2354_n1288# 0.051412f
C39 drain_left.t14 a_n2354_n1288# 0.051412f
C40 drain_left.n11 a_n2354_n1288# 0.325002f
C41 drain_left.t6 a_n2354_n1288# 0.051412f
C42 drain_left.t0 a_n2354_n1288# 0.051412f
C43 drain_left.n12 a_n2354_n1288# 0.322987f
C44 drain_left.n13 a_n2354_n1288# 0.736752f
C45 drain_left.t15 a_n2354_n1288# 0.051412f
C46 drain_left.t9 a_n2354_n1288# 0.051412f
C47 drain_left.n14 a_n2354_n1288# 0.322987f
C48 drain_left.n15 a_n2354_n1288# 0.362832f
C49 drain_left.t1 a_n2354_n1288# 0.051412f
C50 drain_left.t21 a_n2354_n1288# 0.051412f
C51 drain_left.n16 a_n2354_n1288# 0.322987f
C52 drain_left.n17 a_n2354_n1288# 0.362832f
C53 drain_left.t10 a_n2354_n1288# 0.051412f
C54 drain_left.t4 a_n2354_n1288# 0.051412f
C55 drain_left.n18 a_n2354_n1288# 0.322987f
C56 drain_left.n19 a_n2354_n1288# 0.362832f
C57 drain_left.t23 a_n2354_n1288# 0.051412f
C58 drain_left.t18 a_n2354_n1288# 0.051412f
C59 drain_left.n20 a_n2354_n1288# 0.322987f
C60 drain_left.n21 a_n2354_n1288# 0.633597f
C61 plus.n0 a_n2354_n1288# 0.050595f
C62 plus.t0 a_n2354_n1288# 0.089328f
C63 plus.t19 a_n2354_n1288# 0.089328f
C64 plus.n1 a_n2354_n1288# 0.062388f
C65 plus.n2 a_n2354_n1288# 0.050595f
C66 plus.t13 a_n2354_n1288# 0.089328f
C67 plus.t2 a_n2354_n1288# 0.089328f
C68 plus.t22 a_n2354_n1288# 0.089328f
C69 plus.n3 a_n2354_n1288# 0.062388f
C70 plus.n4 a_n2354_n1288# 0.050595f
C71 plus.t14 a_n2354_n1288# 0.089328f
C72 plus.t8 a_n2354_n1288# 0.089328f
C73 plus.n5 a_n2354_n1288# 0.062388f
C74 plus.n6 a_n2354_n1288# 0.050595f
C75 plus.t23 a_n2354_n1288# 0.089328f
C76 plus.t17 a_n2354_n1288# 0.089328f
C77 plus.n7 a_n2354_n1288# 0.019436f
C78 plus.t4 a_n2354_n1288# 0.095986f
C79 plus.t9 a_n2354_n1288# 0.089328f
C80 plus.n8 a_n2354_n1288# 0.062388f
C81 plus.n9 a_n2354_n1288# 0.077106f
C82 plus.n10 a_n2354_n1288# 0.108297f
C83 plus.n11 a_n2354_n1288# 0.050595f
C84 plus.n12 a_n2354_n1288# 0.018188f
C85 plus.n13 a_n2354_n1288# 0.062388f
C86 plus.n14 a_n2354_n1288# 0.020839f
C87 plus.n15 a_n2354_n1288# 0.062388f
C88 plus.n16 a_n2354_n1288# 0.020839f
C89 plus.n17 a_n2354_n1288# 0.050595f
C90 plus.n18 a_n2354_n1288# 0.050595f
C91 plus.n19 a_n2354_n1288# 0.020839f
C92 plus.n20 a_n2354_n1288# 0.062388f
C93 plus.n21 a_n2354_n1288# 0.018812f
C94 plus.n22 a_n2354_n1288# 0.018812f
C95 plus.n23 a_n2354_n1288# 0.050595f
C96 plus.n24 a_n2354_n1288# 0.050595f
C97 plus.n25 a_n2354_n1288# 0.020839f
C98 plus.n26 a_n2354_n1288# 0.062388f
C99 plus.n27 a_n2354_n1288# 0.020839f
C100 plus.n28 a_n2354_n1288# 0.062388f
C101 plus.n29 a_n2354_n1288# 0.020839f
C102 plus.n30 a_n2354_n1288# 0.050595f
C103 plus.n31 a_n2354_n1288# 0.050595f
C104 plus.n32 a_n2354_n1288# 0.018188f
C105 plus.n33 a_n2354_n1288# 0.019436f
C106 plus.n34 a_n2354_n1288# 0.062388f
C107 plus.t5 a_n2354_n1288# 0.095986f
C108 plus.n35 a_n2354_n1288# 0.077038f
C109 plus.n36 a_n2354_n1288# 0.357952f
C110 plus.n37 a_n2354_n1288# 0.050595f
C111 plus.t11 a_n2354_n1288# 0.095986f
C112 plus.t21 a_n2354_n1288# 0.089328f
C113 plus.t6 a_n2354_n1288# 0.089328f
C114 plus.n38 a_n2354_n1288# 0.062388f
C115 plus.n39 a_n2354_n1288# 0.050595f
C116 plus.t16 a_n2354_n1288# 0.089328f
C117 plus.t18 a_n2354_n1288# 0.089328f
C118 plus.t3 a_n2354_n1288# 0.089328f
C119 plus.n40 a_n2354_n1288# 0.062388f
C120 plus.n41 a_n2354_n1288# 0.050595f
C121 plus.t12 a_n2354_n1288# 0.089328f
C122 plus.t15 a_n2354_n1288# 0.089328f
C123 plus.n42 a_n2354_n1288# 0.062388f
C124 plus.n43 a_n2354_n1288# 0.050595f
C125 plus.t1 a_n2354_n1288# 0.089328f
C126 plus.t7 a_n2354_n1288# 0.089328f
C127 plus.n44 a_n2354_n1288# 0.019436f
C128 plus.t10 a_n2354_n1288# 0.089328f
C129 plus.n45 a_n2354_n1288# 0.062388f
C130 plus.t20 a_n2354_n1288# 0.095986f
C131 plus.n46 a_n2354_n1288# 0.077106f
C132 plus.n47 a_n2354_n1288# 0.108297f
C133 plus.n48 a_n2354_n1288# 0.050595f
C134 plus.n49 a_n2354_n1288# 0.018188f
C135 plus.n50 a_n2354_n1288# 0.062388f
C136 plus.n51 a_n2354_n1288# 0.020839f
C137 plus.n52 a_n2354_n1288# 0.062388f
C138 plus.n53 a_n2354_n1288# 0.020839f
C139 plus.n54 a_n2354_n1288# 0.050595f
C140 plus.n55 a_n2354_n1288# 0.050595f
C141 plus.n56 a_n2354_n1288# 0.020839f
C142 plus.n57 a_n2354_n1288# 0.062388f
C143 plus.n58 a_n2354_n1288# 0.018812f
C144 plus.n59 a_n2354_n1288# 0.018812f
C145 plus.n60 a_n2354_n1288# 0.050595f
C146 plus.n61 a_n2354_n1288# 0.050595f
C147 plus.n62 a_n2354_n1288# 0.020839f
C148 plus.n63 a_n2354_n1288# 0.062388f
C149 plus.n64 a_n2354_n1288# 0.020839f
C150 plus.n65 a_n2354_n1288# 0.062388f
C151 plus.n66 a_n2354_n1288# 0.020839f
C152 plus.n67 a_n2354_n1288# 0.050595f
C153 plus.n68 a_n2354_n1288# 0.050595f
C154 plus.n69 a_n2354_n1288# 0.018188f
C155 plus.n70 a_n2354_n1288# 0.019436f
C156 plus.n71 a_n2354_n1288# 0.062388f
C157 plus.n72 a_n2354_n1288# 0.077038f
C158 plus.n73 a_n2354_n1288# 1.28201f
C159 drain_right.t22 a_n2354_n1288# 0.043003f
C160 drain_right.t5 a_n2354_n1288# 0.043003f
C161 drain_right.n0 a_n2354_n1288# 0.271843f
C162 drain_right.t10 a_n2354_n1288# 0.043003f
C163 drain_right.t17 a_n2354_n1288# 0.043003f
C164 drain_right.n1 a_n2354_n1288# 0.270158f
C165 drain_right.n2 a_n2354_n1288# 0.616251f
C166 drain_right.t4 a_n2354_n1288# 0.043003f
C167 drain_right.t6 a_n2354_n1288# 0.043003f
C168 drain_right.n3 a_n2354_n1288# 0.270158f
C169 drain_right.n4 a_n2354_n1288# 0.277746f
C170 drain_right.t12 a_n2354_n1288# 0.043003f
C171 drain_right.t23 a_n2354_n1288# 0.043003f
C172 drain_right.n5 a_n2354_n1288# 0.271843f
C173 drain_right.t8 a_n2354_n1288# 0.043003f
C174 drain_right.t11 a_n2354_n1288# 0.043003f
C175 drain_right.n6 a_n2354_n1288# 0.270158f
C176 drain_right.n7 a_n2354_n1288# 0.616251f
C177 drain_right.t15 a_n2354_n1288# 0.043003f
C178 drain_right.t16 a_n2354_n1288# 0.043003f
C179 drain_right.n8 a_n2354_n1288# 0.270158f
C180 drain_right.n9 a_n2354_n1288# 0.277746f
C181 drain_right.n10 a_n2354_n1288# 0.859694f
C182 drain_right.t1 a_n2354_n1288# 0.043003f
C183 drain_right.t7 a_n2354_n1288# 0.043003f
C184 drain_right.n11 a_n2354_n1288# 0.271844f
C185 drain_right.t9 a_n2354_n1288# 0.043003f
C186 drain_right.t20 a_n2354_n1288# 0.043003f
C187 drain_right.n12 a_n2354_n1288# 0.270159f
C188 drain_right.n13 a_n2354_n1288# 0.616249f
C189 drain_right.t21 a_n2354_n1288# 0.043003f
C190 drain_right.t3 a_n2354_n1288# 0.043003f
C191 drain_right.n14 a_n2354_n1288# 0.270159f
C192 drain_right.n15 a_n2354_n1288# 0.303487f
C193 drain_right.t0 a_n2354_n1288# 0.043003f
C194 drain_right.t14 a_n2354_n1288# 0.043003f
C195 drain_right.n16 a_n2354_n1288# 0.270159f
C196 drain_right.n17 a_n2354_n1288# 0.303487f
C197 drain_right.t13 a_n2354_n1288# 0.043003f
C198 drain_right.t19 a_n2354_n1288# 0.043003f
C199 drain_right.n18 a_n2354_n1288# 0.270159f
C200 drain_right.n19 a_n2354_n1288# 0.303487f
C201 drain_right.t18 a_n2354_n1288# 0.043003f
C202 drain_right.t2 a_n2354_n1288# 0.043003f
C203 drain_right.n20 a_n2354_n1288# 0.270159f
C204 drain_right.n21 a_n2354_n1288# 0.529966f
C205 source.n0 a_n2354_n1288# 0.051457f
C206 source.n1 a_n2354_n1288# 0.113855f
C207 source.t23 a_n2354_n1288# 0.085443f
C208 source.n2 a_n2354_n1288# 0.089108f
C209 source.n3 a_n2354_n1288# 0.028725f
C210 source.n4 a_n2354_n1288# 0.018945f
C211 source.n5 a_n2354_n1288# 0.250965f
C212 source.n6 a_n2354_n1288# 0.056409f
C213 source.n7 a_n2354_n1288# 0.532297f
C214 source.t17 a_n2354_n1288# 0.055719f
C215 source.t12 a_n2354_n1288# 0.055719f
C216 source.n8 a_n2354_n1288# 0.297875f
C217 source.n9 a_n2354_n1288# 0.397487f
C218 source.t14 a_n2354_n1288# 0.055719f
C219 source.t8 a_n2354_n1288# 0.055719f
C220 source.n10 a_n2354_n1288# 0.297875f
C221 source.n11 a_n2354_n1288# 0.397487f
C222 source.t10 a_n2354_n1288# 0.055719f
C223 source.t7 a_n2354_n1288# 0.055719f
C224 source.n12 a_n2354_n1288# 0.297875f
C225 source.n13 a_n2354_n1288# 0.397487f
C226 source.t2 a_n2354_n1288# 0.055719f
C227 source.t4 a_n2354_n1288# 0.055719f
C228 source.n14 a_n2354_n1288# 0.297875f
C229 source.n15 a_n2354_n1288# 0.397487f
C230 source.t9 a_n2354_n1288# 0.055719f
C231 source.t11 a_n2354_n1288# 0.055719f
C232 source.n16 a_n2354_n1288# 0.297875f
C233 source.n17 a_n2354_n1288# 0.397487f
C234 source.n18 a_n2354_n1288# 0.051457f
C235 source.n19 a_n2354_n1288# 0.113855f
C236 source.t19 a_n2354_n1288# 0.085443f
C237 source.n20 a_n2354_n1288# 0.089108f
C238 source.n21 a_n2354_n1288# 0.028725f
C239 source.n22 a_n2354_n1288# 0.018945f
C240 source.n23 a_n2354_n1288# 0.250965f
C241 source.n24 a_n2354_n1288# 0.056409f
C242 source.n25 a_n2354_n1288# 0.144093f
C243 source.n26 a_n2354_n1288# 0.051457f
C244 source.n27 a_n2354_n1288# 0.113855f
C245 source.t42 a_n2354_n1288# 0.085443f
C246 source.n28 a_n2354_n1288# 0.089108f
C247 source.n29 a_n2354_n1288# 0.028725f
C248 source.n30 a_n2354_n1288# 0.018945f
C249 source.n31 a_n2354_n1288# 0.250965f
C250 source.n32 a_n2354_n1288# 0.056409f
C251 source.n33 a_n2354_n1288# 0.144093f
C252 source.t44 a_n2354_n1288# 0.055719f
C253 source.t36 a_n2354_n1288# 0.055719f
C254 source.n34 a_n2354_n1288# 0.297875f
C255 source.n35 a_n2354_n1288# 0.397487f
C256 source.t29 a_n2354_n1288# 0.055719f
C257 source.t30 a_n2354_n1288# 0.055719f
C258 source.n36 a_n2354_n1288# 0.297875f
C259 source.n37 a_n2354_n1288# 0.397487f
C260 source.t43 a_n2354_n1288# 0.055719f
C261 source.t38 a_n2354_n1288# 0.055719f
C262 source.n38 a_n2354_n1288# 0.297875f
C263 source.n39 a_n2354_n1288# 0.397487f
C264 source.t45 a_n2354_n1288# 0.055719f
C265 source.t24 a_n2354_n1288# 0.055719f
C266 source.n40 a_n2354_n1288# 0.297875f
C267 source.n41 a_n2354_n1288# 0.397487f
C268 source.t32 a_n2354_n1288# 0.055719f
C269 source.t25 a_n2354_n1288# 0.055719f
C270 source.n42 a_n2354_n1288# 0.297875f
C271 source.n43 a_n2354_n1288# 0.397487f
C272 source.n44 a_n2354_n1288# 0.051457f
C273 source.n45 a_n2354_n1288# 0.113855f
C274 source.t46 a_n2354_n1288# 0.085443f
C275 source.n46 a_n2354_n1288# 0.089108f
C276 source.n47 a_n2354_n1288# 0.028725f
C277 source.n48 a_n2354_n1288# 0.018945f
C278 source.n49 a_n2354_n1288# 0.250965f
C279 source.n50 a_n2354_n1288# 0.056409f
C280 source.n51 a_n2354_n1288# 0.860983f
C281 source.n52 a_n2354_n1288# 0.051457f
C282 source.n53 a_n2354_n1288# 0.113855f
C283 source.t21 a_n2354_n1288# 0.085443f
C284 source.n54 a_n2354_n1288# 0.089108f
C285 source.n55 a_n2354_n1288# 0.028725f
C286 source.n56 a_n2354_n1288# 0.018945f
C287 source.n57 a_n2354_n1288# 0.250965f
C288 source.n58 a_n2354_n1288# 0.056409f
C289 source.n59 a_n2354_n1288# 0.860983f
C290 source.t3 a_n2354_n1288# 0.055719f
C291 source.t13 a_n2354_n1288# 0.055719f
C292 source.n60 a_n2354_n1288# 0.297873f
C293 source.n61 a_n2354_n1288# 0.397489f
C294 source.t20 a_n2354_n1288# 0.055719f
C295 source.t18 a_n2354_n1288# 0.055719f
C296 source.n62 a_n2354_n1288# 0.297873f
C297 source.n63 a_n2354_n1288# 0.397489f
C298 source.t6 a_n2354_n1288# 0.055719f
C299 source.t1 a_n2354_n1288# 0.055719f
C300 source.n64 a_n2354_n1288# 0.297873f
C301 source.n65 a_n2354_n1288# 0.397489f
C302 source.t15 a_n2354_n1288# 0.055719f
C303 source.t5 a_n2354_n1288# 0.055719f
C304 source.n66 a_n2354_n1288# 0.297873f
C305 source.n67 a_n2354_n1288# 0.397489f
C306 source.t0 a_n2354_n1288# 0.055719f
C307 source.t16 a_n2354_n1288# 0.055719f
C308 source.n68 a_n2354_n1288# 0.297873f
C309 source.n69 a_n2354_n1288# 0.397489f
C310 source.n70 a_n2354_n1288# 0.051457f
C311 source.n71 a_n2354_n1288# 0.113855f
C312 source.t22 a_n2354_n1288# 0.085443f
C313 source.n72 a_n2354_n1288# 0.089108f
C314 source.n73 a_n2354_n1288# 0.028725f
C315 source.n74 a_n2354_n1288# 0.018945f
C316 source.n75 a_n2354_n1288# 0.250965f
C317 source.n76 a_n2354_n1288# 0.056409f
C318 source.n77 a_n2354_n1288# 0.144093f
C319 source.n78 a_n2354_n1288# 0.051457f
C320 source.n79 a_n2354_n1288# 0.113855f
C321 source.t40 a_n2354_n1288# 0.085443f
C322 source.n80 a_n2354_n1288# 0.089108f
C323 source.n81 a_n2354_n1288# 0.028725f
C324 source.n82 a_n2354_n1288# 0.018945f
C325 source.n83 a_n2354_n1288# 0.250965f
C326 source.n84 a_n2354_n1288# 0.056409f
C327 source.n85 a_n2354_n1288# 0.144093f
C328 source.t33 a_n2354_n1288# 0.055719f
C329 source.t39 a_n2354_n1288# 0.055719f
C330 source.n86 a_n2354_n1288# 0.297873f
C331 source.n87 a_n2354_n1288# 0.397489f
C332 source.t37 a_n2354_n1288# 0.055719f
C333 source.t34 a_n2354_n1288# 0.055719f
C334 source.n88 a_n2354_n1288# 0.297873f
C335 source.n89 a_n2354_n1288# 0.397489f
C336 source.t28 a_n2354_n1288# 0.055719f
C337 source.t35 a_n2354_n1288# 0.055719f
C338 source.n90 a_n2354_n1288# 0.297873f
C339 source.n91 a_n2354_n1288# 0.397489f
C340 source.t47 a_n2354_n1288# 0.055719f
C341 source.t41 a_n2354_n1288# 0.055719f
C342 source.n92 a_n2354_n1288# 0.297873f
C343 source.n93 a_n2354_n1288# 0.397489f
C344 source.t26 a_n2354_n1288# 0.055719f
C345 source.t31 a_n2354_n1288# 0.055719f
C346 source.n94 a_n2354_n1288# 0.297873f
C347 source.n95 a_n2354_n1288# 0.397489f
C348 source.n96 a_n2354_n1288# 0.051457f
C349 source.n97 a_n2354_n1288# 0.113855f
C350 source.t27 a_n2354_n1288# 0.085443f
C351 source.n98 a_n2354_n1288# 0.089108f
C352 source.n99 a_n2354_n1288# 0.028725f
C353 source.n100 a_n2354_n1288# 0.018945f
C354 source.n101 a_n2354_n1288# 0.250965f
C355 source.n102 a_n2354_n1288# 0.056409f
C356 source.n103 a_n2354_n1288# 0.343108f
C357 source.n104 a_n2354_n1288# 0.871637f
C358 minus.n0 a_n2354_n1288# 0.03751f
C359 minus.t5 a_n2354_n1288# 0.071162f
C360 minus.t21 a_n2354_n1288# 0.066226f
C361 minus.t10 a_n2354_n1288# 0.066226f
C362 minus.n1 a_n2354_n1288# 0.046253f
C363 minus.n2 a_n2354_n1288# 0.03751f
C364 minus.t4 a_n2354_n1288# 0.066226f
C365 minus.t23 a_n2354_n1288# 0.066226f
C366 minus.t9 a_n2354_n1288# 0.066226f
C367 minus.n3 a_n2354_n1288# 0.046253f
C368 minus.n4 a_n2354_n1288# 0.03751f
C369 minus.t2 a_n2354_n1288# 0.066226f
C370 minus.t20 a_n2354_n1288# 0.066226f
C371 minus.n5 a_n2354_n1288# 0.046253f
C372 minus.n6 a_n2354_n1288# 0.03751f
C373 minus.t14 a_n2354_n1288# 0.066226f
C374 minus.t3 a_n2354_n1288# 0.066226f
C375 minus.n7 a_n2354_n1288# 0.014409f
C376 minus.t22 a_n2354_n1288# 0.066226f
C377 minus.n8 a_n2354_n1288# 0.046253f
C378 minus.t16 a_n2354_n1288# 0.071162f
C379 minus.n9 a_n2354_n1288# 0.057165f
C380 minus.n10 a_n2354_n1288# 0.080289f
C381 minus.n11 a_n2354_n1288# 0.03751f
C382 minus.n12 a_n2354_n1288# 0.013484f
C383 minus.n13 a_n2354_n1288# 0.046253f
C384 minus.n14 a_n2354_n1288# 0.01545f
C385 minus.n15 a_n2354_n1288# 0.046253f
C386 minus.n16 a_n2354_n1288# 0.01545f
C387 minus.n17 a_n2354_n1288# 0.03751f
C388 minus.n18 a_n2354_n1288# 0.03751f
C389 minus.n19 a_n2354_n1288# 0.01545f
C390 minus.n20 a_n2354_n1288# 0.046253f
C391 minus.n21 a_n2354_n1288# 0.013947f
C392 minus.n22 a_n2354_n1288# 0.013947f
C393 minus.n23 a_n2354_n1288# 0.03751f
C394 minus.n24 a_n2354_n1288# 0.03751f
C395 minus.n25 a_n2354_n1288# 0.01545f
C396 minus.n26 a_n2354_n1288# 0.046253f
C397 minus.n27 a_n2354_n1288# 0.01545f
C398 minus.n28 a_n2354_n1288# 0.046253f
C399 minus.n29 a_n2354_n1288# 0.01545f
C400 minus.n30 a_n2354_n1288# 0.03751f
C401 minus.n31 a_n2354_n1288# 0.03751f
C402 minus.n32 a_n2354_n1288# 0.013484f
C403 minus.n33 a_n2354_n1288# 0.014409f
C404 minus.n34 a_n2354_n1288# 0.046253f
C405 minus.n35 a_n2354_n1288# 0.057115f
C406 minus.n36 a_n2354_n1288# 0.998819f
C407 minus.n37 a_n2354_n1288# 0.03751f
C408 minus.t11 a_n2354_n1288# 0.066226f
C409 minus.t12 a_n2354_n1288# 0.066226f
C410 minus.n38 a_n2354_n1288# 0.046253f
C411 minus.n39 a_n2354_n1288# 0.03751f
C412 minus.t15 a_n2354_n1288# 0.066226f
C413 minus.t7 a_n2354_n1288# 0.066226f
C414 minus.t8 a_n2354_n1288# 0.066226f
C415 minus.n40 a_n2354_n1288# 0.046253f
C416 minus.n41 a_n2354_n1288# 0.03751f
C417 minus.t17 a_n2354_n1288# 0.066226f
C418 minus.t19 a_n2354_n1288# 0.066226f
C419 minus.n42 a_n2354_n1288# 0.046253f
C420 minus.n43 a_n2354_n1288# 0.03751f
C421 minus.t6 a_n2354_n1288# 0.066226f
C422 minus.t13 a_n2354_n1288# 0.066226f
C423 minus.n44 a_n2354_n1288# 0.014409f
C424 minus.t1 a_n2354_n1288# 0.071162f
C425 minus.t18 a_n2354_n1288# 0.066226f
C426 minus.n45 a_n2354_n1288# 0.046253f
C427 minus.n46 a_n2354_n1288# 0.057165f
C428 minus.n47 a_n2354_n1288# 0.080289f
C429 minus.n48 a_n2354_n1288# 0.03751f
C430 minus.n49 a_n2354_n1288# 0.013484f
C431 minus.n50 a_n2354_n1288# 0.046253f
C432 minus.n51 a_n2354_n1288# 0.01545f
C433 minus.n52 a_n2354_n1288# 0.046253f
C434 minus.n53 a_n2354_n1288# 0.01545f
C435 minus.n54 a_n2354_n1288# 0.03751f
C436 minus.n55 a_n2354_n1288# 0.03751f
C437 minus.n56 a_n2354_n1288# 0.01545f
C438 minus.n57 a_n2354_n1288# 0.046253f
C439 minus.n58 a_n2354_n1288# 0.013947f
C440 minus.n59 a_n2354_n1288# 0.013947f
C441 minus.n60 a_n2354_n1288# 0.03751f
C442 minus.n61 a_n2354_n1288# 0.03751f
C443 minus.n62 a_n2354_n1288# 0.01545f
C444 minus.n63 a_n2354_n1288# 0.046253f
C445 minus.n64 a_n2354_n1288# 0.01545f
C446 minus.n65 a_n2354_n1288# 0.046253f
C447 minus.n66 a_n2354_n1288# 0.01545f
C448 minus.n67 a_n2354_n1288# 0.03751f
C449 minus.n68 a_n2354_n1288# 0.03751f
C450 minus.n69 a_n2354_n1288# 0.013484f
C451 minus.n70 a_n2354_n1288# 0.014409f
C452 minus.n71 a_n2354_n1288# 0.046253f
C453 minus.t0 a_n2354_n1288# 0.071162f
C454 minus.n72 a_n2354_n1288# 0.057115f
C455 minus.n73 a_n2354_n1288# 0.242595f
C456 minus.n74 a_n2354_n1288# 1.23259f
.ends

