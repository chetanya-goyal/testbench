* NGSPICE file created from diffpair241.ext - technology: sky130A

.subckt diffpair241 minus drain_right drain_left source plus
X0 drain_right minus source a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X1 source plus drain_left a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X2 source minus drain_right a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X3 a_n1106_n2092# a_n1106_n2092# a_n1106_n2092# a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=22.8 ps=103.6 w=6 l=0.15
X4 drain_left plus source a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X5 drain_left plus source a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X6 drain_right minus source a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X7 a_n1106_n2092# a_n1106_n2092# a_n1106_n2092# a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X8 source plus drain_left a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X9 a_n1106_n2092# a_n1106_n2092# a_n1106_n2092# a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X10 a_n1106_n2092# a_n1106_n2092# a_n1106_n2092# a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X11 source minus drain_right a_n1106_n2092# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
.ends

