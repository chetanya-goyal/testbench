* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right.t19 minus.t0 source.t23 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X1 drain_right.t18 minus.t1 source.t22 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X2 drain_right.t17 minus.t2 source.t24 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X3 source.t30 minus.t3 drain_right.t16 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X4 source.t13 plus.t0 drain_left.t19 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X5 source.t9 plus.t1 drain_left.t18 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X6 source.t26 minus.t4 drain_right.t15 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X7 source.t10 plus.t2 drain_left.t17 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X8 source.t12 plus.t3 drain_left.t16 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X9 source.t35 minus.t5 drain_right.t14 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X10 source.t8 plus.t4 drain_left.t15 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X11 source.t21 minus.t6 drain_right.t13 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X12 drain_left.t14 plus.t5 source.t17 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X13 drain_right.t12 minus.t7 source.t33 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X14 drain_right.t11 minus.t8 source.t28 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X15 source.t31 minus.t9 drain_right.t10 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X16 drain_left.t13 plus.t6 source.t3 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X17 a_n2542_n1288# a_n2542_n1288# a_n2542_n1288# a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.5
X18 drain_left.t12 plus.t7 source.t1 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X19 drain_left.t11 plus.t8 source.t2 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X20 source.t5 plus.t9 drain_left.t10 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X21 source.t29 minus.t10 drain_right.t9 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X22 a_n2542_n1288# a_n2542_n1288# a_n2542_n1288# a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X23 source.t39 minus.t11 drain_right.t8 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X24 drain_right.t7 minus.t12 source.t34 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X25 source.t11 plus.t10 drain_left.t9 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X26 drain_left.t8 plus.t11 source.t14 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X27 drain_right.t6 minus.t13 source.t38 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X28 drain_right.t5 minus.t14 source.t32 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X29 source.t0 plus.t12 drain_left.t7 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X30 drain_left.t6 plus.t13 source.t15 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X31 drain_right.t4 minus.t15 source.t20 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X32 source.t27 minus.t16 drain_right.t3 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X33 a_n2542_n1288# a_n2542_n1288# a_n2542_n1288# a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X34 source.t25 minus.t17 drain_right.t2 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X35 drain_left.t5 plus.t14 source.t7 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X36 source.t36 minus.t18 drain_right.t1 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X37 source.t16 plus.t15 drain_left.t4 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X38 drain_right.t0 minus.t19 source.t37 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X39 drain_left.t3 plus.t16 source.t19 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X40 source.t4 plus.t17 drain_left.t2 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X41 a_n2542_n1288# a_n2542_n1288# a_n2542_n1288# a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X42 drain_left.t1 plus.t18 source.t18 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X43 drain_left.t0 plus.t19 source.t6 a_n2542_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
R0 minus.n6 minus.t13 195.948
R1 minus.n34 minus.t18 195.948
R2 minus.n7 minus.t4 174.966
R3 minus.n5 minus.t8 174.966
R4 minus.n13 minus.t17 174.966
R5 minus.n14 minus.t7 174.966
R6 minus.n18 minus.t10 174.966
R7 minus.n19 minus.t1 174.966
R8 minus.n1 minus.t11 174.966
R9 minus.n25 minus.t15 174.966
R10 minus.n26 minus.t5 174.966
R11 minus.n35 minus.t0 174.966
R12 minus.n33 minus.t16 174.966
R13 minus.n41 minus.t19 174.966
R14 minus.n42 minus.t9 174.966
R15 minus.n46 minus.t2 174.966
R16 minus.n47 minus.t6 174.966
R17 minus.n29 minus.t14 174.966
R18 minus.n53 minus.t3 174.966
R19 minus.n54 minus.t12 174.966
R20 minus.n27 minus.n26 161.3
R21 minus.n25 minus.n0 161.3
R22 minus.n24 minus.n23 161.3
R23 minus.n22 minus.n1 161.3
R24 minus.n21 minus.n20 161.3
R25 minus.n19 minus.n2 161.3
R26 minus.n18 minus.n17 161.3
R27 minus.n16 minus.n3 161.3
R28 minus.n15 minus.n14 161.3
R29 minus.n13 minus.n4 161.3
R30 minus.n12 minus.n11 161.3
R31 minus.n10 minus.n5 161.3
R32 minus.n9 minus.n8 161.3
R33 minus.n55 minus.n54 161.3
R34 minus.n53 minus.n28 161.3
R35 minus.n52 minus.n51 161.3
R36 minus.n50 minus.n29 161.3
R37 minus.n49 minus.n48 161.3
R38 minus.n47 minus.n30 161.3
R39 minus.n46 minus.n45 161.3
R40 minus.n44 minus.n31 161.3
R41 minus.n43 minus.n42 161.3
R42 minus.n41 minus.n32 161.3
R43 minus.n40 minus.n39 161.3
R44 minus.n38 minus.n33 161.3
R45 minus.n37 minus.n36 161.3
R46 minus.n9 minus.n6 70.4033
R47 minus.n37 minus.n34 70.4033
R48 minus.n14 minus.n13 48.2005
R49 minus.n19 minus.n18 48.2005
R50 minus.n26 minus.n25 48.2005
R51 minus.n42 minus.n41 48.2005
R52 minus.n47 minus.n46 48.2005
R53 minus.n54 minus.n53 48.2005
R54 minus.n12 minus.n5 47.4702
R55 minus.n20 minus.n1 47.4702
R56 minus.n40 minus.n33 47.4702
R57 minus.n48 minus.n29 47.4702
R58 minus.n56 minus.n27 31.2657
R59 minus.n8 minus.n5 25.5611
R60 minus.n24 minus.n1 25.5611
R61 minus.n36 minus.n33 25.5611
R62 minus.n52 minus.n29 25.5611
R63 minus.n18 minus.n3 24.1005
R64 minus.n14 minus.n3 24.1005
R65 minus.n42 minus.n31 24.1005
R66 minus.n46 minus.n31 24.1005
R67 minus.n8 minus.n7 22.6399
R68 minus.n25 minus.n24 22.6399
R69 minus.n36 minus.n35 22.6399
R70 minus.n53 minus.n52 22.6399
R71 minus.n7 minus.n6 20.9576
R72 minus.n35 minus.n34 20.9576
R73 minus.n56 minus.n55 6.59141
R74 minus.n13 minus.n12 0.730803
R75 minus.n20 minus.n19 0.730803
R76 minus.n41 minus.n40 0.730803
R77 minus.n48 minus.n47 0.730803
R78 minus.n27 minus.n0 0.189894
R79 minus.n23 minus.n0 0.189894
R80 minus.n23 minus.n22 0.189894
R81 minus.n22 minus.n21 0.189894
R82 minus.n21 minus.n2 0.189894
R83 minus.n17 minus.n2 0.189894
R84 minus.n17 minus.n16 0.189894
R85 minus.n16 minus.n15 0.189894
R86 minus.n15 minus.n4 0.189894
R87 minus.n11 minus.n4 0.189894
R88 minus.n11 minus.n10 0.189894
R89 minus.n10 minus.n9 0.189894
R90 minus.n38 minus.n37 0.189894
R91 minus.n39 minus.n38 0.189894
R92 minus.n39 minus.n32 0.189894
R93 minus.n43 minus.n32 0.189894
R94 minus.n44 minus.n43 0.189894
R95 minus.n45 minus.n44 0.189894
R96 minus.n45 minus.n30 0.189894
R97 minus.n49 minus.n30 0.189894
R98 minus.n50 minus.n49 0.189894
R99 minus.n51 minus.n50 0.189894
R100 minus.n51 minus.n28 0.189894
R101 minus.n55 minus.n28 0.189894
R102 minus minus.n56 0.188
R103 source.n90 source.n88 289.615
R104 source.n74 source.n72 289.615
R105 source.n66 source.n64 289.615
R106 source.n50 source.n48 289.615
R107 source.n2 source.n0 289.615
R108 source.n18 source.n16 289.615
R109 source.n26 source.n24 289.615
R110 source.n42 source.n40 289.615
R111 source.n91 source.n90 185
R112 source.n75 source.n74 185
R113 source.n67 source.n66 185
R114 source.n51 source.n50 185
R115 source.n3 source.n2 185
R116 source.n19 source.n18 185
R117 source.n27 source.n26 185
R118 source.n43 source.n42 185
R119 source.t34 source.n89 167.117
R120 source.t36 source.n73 167.117
R121 source.t18 source.n65 167.117
R122 source.t11 source.n49 167.117
R123 source.t14 source.n1 167.117
R124 source.t12 source.n17 167.117
R125 source.t38 source.n25 167.117
R126 source.t35 source.n41 167.117
R127 source.n9 source.n8 84.1169
R128 source.n11 source.n10 84.1169
R129 source.n13 source.n12 84.1169
R130 source.n15 source.n14 84.1169
R131 source.n33 source.n32 84.1169
R132 source.n35 source.n34 84.1169
R133 source.n37 source.n36 84.1169
R134 source.n39 source.n38 84.1169
R135 source.n87 source.n86 84.1168
R136 source.n85 source.n84 84.1168
R137 source.n83 source.n82 84.1168
R138 source.n81 source.n80 84.1168
R139 source.n63 source.n62 84.1168
R140 source.n61 source.n60 84.1168
R141 source.n59 source.n58 84.1168
R142 source.n57 source.n56 84.1168
R143 source.n90 source.t34 52.3082
R144 source.n74 source.t36 52.3082
R145 source.n66 source.t18 52.3082
R146 source.n50 source.t11 52.3082
R147 source.n2 source.t14 52.3082
R148 source.n18 source.t12 52.3082
R149 source.n26 source.t38 52.3082
R150 source.n42 source.t35 52.3082
R151 source.n95 source.n94 31.4096
R152 source.n79 source.n78 31.4096
R153 source.n71 source.n70 31.4096
R154 source.n55 source.n54 31.4096
R155 source.n7 source.n6 31.4096
R156 source.n23 source.n22 31.4096
R157 source.n31 source.n30 31.4096
R158 source.n47 source.n46 31.4096
R159 source.n55 source.n47 14.4275
R160 source.n86 source.t32 9.9005
R161 source.n86 source.t30 9.9005
R162 source.n84 source.t24 9.9005
R163 source.n84 source.t21 9.9005
R164 source.n82 source.t37 9.9005
R165 source.n82 source.t31 9.9005
R166 source.n80 source.t23 9.9005
R167 source.n80 source.t27 9.9005
R168 source.n62 source.t7 9.9005
R169 source.n62 source.t9 9.9005
R170 source.n60 source.t2 9.9005
R171 source.n60 source.t8 9.9005
R172 source.n58 source.t17 9.9005
R173 source.n58 source.t13 9.9005
R174 source.n56 source.t3 9.9005
R175 source.n56 source.t0 9.9005
R176 source.n8 source.t19 9.9005
R177 source.n8 source.t10 9.9005
R178 source.n10 source.t6 9.9005
R179 source.n10 source.t5 9.9005
R180 source.n12 source.t1 9.9005
R181 source.n12 source.t16 9.9005
R182 source.n14 source.t15 9.9005
R183 source.n14 source.t4 9.9005
R184 source.n32 source.t28 9.9005
R185 source.n32 source.t26 9.9005
R186 source.n34 source.t33 9.9005
R187 source.n34 source.t25 9.9005
R188 source.n36 source.t22 9.9005
R189 source.n36 source.t29 9.9005
R190 source.n38 source.t20 9.9005
R191 source.n38 source.t39 9.9005
R192 source.n91 source.n89 9.71174
R193 source.n75 source.n73 9.71174
R194 source.n67 source.n65 9.71174
R195 source.n51 source.n49 9.71174
R196 source.n3 source.n1 9.71174
R197 source.n19 source.n17 9.71174
R198 source.n27 source.n25 9.71174
R199 source.n43 source.n41 9.71174
R200 source.n94 source.n93 9.45567
R201 source.n78 source.n77 9.45567
R202 source.n70 source.n69 9.45567
R203 source.n54 source.n53 9.45567
R204 source.n6 source.n5 9.45567
R205 source.n22 source.n21 9.45567
R206 source.n30 source.n29 9.45567
R207 source.n46 source.n45 9.45567
R208 source.n93 source.n92 9.3005
R209 source.n77 source.n76 9.3005
R210 source.n69 source.n68 9.3005
R211 source.n53 source.n52 9.3005
R212 source.n5 source.n4 9.3005
R213 source.n21 source.n20 9.3005
R214 source.n29 source.n28 9.3005
R215 source.n45 source.n44 9.3005
R216 source.n96 source.n7 8.8068
R217 source.n94 source.n88 8.14595
R218 source.n78 source.n72 8.14595
R219 source.n70 source.n64 8.14595
R220 source.n54 source.n48 8.14595
R221 source.n6 source.n0 8.14595
R222 source.n22 source.n16 8.14595
R223 source.n30 source.n24 8.14595
R224 source.n46 source.n40 8.14595
R225 source.n92 source.n91 7.3702
R226 source.n76 source.n75 7.3702
R227 source.n68 source.n67 7.3702
R228 source.n52 source.n51 7.3702
R229 source.n4 source.n3 7.3702
R230 source.n20 source.n19 7.3702
R231 source.n28 source.n27 7.3702
R232 source.n44 source.n43 7.3702
R233 source.n92 source.n88 5.81868
R234 source.n76 source.n72 5.81868
R235 source.n68 source.n64 5.81868
R236 source.n52 source.n48 5.81868
R237 source.n4 source.n0 5.81868
R238 source.n20 source.n16 5.81868
R239 source.n28 source.n24 5.81868
R240 source.n44 source.n40 5.81868
R241 source.n96 source.n95 5.62119
R242 source.n93 source.n89 3.44771
R243 source.n77 source.n73 3.44771
R244 source.n69 source.n65 3.44771
R245 source.n53 source.n49 3.44771
R246 source.n5 source.n1 3.44771
R247 source.n21 source.n17 3.44771
R248 source.n29 source.n25 3.44771
R249 source.n45 source.n41 3.44771
R250 source.n47 source.n39 0.716017
R251 source.n39 source.n37 0.716017
R252 source.n37 source.n35 0.716017
R253 source.n35 source.n33 0.716017
R254 source.n33 source.n31 0.716017
R255 source.n23 source.n15 0.716017
R256 source.n15 source.n13 0.716017
R257 source.n13 source.n11 0.716017
R258 source.n11 source.n9 0.716017
R259 source.n9 source.n7 0.716017
R260 source.n57 source.n55 0.716017
R261 source.n59 source.n57 0.716017
R262 source.n61 source.n59 0.716017
R263 source.n63 source.n61 0.716017
R264 source.n71 source.n63 0.716017
R265 source.n81 source.n79 0.716017
R266 source.n83 source.n81 0.716017
R267 source.n85 source.n83 0.716017
R268 source.n87 source.n85 0.716017
R269 source.n95 source.n87 0.716017
R270 source.n31 source.n23 0.470328
R271 source.n79 source.n71 0.470328
R272 source source.n96 0.188
R273 drain_right.n10 drain_right.n8 101.511
R274 drain_right.n6 drain_right.n4 101.511
R275 drain_right.n2 drain_right.n0 101.511
R276 drain_right.n10 drain_right.n9 100.796
R277 drain_right.n12 drain_right.n11 100.796
R278 drain_right.n14 drain_right.n13 100.796
R279 drain_right.n16 drain_right.n15 100.796
R280 drain_right.n7 drain_right.n3 100.796
R281 drain_right.n6 drain_right.n5 100.796
R282 drain_right.n2 drain_right.n1 100.796
R283 drain_right drain_right.n7 24.9622
R284 drain_right.n3 drain_right.t10 9.9005
R285 drain_right.n3 drain_right.t17 9.9005
R286 drain_right.n4 drain_right.t16 9.9005
R287 drain_right.n4 drain_right.t7 9.9005
R288 drain_right.n5 drain_right.t13 9.9005
R289 drain_right.n5 drain_right.t5 9.9005
R290 drain_right.n1 drain_right.t3 9.9005
R291 drain_right.n1 drain_right.t0 9.9005
R292 drain_right.n0 drain_right.t1 9.9005
R293 drain_right.n0 drain_right.t19 9.9005
R294 drain_right.n8 drain_right.t15 9.9005
R295 drain_right.n8 drain_right.t6 9.9005
R296 drain_right.n9 drain_right.t2 9.9005
R297 drain_right.n9 drain_right.t11 9.9005
R298 drain_right.n11 drain_right.t9 9.9005
R299 drain_right.n11 drain_right.t12 9.9005
R300 drain_right.n13 drain_right.t8 9.9005
R301 drain_right.n13 drain_right.t18 9.9005
R302 drain_right.n15 drain_right.t14 9.9005
R303 drain_right.n15 drain_right.t4 9.9005
R304 drain_right drain_right.n16 6.36873
R305 drain_right.n16 drain_right.n14 0.716017
R306 drain_right.n14 drain_right.n12 0.716017
R307 drain_right.n12 drain_right.n10 0.716017
R308 drain_right.n7 drain_right.n6 0.660671
R309 drain_right.n7 drain_right.n2 0.660671
R310 plus.n8 plus.t3 195.948
R311 plus.n36 plus.t18 195.948
R312 plus.n26 plus.t11 174.966
R313 plus.n25 plus.t2 174.966
R314 plus.n1 plus.t16 174.966
R315 plus.n19 plus.t9 174.966
R316 plus.n18 plus.t19 174.966
R317 plus.n4 plus.t15 174.966
R318 plus.n13 plus.t7 174.966
R319 plus.n11 plus.t17 174.966
R320 plus.n7 plus.t13 174.966
R321 plus.n54 plus.t10 174.966
R322 plus.n53 plus.t6 174.966
R323 plus.n29 plus.t12 174.966
R324 plus.n47 plus.t5 174.966
R325 plus.n46 plus.t0 174.966
R326 plus.n32 plus.t8 174.966
R327 plus.n41 plus.t4 174.966
R328 plus.n39 plus.t14 174.966
R329 plus.n35 plus.t1 174.966
R330 plus.n10 plus.n9 161.3
R331 plus.n11 plus.n6 161.3
R332 plus.n12 plus.n5 161.3
R333 plus.n14 plus.n13 161.3
R334 plus.n15 plus.n4 161.3
R335 plus.n17 plus.n16 161.3
R336 plus.n18 plus.n3 161.3
R337 plus.n19 plus.n2 161.3
R338 plus.n21 plus.n20 161.3
R339 plus.n22 plus.n1 161.3
R340 plus.n24 plus.n23 161.3
R341 plus.n25 plus.n0 161.3
R342 plus.n27 plus.n26 161.3
R343 plus.n38 plus.n37 161.3
R344 plus.n39 plus.n34 161.3
R345 plus.n40 plus.n33 161.3
R346 plus.n42 plus.n41 161.3
R347 plus.n43 plus.n32 161.3
R348 plus.n45 plus.n44 161.3
R349 plus.n46 plus.n31 161.3
R350 plus.n47 plus.n30 161.3
R351 plus.n49 plus.n48 161.3
R352 plus.n50 plus.n29 161.3
R353 plus.n52 plus.n51 161.3
R354 plus.n53 plus.n28 161.3
R355 plus.n55 plus.n54 161.3
R356 plus.n9 plus.n8 70.4033
R357 plus.n37 plus.n36 70.4033
R358 plus.n26 plus.n25 48.2005
R359 plus.n19 plus.n18 48.2005
R360 plus.n13 plus.n4 48.2005
R361 plus.n54 plus.n53 48.2005
R362 plus.n47 plus.n46 48.2005
R363 plus.n41 plus.n32 48.2005
R364 plus.n20 plus.n1 47.4702
R365 plus.n12 plus.n11 47.4702
R366 plus.n48 plus.n29 47.4702
R367 plus.n40 plus.n39 47.4702
R368 plus plus.n55 28.9346
R369 plus.n24 plus.n1 25.5611
R370 plus.n11 plus.n10 25.5611
R371 plus.n52 plus.n29 25.5611
R372 plus.n39 plus.n38 25.5611
R373 plus.n17 plus.n4 24.1005
R374 plus.n18 plus.n17 24.1005
R375 plus.n46 plus.n45 24.1005
R376 plus.n45 plus.n32 24.1005
R377 plus.n25 plus.n24 22.6399
R378 plus.n10 plus.n7 22.6399
R379 plus.n53 plus.n52 22.6399
R380 plus.n38 plus.n35 22.6399
R381 plus.n8 plus.n7 20.9576
R382 plus.n36 plus.n35 20.9576
R383 plus plus.n27 8.44747
R384 plus.n20 plus.n19 0.730803
R385 plus.n13 plus.n12 0.730803
R386 plus.n48 plus.n47 0.730803
R387 plus.n41 plus.n40 0.730803
R388 plus.n9 plus.n6 0.189894
R389 plus.n6 plus.n5 0.189894
R390 plus.n14 plus.n5 0.189894
R391 plus.n15 plus.n14 0.189894
R392 plus.n16 plus.n15 0.189894
R393 plus.n16 plus.n3 0.189894
R394 plus.n3 plus.n2 0.189894
R395 plus.n21 plus.n2 0.189894
R396 plus.n22 plus.n21 0.189894
R397 plus.n23 plus.n22 0.189894
R398 plus.n23 plus.n0 0.189894
R399 plus.n27 plus.n0 0.189894
R400 plus.n55 plus.n28 0.189894
R401 plus.n51 plus.n28 0.189894
R402 plus.n51 plus.n50 0.189894
R403 plus.n50 plus.n49 0.189894
R404 plus.n49 plus.n30 0.189894
R405 plus.n31 plus.n30 0.189894
R406 plus.n44 plus.n31 0.189894
R407 plus.n44 plus.n43 0.189894
R408 plus.n43 plus.n42 0.189894
R409 plus.n42 plus.n33 0.189894
R410 plus.n34 plus.n33 0.189894
R411 plus.n37 plus.n34 0.189894
R412 drain_left.n10 drain_left.n8 101.511
R413 drain_left.n6 drain_left.n4 101.511
R414 drain_left.n2 drain_left.n0 101.511
R415 drain_left.n16 drain_left.n15 100.796
R416 drain_left.n14 drain_left.n13 100.796
R417 drain_left.n12 drain_left.n11 100.796
R418 drain_left.n10 drain_left.n9 100.796
R419 drain_left.n7 drain_left.n3 100.796
R420 drain_left.n6 drain_left.n5 100.796
R421 drain_left.n2 drain_left.n1 100.796
R422 drain_left drain_left.n7 25.5155
R423 drain_left.n3 drain_left.t19 9.9005
R424 drain_left.n3 drain_left.t11 9.9005
R425 drain_left.n4 drain_left.t18 9.9005
R426 drain_left.n4 drain_left.t1 9.9005
R427 drain_left.n5 drain_left.t15 9.9005
R428 drain_left.n5 drain_left.t5 9.9005
R429 drain_left.n1 drain_left.t7 9.9005
R430 drain_left.n1 drain_left.t14 9.9005
R431 drain_left.n0 drain_left.t9 9.9005
R432 drain_left.n0 drain_left.t13 9.9005
R433 drain_left.n15 drain_left.t17 9.9005
R434 drain_left.n15 drain_left.t8 9.9005
R435 drain_left.n13 drain_left.t10 9.9005
R436 drain_left.n13 drain_left.t3 9.9005
R437 drain_left.n11 drain_left.t4 9.9005
R438 drain_left.n11 drain_left.t0 9.9005
R439 drain_left.n9 drain_left.t2 9.9005
R440 drain_left.n9 drain_left.t12 9.9005
R441 drain_left.n8 drain_left.t16 9.9005
R442 drain_left.n8 drain_left.t6 9.9005
R443 drain_left drain_left.n16 6.36873
R444 drain_left.n12 drain_left.n10 0.716017
R445 drain_left.n14 drain_left.n12 0.716017
R446 drain_left.n16 drain_left.n14 0.716017
R447 drain_left.n7 drain_left.n6 0.660671
R448 drain_left.n7 drain_left.n2 0.660671
C0 minus drain_left 0.179153f
C1 source minus 2.76186f
C2 minus drain_right 2.24303f
C3 minus plus 4.47617f
C4 source drain_left 7.85654f
C5 drain_right drain_left 1.3588f
C6 drain_left plus 2.49468f
C7 source drain_right 7.857871f
C8 source plus 2.77583f
C9 drain_right plus 0.415087f
C10 drain_right a_n2542_n1288# 4.95758f
C11 drain_left a_n2542_n1288# 5.34866f
C12 source a_n2542_n1288# 3.378014f
C13 minus a_n2542_n1288# 9.301064f
C14 plus a_n2542_n1288# 10.67516f
C15 drain_left.t9 a_n2542_n1288# 0.045619f
C16 drain_left.t13 a_n2542_n1288# 0.045619f
C17 drain_left.n0 a_n2542_n1288# 0.289171f
C18 drain_left.t7 a_n2542_n1288# 0.045619f
C19 drain_left.t14 a_n2542_n1288# 0.045619f
C20 drain_left.n1 a_n2542_n1288# 0.286594f
C21 drain_left.n2 a_n2542_n1288# 0.712962f
C22 drain_left.t19 a_n2542_n1288# 0.045619f
C23 drain_left.t11 a_n2542_n1288# 0.045619f
C24 drain_left.n3 a_n2542_n1288# 0.286594f
C25 drain_left.t18 a_n2542_n1288# 0.045619f
C26 drain_left.t1 a_n2542_n1288# 0.045619f
C27 drain_left.n4 a_n2542_n1288# 0.289171f
C28 drain_left.t15 a_n2542_n1288# 0.045619f
C29 drain_left.t5 a_n2542_n1288# 0.045619f
C30 drain_left.n5 a_n2542_n1288# 0.286594f
C31 drain_left.n6 a_n2542_n1288# 0.712962f
C32 drain_left.n7 a_n2542_n1288# 1.32592f
C33 drain_left.t16 a_n2542_n1288# 0.045619f
C34 drain_left.t6 a_n2542_n1288# 0.045619f
C35 drain_left.n8 a_n2542_n1288# 0.289172f
C36 drain_left.t2 a_n2542_n1288# 0.045619f
C37 drain_left.t12 a_n2542_n1288# 0.045619f
C38 drain_left.n9 a_n2542_n1288# 0.286595f
C39 drain_left.n10 a_n2542_n1288# 0.717093f
C40 drain_left.t4 a_n2542_n1288# 0.045619f
C41 drain_left.t0 a_n2542_n1288# 0.045619f
C42 drain_left.n11 a_n2542_n1288# 0.286595f
C43 drain_left.n12 a_n2542_n1288# 0.354022f
C44 drain_left.t10 a_n2542_n1288# 0.045619f
C45 drain_left.t3 a_n2542_n1288# 0.045619f
C46 drain_left.n13 a_n2542_n1288# 0.286595f
C47 drain_left.n14 a_n2542_n1288# 0.354022f
C48 drain_left.t17 a_n2542_n1288# 0.045619f
C49 drain_left.t8 a_n2542_n1288# 0.045619f
C50 drain_left.n15 a_n2542_n1288# 0.286595f
C51 drain_left.n16 a_n2542_n1288# 0.602008f
C52 plus.n0 a_n2542_n1288# 0.0475f
C53 plus.t11 a_n2542_n1288# 0.147095f
C54 plus.t2 a_n2542_n1288# 0.147095f
C55 plus.t16 a_n2542_n1288# 0.147095f
C56 plus.n1 a_n2542_n1288# 0.110937f
C57 plus.n2 a_n2542_n1288# 0.0475f
C58 plus.t9 a_n2542_n1288# 0.147095f
C59 plus.t19 a_n2542_n1288# 0.147095f
C60 plus.n3 a_n2542_n1288# 0.0475f
C61 plus.t15 a_n2542_n1288# 0.147095f
C62 plus.n4 a_n2542_n1288# 0.11079f
C63 plus.n5 a_n2542_n1288# 0.0475f
C64 plus.t7 a_n2542_n1288# 0.147095f
C65 plus.t17 a_n2542_n1288# 0.147095f
C66 plus.n6 a_n2542_n1288# 0.0475f
C67 plus.t13 a_n2542_n1288# 0.147095f
C68 plus.n7 a_n2542_n1288# 0.110497f
C69 plus.t3 a_n2542_n1288# 0.158448f
C70 plus.n8 a_n2542_n1288# 0.094969f
C71 plus.n9 a_n2542_n1288# 0.155901f
C72 plus.n10 a_n2542_n1288# 0.010779f
C73 plus.n11 a_n2542_n1288# 0.110937f
C74 plus.n12 a_n2542_n1288# 0.010779f
C75 plus.n13 a_n2542_n1288# 0.106104f
C76 plus.n14 a_n2542_n1288# 0.0475f
C77 plus.n15 a_n2542_n1288# 0.0475f
C78 plus.n16 a_n2542_n1288# 0.0475f
C79 plus.n17 a_n2542_n1288# 0.010779f
C80 plus.n18 a_n2542_n1288# 0.11079f
C81 plus.n19 a_n2542_n1288# 0.106104f
C82 plus.n20 a_n2542_n1288# 0.010779f
C83 plus.n21 a_n2542_n1288# 0.0475f
C84 plus.n22 a_n2542_n1288# 0.0475f
C85 plus.n23 a_n2542_n1288# 0.0475f
C86 plus.n24 a_n2542_n1288# 0.010779f
C87 plus.n25 a_n2542_n1288# 0.110497f
C88 plus.n26 a_n2542_n1288# 0.105958f
C89 plus.n27 a_n2542_n1288# 0.350313f
C90 plus.n28 a_n2542_n1288# 0.0475f
C91 plus.t10 a_n2542_n1288# 0.147095f
C92 plus.t6 a_n2542_n1288# 0.147095f
C93 plus.t12 a_n2542_n1288# 0.147095f
C94 plus.n29 a_n2542_n1288# 0.110937f
C95 plus.n30 a_n2542_n1288# 0.0475f
C96 plus.t5 a_n2542_n1288# 0.147095f
C97 plus.n31 a_n2542_n1288# 0.0475f
C98 plus.t0 a_n2542_n1288# 0.147095f
C99 plus.t8 a_n2542_n1288# 0.147095f
C100 plus.n32 a_n2542_n1288# 0.11079f
C101 plus.n33 a_n2542_n1288# 0.0475f
C102 plus.t4 a_n2542_n1288# 0.147095f
C103 plus.n34 a_n2542_n1288# 0.0475f
C104 plus.t14 a_n2542_n1288# 0.147095f
C105 plus.t1 a_n2542_n1288# 0.147095f
C106 plus.n35 a_n2542_n1288# 0.110497f
C107 plus.t18 a_n2542_n1288# 0.158448f
C108 plus.n36 a_n2542_n1288# 0.094969f
C109 plus.n37 a_n2542_n1288# 0.155901f
C110 plus.n38 a_n2542_n1288# 0.010779f
C111 plus.n39 a_n2542_n1288# 0.110937f
C112 plus.n40 a_n2542_n1288# 0.010779f
C113 plus.n41 a_n2542_n1288# 0.106104f
C114 plus.n42 a_n2542_n1288# 0.0475f
C115 plus.n43 a_n2542_n1288# 0.0475f
C116 plus.n44 a_n2542_n1288# 0.0475f
C117 plus.n45 a_n2542_n1288# 0.010779f
C118 plus.n46 a_n2542_n1288# 0.11079f
C119 plus.n47 a_n2542_n1288# 0.106104f
C120 plus.n48 a_n2542_n1288# 0.010779f
C121 plus.n49 a_n2542_n1288# 0.0475f
C122 plus.n50 a_n2542_n1288# 0.0475f
C123 plus.n51 a_n2542_n1288# 0.0475f
C124 plus.n52 a_n2542_n1288# 0.010779f
C125 plus.n53 a_n2542_n1288# 0.110497f
C126 plus.n54 a_n2542_n1288# 0.105958f
C127 plus.n55 a_n2542_n1288# 1.26423f
C128 drain_right.t1 a_n2542_n1288# 0.04479f
C129 drain_right.t19 a_n2542_n1288# 0.04479f
C130 drain_right.n0 a_n2542_n1288# 0.283912f
C131 drain_right.t3 a_n2542_n1288# 0.04479f
C132 drain_right.t0 a_n2542_n1288# 0.04479f
C133 drain_right.n1 a_n2542_n1288# 0.281381f
C134 drain_right.n2 a_n2542_n1288# 0.699995f
C135 drain_right.t10 a_n2542_n1288# 0.04479f
C136 drain_right.t17 a_n2542_n1288# 0.04479f
C137 drain_right.n3 a_n2542_n1288# 0.281381f
C138 drain_right.t16 a_n2542_n1288# 0.04479f
C139 drain_right.t7 a_n2542_n1288# 0.04479f
C140 drain_right.n4 a_n2542_n1288# 0.283912f
C141 drain_right.t13 a_n2542_n1288# 0.04479f
C142 drain_right.t5 a_n2542_n1288# 0.04479f
C143 drain_right.n5 a_n2542_n1288# 0.281381f
C144 drain_right.n6 a_n2542_n1288# 0.699995f
C145 drain_right.n7 a_n2542_n1288# 1.24666f
C146 drain_right.t15 a_n2542_n1288# 0.04479f
C147 drain_right.t6 a_n2542_n1288# 0.04479f
C148 drain_right.n8 a_n2542_n1288# 0.283913f
C149 drain_right.t2 a_n2542_n1288# 0.04479f
C150 drain_right.t11 a_n2542_n1288# 0.04479f
C151 drain_right.n9 a_n2542_n1288# 0.281383f
C152 drain_right.n10 a_n2542_n1288# 0.704052f
C153 drain_right.t9 a_n2542_n1288# 0.04479f
C154 drain_right.t12 a_n2542_n1288# 0.04479f
C155 drain_right.n11 a_n2542_n1288# 0.281383f
C156 drain_right.n12 a_n2542_n1288# 0.347584f
C157 drain_right.t8 a_n2542_n1288# 0.04479f
C158 drain_right.t18 a_n2542_n1288# 0.04479f
C159 drain_right.n13 a_n2542_n1288# 0.281383f
C160 drain_right.n14 a_n2542_n1288# 0.347584f
C161 drain_right.t14 a_n2542_n1288# 0.04479f
C162 drain_right.t4 a_n2542_n1288# 0.04479f
C163 drain_right.n15 a_n2542_n1288# 0.281383f
C164 drain_right.n16 a_n2542_n1288# 0.59106f
C165 source.n0 a_n2542_n1288# 0.04699f
C166 source.n1 a_n2542_n1288# 0.10397f
C167 source.t14 a_n2542_n1288# 0.078025f
C168 source.n2 a_n2542_n1288# 0.081371f
C169 source.n3 a_n2542_n1288# 0.026231f
C170 source.n4 a_n2542_n1288# 0.0173f
C171 source.n5 a_n2542_n1288# 0.229176f
C172 source.n6 a_n2542_n1288# 0.051512f
C173 source.n7 a_n2542_n1288# 0.51782f
C174 source.t19 a_n2542_n1288# 0.050882f
C175 source.t10 a_n2542_n1288# 0.050882f
C176 source.n8 a_n2542_n1288# 0.272014f
C177 source.n9 a_n2542_n1288# 0.398748f
C178 source.t6 a_n2542_n1288# 0.050882f
C179 source.t5 a_n2542_n1288# 0.050882f
C180 source.n10 a_n2542_n1288# 0.272014f
C181 source.n11 a_n2542_n1288# 0.398748f
C182 source.t1 a_n2542_n1288# 0.050882f
C183 source.t16 a_n2542_n1288# 0.050882f
C184 source.n12 a_n2542_n1288# 0.272014f
C185 source.n13 a_n2542_n1288# 0.398748f
C186 source.t15 a_n2542_n1288# 0.050882f
C187 source.t4 a_n2542_n1288# 0.050882f
C188 source.n14 a_n2542_n1288# 0.272014f
C189 source.n15 a_n2542_n1288# 0.398748f
C190 source.n16 a_n2542_n1288# 0.04699f
C191 source.n17 a_n2542_n1288# 0.10397f
C192 source.t12 a_n2542_n1288# 0.078025f
C193 source.n18 a_n2542_n1288# 0.081371f
C194 source.n19 a_n2542_n1288# 0.026231f
C195 source.n20 a_n2542_n1288# 0.0173f
C196 source.n21 a_n2542_n1288# 0.229176f
C197 source.n22 a_n2542_n1288# 0.051512f
C198 source.n23 a_n2542_n1288# 0.149469f
C199 source.n24 a_n2542_n1288# 0.04699f
C200 source.n25 a_n2542_n1288# 0.10397f
C201 source.t38 a_n2542_n1288# 0.078025f
C202 source.n26 a_n2542_n1288# 0.081371f
C203 source.n27 a_n2542_n1288# 0.026231f
C204 source.n28 a_n2542_n1288# 0.0173f
C205 source.n29 a_n2542_n1288# 0.229176f
C206 source.n30 a_n2542_n1288# 0.051512f
C207 source.n31 a_n2542_n1288# 0.149469f
C208 source.t28 a_n2542_n1288# 0.050882f
C209 source.t26 a_n2542_n1288# 0.050882f
C210 source.n32 a_n2542_n1288# 0.272014f
C211 source.n33 a_n2542_n1288# 0.398748f
C212 source.t33 a_n2542_n1288# 0.050882f
C213 source.t25 a_n2542_n1288# 0.050882f
C214 source.n34 a_n2542_n1288# 0.272014f
C215 source.n35 a_n2542_n1288# 0.398748f
C216 source.t22 a_n2542_n1288# 0.050882f
C217 source.t29 a_n2542_n1288# 0.050882f
C218 source.n36 a_n2542_n1288# 0.272014f
C219 source.n37 a_n2542_n1288# 0.398748f
C220 source.t20 a_n2542_n1288# 0.050882f
C221 source.t39 a_n2542_n1288# 0.050882f
C222 source.n38 a_n2542_n1288# 0.272014f
C223 source.n39 a_n2542_n1288# 0.398748f
C224 source.n40 a_n2542_n1288# 0.04699f
C225 source.n41 a_n2542_n1288# 0.10397f
C226 source.t35 a_n2542_n1288# 0.078025f
C227 source.n42 a_n2542_n1288# 0.081371f
C228 source.n43 a_n2542_n1288# 0.026231f
C229 source.n44 a_n2542_n1288# 0.0173f
C230 source.n45 a_n2542_n1288# 0.229176f
C231 source.n46 a_n2542_n1288# 0.051512f
C232 source.n47 a_n2542_n1288# 0.822004f
C233 source.n48 a_n2542_n1288# 0.04699f
C234 source.n49 a_n2542_n1288# 0.10397f
C235 source.t11 a_n2542_n1288# 0.078025f
C236 source.n50 a_n2542_n1288# 0.081371f
C237 source.n51 a_n2542_n1288# 0.026231f
C238 source.n52 a_n2542_n1288# 0.0173f
C239 source.n53 a_n2542_n1288# 0.229176f
C240 source.n54 a_n2542_n1288# 0.051512f
C241 source.n55 a_n2542_n1288# 0.822004f
C242 source.t3 a_n2542_n1288# 0.050882f
C243 source.t0 a_n2542_n1288# 0.050882f
C244 source.n56 a_n2542_n1288# 0.272012f
C245 source.n57 a_n2542_n1288# 0.39875f
C246 source.t17 a_n2542_n1288# 0.050882f
C247 source.t13 a_n2542_n1288# 0.050882f
C248 source.n58 a_n2542_n1288# 0.272012f
C249 source.n59 a_n2542_n1288# 0.39875f
C250 source.t2 a_n2542_n1288# 0.050882f
C251 source.t8 a_n2542_n1288# 0.050882f
C252 source.n60 a_n2542_n1288# 0.272012f
C253 source.n61 a_n2542_n1288# 0.39875f
C254 source.t7 a_n2542_n1288# 0.050882f
C255 source.t9 a_n2542_n1288# 0.050882f
C256 source.n62 a_n2542_n1288# 0.272012f
C257 source.n63 a_n2542_n1288# 0.39875f
C258 source.n64 a_n2542_n1288# 0.04699f
C259 source.n65 a_n2542_n1288# 0.10397f
C260 source.t18 a_n2542_n1288# 0.078025f
C261 source.n66 a_n2542_n1288# 0.081371f
C262 source.n67 a_n2542_n1288# 0.026231f
C263 source.n68 a_n2542_n1288# 0.0173f
C264 source.n69 a_n2542_n1288# 0.229176f
C265 source.n70 a_n2542_n1288# 0.051512f
C266 source.n71 a_n2542_n1288# 0.149469f
C267 source.n72 a_n2542_n1288# 0.04699f
C268 source.n73 a_n2542_n1288# 0.10397f
C269 source.t36 a_n2542_n1288# 0.078025f
C270 source.n74 a_n2542_n1288# 0.081371f
C271 source.n75 a_n2542_n1288# 0.026231f
C272 source.n76 a_n2542_n1288# 0.0173f
C273 source.n77 a_n2542_n1288# 0.229176f
C274 source.n78 a_n2542_n1288# 0.051512f
C275 source.n79 a_n2542_n1288# 0.149469f
C276 source.t23 a_n2542_n1288# 0.050882f
C277 source.t27 a_n2542_n1288# 0.050882f
C278 source.n80 a_n2542_n1288# 0.272012f
C279 source.n81 a_n2542_n1288# 0.39875f
C280 source.t37 a_n2542_n1288# 0.050882f
C281 source.t31 a_n2542_n1288# 0.050882f
C282 source.n82 a_n2542_n1288# 0.272012f
C283 source.n83 a_n2542_n1288# 0.39875f
C284 source.t24 a_n2542_n1288# 0.050882f
C285 source.t21 a_n2542_n1288# 0.050882f
C286 source.n84 a_n2542_n1288# 0.272012f
C287 source.n85 a_n2542_n1288# 0.39875f
C288 source.t32 a_n2542_n1288# 0.050882f
C289 source.t30 a_n2542_n1288# 0.050882f
C290 source.n86 a_n2542_n1288# 0.272012f
C291 source.n87 a_n2542_n1288# 0.39875f
C292 source.n88 a_n2542_n1288# 0.04699f
C293 source.n89 a_n2542_n1288# 0.10397f
C294 source.t34 a_n2542_n1288# 0.078025f
C295 source.n90 a_n2542_n1288# 0.081371f
C296 source.n91 a_n2542_n1288# 0.026231f
C297 source.n92 a_n2542_n1288# 0.0173f
C298 source.n93 a_n2542_n1288# 0.229176f
C299 source.n94 a_n2542_n1288# 0.051512f
C300 source.n95 a_n2542_n1288# 0.345419f
C301 source.n96 a_n2542_n1288# 0.803668f
C302 minus.n0 a_n2542_n1288# 0.045599f
C303 minus.t11 a_n2542_n1288# 0.141208f
C304 minus.n1 a_n2542_n1288# 0.106497f
C305 minus.n2 a_n2542_n1288# 0.045599f
C306 minus.n3 a_n2542_n1288# 0.010347f
C307 minus.t10 a_n2542_n1288# 0.141208f
C308 minus.n4 a_n2542_n1288# 0.045599f
C309 minus.t8 a_n2542_n1288# 0.141208f
C310 minus.n5 a_n2542_n1288# 0.106497f
C311 minus.t13 a_n2542_n1288# 0.152107f
C312 minus.n6 a_n2542_n1288# 0.091168f
C313 minus.t4 a_n2542_n1288# 0.141208f
C314 minus.n7 a_n2542_n1288# 0.106075f
C315 minus.n8 a_n2542_n1288# 0.010347f
C316 minus.n9 a_n2542_n1288# 0.149661f
C317 minus.n10 a_n2542_n1288# 0.045599f
C318 minus.n11 a_n2542_n1288# 0.045599f
C319 minus.n12 a_n2542_n1288# 0.010347f
C320 minus.t17 a_n2542_n1288# 0.141208f
C321 minus.n13 a_n2542_n1288# 0.101858f
C322 minus.t7 a_n2542_n1288# 0.141208f
C323 minus.n14 a_n2542_n1288# 0.106356f
C324 minus.n15 a_n2542_n1288# 0.045599f
C325 minus.n16 a_n2542_n1288# 0.045599f
C326 minus.n17 a_n2542_n1288# 0.045599f
C327 minus.n18 a_n2542_n1288# 0.106356f
C328 minus.t1 a_n2542_n1288# 0.141208f
C329 minus.n19 a_n2542_n1288# 0.101858f
C330 minus.n20 a_n2542_n1288# 0.010347f
C331 minus.n21 a_n2542_n1288# 0.045599f
C332 minus.n22 a_n2542_n1288# 0.045599f
C333 minus.n23 a_n2542_n1288# 0.045599f
C334 minus.n24 a_n2542_n1288# 0.010347f
C335 minus.t15 a_n2542_n1288# 0.141208f
C336 minus.n25 a_n2542_n1288# 0.106075f
C337 minus.t5 a_n2542_n1288# 0.141208f
C338 minus.n26 a_n2542_n1288# 0.101717f
C339 minus.n27 a_n2542_n1288# 1.27574f
C340 minus.n28 a_n2542_n1288# 0.045599f
C341 minus.t14 a_n2542_n1288# 0.141208f
C342 minus.n29 a_n2542_n1288# 0.106497f
C343 minus.n30 a_n2542_n1288# 0.045599f
C344 minus.n31 a_n2542_n1288# 0.010347f
C345 minus.n32 a_n2542_n1288# 0.045599f
C346 minus.t16 a_n2542_n1288# 0.141208f
C347 minus.n33 a_n2542_n1288# 0.106497f
C348 minus.t18 a_n2542_n1288# 0.152107f
C349 minus.n34 a_n2542_n1288# 0.091168f
C350 minus.t0 a_n2542_n1288# 0.141208f
C351 minus.n35 a_n2542_n1288# 0.106075f
C352 minus.n36 a_n2542_n1288# 0.010347f
C353 minus.n37 a_n2542_n1288# 0.149661f
C354 minus.n38 a_n2542_n1288# 0.045599f
C355 minus.n39 a_n2542_n1288# 0.045599f
C356 minus.n40 a_n2542_n1288# 0.010347f
C357 minus.t19 a_n2542_n1288# 0.141208f
C358 minus.n41 a_n2542_n1288# 0.101858f
C359 minus.t9 a_n2542_n1288# 0.141208f
C360 minus.n42 a_n2542_n1288# 0.106356f
C361 minus.n43 a_n2542_n1288# 0.045599f
C362 minus.n44 a_n2542_n1288# 0.045599f
C363 minus.n45 a_n2542_n1288# 0.045599f
C364 minus.t2 a_n2542_n1288# 0.141208f
C365 minus.n46 a_n2542_n1288# 0.106356f
C366 minus.t6 a_n2542_n1288# 0.141208f
C367 minus.n47 a_n2542_n1288# 0.101858f
C368 minus.n48 a_n2542_n1288# 0.010347f
C369 minus.n49 a_n2542_n1288# 0.045599f
C370 minus.n50 a_n2542_n1288# 0.045599f
C371 minus.n51 a_n2542_n1288# 0.045599f
C372 minus.n52 a_n2542_n1288# 0.010347f
C373 minus.t3 a_n2542_n1288# 0.141208f
C374 minus.n53 a_n2542_n1288# 0.106075f
C375 minus.t12 a_n2542_n1288# 0.141208f
C376 minus.n54 a_n2542_n1288# 0.101717f
C377 minus.n55 a_n2542_n1288# 0.307893f
C378 minus.n56 a_n2542_n1288# 1.56557f
.ends

