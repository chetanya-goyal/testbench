* NGSPICE file created from diffpair475.ext - technology: sky130A

.subckt diffpair475 minus drain_right drain_left source plus
X0 drain_right.t11 minus.t0 source.t18 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X1 a_n2298_n3288# a_n2298_n3288# a_n2298_n3288# a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.8
X2 drain_right.t10 minus.t1 source.t10 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X3 source.t23 plus.t0 drain_left.t11 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X4 source.t8 plus.t1 drain_left.t10 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X5 a_n2298_n3288# a_n2298_n3288# a_n2298_n3288# a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.8
X6 drain_right.t9 minus.t2 source.t20 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X7 drain_right.t8 minus.t3 source.t12 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X8 source.t16 minus.t4 drain_right.t7 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X9 drain_right.t6 minus.t5 source.t17 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X10 source.t15 minus.t6 drain_right.t5 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
X11 a_n2298_n3288# a_n2298_n3288# a_n2298_n3288# a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.8
X12 drain_left.t9 plus.t2 source.t5 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X13 source.t14 minus.t7 drain_right.t4 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X14 drain_left.t8 plus.t3 source.t9 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X15 drain_right.t3 minus.t8 source.t13 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X16 source.t19 minus.t9 drain_right.t2 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X17 a_n2298_n3288# a_n2298_n3288# a_n2298_n3288# a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.8
X18 drain_left.t7 plus.t4 source.t4 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X19 drain_left.t6 plus.t5 source.t22 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X20 source.t6 plus.t6 drain_left.t5 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X21 drain_left.t4 plus.t7 source.t7 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X22 source.t0 plus.t8 drain_left.t3 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X23 drain_left.t2 plus.t9 source.t2 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X24 source.t11 minus.t10 drain_right.t1 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X25 source.t1 plus.t10 drain_left.t1 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
X26 source.t21 minus.t11 drain_right.t0 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
X27 source.t3 plus.t11 drain_left.t0 a_n2298_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
R0 minus.n4 minus.t5 432
R1 minus.n20 minus.t11 432
R2 minus.n3 minus.t4 410.604
R3 minus.n7 minus.t3 410.604
R4 minus.n8 minus.t7 410.604
R5 minus.n12 minus.t8 410.604
R6 minus.n14 minus.t6 410.604
R7 minus.n19 minus.t2 410.604
R8 minus.n23 minus.t9 410.604
R9 minus.n24 minus.t1 410.604
R10 minus.n28 minus.t10 410.604
R11 minus.n30 minus.t0 410.604
R12 minus.n15 minus.n14 161.3
R13 minus.n13 minus.n0 161.3
R14 minus.n12 minus.n11 161.3
R15 minus.n10 minus.n1 161.3
R16 minus.n6 minus.n5 161.3
R17 minus.n31 minus.n30 161.3
R18 minus.n29 minus.n16 161.3
R19 minus.n28 minus.n27 161.3
R20 minus.n26 minus.n17 161.3
R21 minus.n22 minus.n21 161.3
R22 minus.n9 minus.n8 80.6037
R23 minus.n7 minus.n2 80.6037
R24 minus.n25 minus.n24 80.6037
R25 minus.n23 minus.n18 80.6037
R26 minus.n8 minus.n7 48.2005
R27 minus.n24 minus.n23 48.2005
R28 minus.n5 minus.n4 44.853
R29 minus.n21 minus.n20 44.853
R30 minus.n7 minus.n6 41.6278
R31 minus.n8 minus.n1 41.6278
R32 minus.n23 minus.n22 41.6278
R33 minus.n24 minus.n17 41.6278
R34 minus.n32 minus.n15 38.027
R35 minus.n14 minus.n13 25.5611
R36 minus.n30 minus.n29 25.5611
R37 minus.n13 minus.n12 22.6399
R38 minus.n29 minus.n28 22.6399
R39 minus.n4 minus.n3 20.5405
R40 minus.n20 minus.n19 20.5405
R41 minus.n32 minus.n31 6.70126
R42 minus.n6 minus.n3 6.57323
R43 minus.n12 minus.n1 6.57323
R44 minus.n22 minus.n19 6.57323
R45 minus.n28 minus.n17 6.57323
R46 minus.n9 minus.n2 0.380177
R47 minus.n25 minus.n18 0.380177
R48 minus.n10 minus.n9 0.285035
R49 minus.n5 minus.n2 0.285035
R50 minus.n21 minus.n18 0.285035
R51 minus.n26 minus.n25 0.285035
R52 minus.n15 minus.n0 0.189894
R53 minus.n11 minus.n0 0.189894
R54 minus.n11 minus.n10 0.189894
R55 minus.n27 minus.n26 0.189894
R56 minus.n27 minus.n16 0.189894
R57 minus.n31 minus.n16 0.189894
R58 minus minus.n32 0.188
R59 source.n538 source.n478 289.615
R60 source.n468 source.n408 289.615
R61 source.n402 source.n342 289.615
R62 source.n332 source.n272 289.615
R63 source.n60 source.n0 289.615
R64 source.n130 source.n70 289.615
R65 source.n196 source.n136 289.615
R66 source.n266 source.n206 289.615
R67 source.n498 source.n497 185
R68 source.n503 source.n502 185
R69 source.n505 source.n504 185
R70 source.n494 source.n493 185
R71 source.n511 source.n510 185
R72 source.n513 source.n512 185
R73 source.n490 source.n489 185
R74 source.n520 source.n519 185
R75 source.n521 source.n488 185
R76 source.n523 source.n522 185
R77 source.n486 source.n485 185
R78 source.n529 source.n528 185
R79 source.n531 source.n530 185
R80 source.n482 source.n481 185
R81 source.n537 source.n536 185
R82 source.n539 source.n538 185
R83 source.n428 source.n427 185
R84 source.n433 source.n432 185
R85 source.n435 source.n434 185
R86 source.n424 source.n423 185
R87 source.n441 source.n440 185
R88 source.n443 source.n442 185
R89 source.n420 source.n419 185
R90 source.n450 source.n449 185
R91 source.n451 source.n418 185
R92 source.n453 source.n452 185
R93 source.n416 source.n415 185
R94 source.n459 source.n458 185
R95 source.n461 source.n460 185
R96 source.n412 source.n411 185
R97 source.n467 source.n466 185
R98 source.n469 source.n468 185
R99 source.n362 source.n361 185
R100 source.n367 source.n366 185
R101 source.n369 source.n368 185
R102 source.n358 source.n357 185
R103 source.n375 source.n374 185
R104 source.n377 source.n376 185
R105 source.n354 source.n353 185
R106 source.n384 source.n383 185
R107 source.n385 source.n352 185
R108 source.n387 source.n386 185
R109 source.n350 source.n349 185
R110 source.n393 source.n392 185
R111 source.n395 source.n394 185
R112 source.n346 source.n345 185
R113 source.n401 source.n400 185
R114 source.n403 source.n402 185
R115 source.n292 source.n291 185
R116 source.n297 source.n296 185
R117 source.n299 source.n298 185
R118 source.n288 source.n287 185
R119 source.n305 source.n304 185
R120 source.n307 source.n306 185
R121 source.n284 source.n283 185
R122 source.n314 source.n313 185
R123 source.n315 source.n282 185
R124 source.n317 source.n316 185
R125 source.n280 source.n279 185
R126 source.n323 source.n322 185
R127 source.n325 source.n324 185
R128 source.n276 source.n275 185
R129 source.n331 source.n330 185
R130 source.n333 source.n332 185
R131 source.n61 source.n60 185
R132 source.n59 source.n58 185
R133 source.n4 source.n3 185
R134 source.n53 source.n52 185
R135 source.n51 source.n50 185
R136 source.n8 source.n7 185
R137 source.n45 source.n44 185
R138 source.n43 source.n10 185
R139 source.n42 source.n41 185
R140 source.n13 source.n11 185
R141 source.n36 source.n35 185
R142 source.n34 source.n33 185
R143 source.n17 source.n16 185
R144 source.n28 source.n27 185
R145 source.n26 source.n25 185
R146 source.n21 source.n20 185
R147 source.n131 source.n130 185
R148 source.n129 source.n128 185
R149 source.n74 source.n73 185
R150 source.n123 source.n122 185
R151 source.n121 source.n120 185
R152 source.n78 source.n77 185
R153 source.n115 source.n114 185
R154 source.n113 source.n80 185
R155 source.n112 source.n111 185
R156 source.n83 source.n81 185
R157 source.n106 source.n105 185
R158 source.n104 source.n103 185
R159 source.n87 source.n86 185
R160 source.n98 source.n97 185
R161 source.n96 source.n95 185
R162 source.n91 source.n90 185
R163 source.n197 source.n196 185
R164 source.n195 source.n194 185
R165 source.n140 source.n139 185
R166 source.n189 source.n188 185
R167 source.n187 source.n186 185
R168 source.n144 source.n143 185
R169 source.n181 source.n180 185
R170 source.n179 source.n146 185
R171 source.n178 source.n177 185
R172 source.n149 source.n147 185
R173 source.n172 source.n171 185
R174 source.n170 source.n169 185
R175 source.n153 source.n152 185
R176 source.n164 source.n163 185
R177 source.n162 source.n161 185
R178 source.n157 source.n156 185
R179 source.n267 source.n266 185
R180 source.n265 source.n264 185
R181 source.n210 source.n209 185
R182 source.n259 source.n258 185
R183 source.n257 source.n256 185
R184 source.n214 source.n213 185
R185 source.n251 source.n250 185
R186 source.n249 source.n216 185
R187 source.n248 source.n247 185
R188 source.n219 source.n217 185
R189 source.n242 source.n241 185
R190 source.n240 source.n239 185
R191 source.n223 source.n222 185
R192 source.n234 source.n233 185
R193 source.n232 source.n231 185
R194 source.n227 source.n226 185
R195 source.n499 source.t18 149.524
R196 source.n429 source.t21 149.524
R197 source.n363 source.t7 149.524
R198 source.n293 source.t3 149.524
R199 source.n22 source.t4 149.524
R200 source.n92 source.t1 149.524
R201 source.n158 source.t17 149.524
R202 source.n228 source.t15 149.524
R203 source.n503 source.n497 104.615
R204 source.n504 source.n503 104.615
R205 source.n504 source.n493 104.615
R206 source.n511 source.n493 104.615
R207 source.n512 source.n511 104.615
R208 source.n512 source.n489 104.615
R209 source.n520 source.n489 104.615
R210 source.n521 source.n520 104.615
R211 source.n522 source.n521 104.615
R212 source.n522 source.n485 104.615
R213 source.n529 source.n485 104.615
R214 source.n530 source.n529 104.615
R215 source.n530 source.n481 104.615
R216 source.n537 source.n481 104.615
R217 source.n538 source.n537 104.615
R218 source.n433 source.n427 104.615
R219 source.n434 source.n433 104.615
R220 source.n434 source.n423 104.615
R221 source.n441 source.n423 104.615
R222 source.n442 source.n441 104.615
R223 source.n442 source.n419 104.615
R224 source.n450 source.n419 104.615
R225 source.n451 source.n450 104.615
R226 source.n452 source.n451 104.615
R227 source.n452 source.n415 104.615
R228 source.n459 source.n415 104.615
R229 source.n460 source.n459 104.615
R230 source.n460 source.n411 104.615
R231 source.n467 source.n411 104.615
R232 source.n468 source.n467 104.615
R233 source.n367 source.n361 104.615
R234 source.n368 source.n367 104.615
R235 source.n368 source.n357 104.615
R236 source.n375 source.n357 104.615
R237 source.n376 source.n375 104.615
R238 source.n376 source.n353 104.615
R239 source.n384 source.n353 104.615
R240 source.n385 source.n384 104.615
R241 source.n386 source.n385 104.615
R242 source.n386 source.n349 104.615
R243 source.n393 source.n349 104.615
R244 source.n394 source.n393 104.615
R245 source.n394 source.n345 104.615
R246 source.n401 source.n345 104.615
R247 source.n402 source.n401 104.615
R248 source.n297 source.n291 104.615
R249 source.n298 source.n297 104.615
R250 source.n298 source.n287 104.615
R251 source.n305 source.n287 104.615
R252 source.n306 source.n305 104.615
R253 source.n306 source.n283 104.615
R254 source.n314 source.n283 104.615
R255 source.n315 source.n314 104.615
R256 source.n316 source.n315 104.615
R257 source.n316 source.n279 104.615
R258 source.n323 source.n279 104.615
R259 source.n324 source.n323 104.615
R260 source.n324 source.n275 104.615
R261 source.n331 source.n275 104.615
R262 source.n332 source.n331 104.615
R263 source.n60 source.n59 104.615
R264 source.n59 source.n3 104.615
R265 source.n52 source.n3 104.615
R266 source.n52 source.n51 104.615
R267 source.n51 source.n7 104.615
R268 source.n44 source.n7 104.615
R269 source.n44 source.n43 104.615
R270 source.n43 source.n42 104.615
R271 source.n42 source.n11 104.615
R272 source.n35 source.n11 104.615
R273 source.n35 source.n34 104.615
R274 source.n34 source.n16 104.615
R275 source.n27 source.n16 104.615
R276 source.n27 source.n26 104.615
R277 source.n26 source.n20 104.615
R278 source.n130 source.n129 104.615
R279 source.n129 source.n73 104.615
R280 source.n122 source.n73 104.615
R281 source.n122 source.n121 104.615
R282 source.n121 source.n77 104.615
R283 source.n114 source.n77 104.615
R284 source.n114 source.n113 104.615
R285 source.n113 source.n112 104.615
R286 source.n112 source.n81 104.615
R287 source.n105 source.n81 104.615
R288 source.n105 source.n104 104.615
R289 source.n104 source.n86 104.615
R290 source.n97 source.n86 104.615
R291 source.n97 source.n96 104.615
R292 source.n96 source.n90 104.615
R293 source.n196 source.n195 104.615
R294 source.n195 source.n139 104.615
R295 source.n188 source.n139 104.615
R296 source.n188 source.n187 104.615
R297 source.n187 source.n143 104.615
R298 source.n180 source.n143 104.615
R299 source.n180 source.n179 104.615
R300 source.n179 source.n178 104.615
R301 source.n178 source.n147 104.615
R302 source.n171 source.n147 104.615
R303 source.n171 source.n170 104.615
R304 source.n170 source.n152 104.615
R305 source.n163 source.n152 104.615
R306 source.n163 source.n162 104.615
R307 source.n162 source.n156 104.615
R308 source.n266 source.n265 104.615
R309 source.n265 source.n209 104.615
R310 source.n258 source.n209 104.615
R311 source.n258 source.n257 104.615
R312 source.n257 source.n213 104.615
R313 source.n250 source.n213 104.615
R314 source.n250 source.n249 104.615
R315 source.n249 source.n248 104.615
R316 source.n248 source.n217 104.615
R317 source.n241 source.n217 104.615
R318 source.n241 source.n240 104.615
R319 source.n240 source.n222 104.615
R320 source.n233 source.n222 104.615
R321 source.n233 source.n232 104.615
R322 source.n232 source.n226 104.615
R323 source.t18 source.n497 52.3082
R324 source.t21 source.n427 52.3082
R325 source.t7 source.n361 52.3082
R326 source.t3 source.n291 52.3082
R327 source.t4 source.n20 52.3082
R328 source.t1 source.n90 52.3082
R329 source.t17 source.n156 52.3082
R330 source.t15 source.n226 52.3082
R331 source.n67 source.n66 42.8739
R332 source.n69 source.n68 42.8739
R333 source.n203 source.n202 42.8739
R334 source.n205 source.n204 42.8739
R335 source.n477 source.n476 42.8737
R336 source.n475 source.n474 42.8737
R337 source.n341 source.n340 42.8737
R338 source.n339 source.n338 42.8737
R339 source.n543 source.n542 29.8581
R340 source.n473 source.n472 29.8581
R341 source.n407 source.n406 29.8581
R342 source.n337 source.n336 29.8581
R343 source.n65 source.n64 29.8581
R344 source.n135 source.n134 29.8581
R345 source.n201 source.n200 29.8581
R346 source.n271 source.n270 29.8581
R347 source.n337 source.n271 22.2619
R348 source.n544 source.n65 16.5119
R349 source.n523 source.n488 13.1884
R350 source.n453 source.n418 13.1884
R351 source.n387 source.n352 13.1884
R352 source.n317 source.n282 13.1884
R353 source.n45 source.n10 13.1884
R354 source.n115 source.n80 13.1884
R355 source.n181 source.n146 13.1884
R356 source.n251 source.n216 13.1884
R357 source.n519 source.n518 12.8005
R358 source.n524 source.n486 12.8005
R359 source.n449 source.n448 12.8005
R360 source.n454 source.n416 12.8005
R361 source.n383 source.n382 12.8005
R362 source.n388 source.n350 12.8005
R363 source.n313 source.n312 12.8005
R364 source.n318 source.n280 12.8005
R365 source.n46 source.n8 12.8005
R366 source.n41 source.n12 12.8005
R367 source.n116 source.n78 12.8005
R368 source.n111 source.n82 12.8005
R369 source.n182 source.n144 12.8005
R370 source.n177 source.n148 12.8005
R371 source.n252 source.n214 12.8005
R372 source.n247 source.n218 12.8005
R373 source.n517 source.n490 12.0247
R374 source.n528 source.n527 12.0247
R375 source.n447 source.n420 12.0247
R376 source.n458 source.n457 12.0247
R377 source.n381 source.n354 12.0247
R378 source.n392 source.n391 12.0247
R379 source.n311 source.n284 12.0247
R380 source.n322 source.n321 12.0247
R381 source.n50 source.n49 12.0247
R382 source.n40 source.n13 12.0247
R383 source.n120 source.n119 12.0247
R384 source.n110 source.n83 12.0247
R385 source.n186 source.n185 12.0247
R386 source.n176 source.n149 12.0247
R387 source.n256 source.n255 12.0247
R388 source.n246 source.n219 12.0247
R389 source.n514 source.n513 11.249
R390 source.n531 source.n484 11.249
R391 source.n444 source.n443 11.249
R392 source.n461 source.n414 11.249
R393 source.n378 source.n377 11.249
R394 source.n395 source.n348 11.249
R395 source.n308 source.n307 11.249
R396 source.n325 source.n278 11.249
R397 source.n53 source.n6 11.249
R398 source.n37 source.n36 11.249
R399 source.n123 source.n76 11.249
R400 source.n107 source.n106 11.249
R401 source.n189 source.n142 11.249
R402 source.n173 source.n172 11.249
R403 source.n259 source.n212 11.249
R404 source.n243 source.n242 11.249
R405 source.n510 source.n492 10.4732
R406 source.n532 source.n482 10.4732
R407 source.n440 source.n422 10.4732
R408 source.n462 source.n412 10.4732
R409 source.n374 source.n356 10.4732
R410 source.n396 source.n346 10.4732
R411 source.n304 source.n286 10.4732
R412 source.n326 source.n276 10.4732
R413 source.n54 source.n4 10.4732
R414 source.n33 source.n15 10.4732
R415 source.n124 source.n74 10.4732
R416 source.n103 source.n85 10.4732
R417 source.n190 source.n140 10.4732
R418 source.n169 source.n151 10.4732
R419 source.n260 source.n210 10.4732
R420 source.n239 source.n221 10.4732
R421 source.n499 source.n498 10.2747
R422 source.n429 source.n428 10.2747
R423 source.n363 source.n362 10.2747
R424 source.n293 source.n292 10.2747
R425 source.n22 source.n21 10.2747
R426 source.n92 source.n91 10.2747
R427 source.n158 source.n157 10.2747
R428 source.n228 source.n227 10.2747
R429 source.n509 source.n494 9.69747
R430 source.n536 source.n535 9.69747
R431 source.n439 source.n424 9.69747
R432 source.n466 source.n465 9.69747
R433 source.n373 source.n358 9.69747
R434 source.n400 source.n399 9.69747
R435 source.n303 source.n288 9.69747
R436 source.n330 source.n329 9.69747
R437 source.n58 source.n57 9.69747
R438 source.n32 source.n17 9.69747
R439 source.n128 source.n127 9.69747
R440 source.n102 source.n87 9.69747
R441 source.n194 source.n193 9.69747
R442 source.n168 source.n153 9.69747
R443 source.n264 source.n263 9.69747
R444 source.n238 source.n223 9.69747
R445 source.n542 source.n541 9.45567
R446 source.n472 source.n471 9.45567
R447 source.n406 source.n405 9.45567
R448 source.n336 source.n335 9.45567
R449 source.n64 source.n63 9.45567
R450 source.n134 source.n133 9.45567
R451 source.n200 source.n199 9.45567
R452 source.n270 source.n269 9.45567
R453 source.n541 source.n540 9.3005
R454 source.n480 source.n479 9.3005
R455 source.n535 source.n534 9.3005
R456 source.n533 source.n532 9.3005
R457 source.n484 source.n483 9.3005
R458 source.n527 source.n526 9.3005
R459 source.n525 source.n524 9.3005
R460 source.n501 source.n500 9.3005
R461 source.n496 source.n495 9.3005
R462 source.n507 source.n506 9.3005
R463 source.n509 source.n508 9.3005
R464 source.n492 source.n491 9.3005
R465 source.n515 source.n514 9.3005
R466 source.n517 source.n516 9.3005
R467 source.n518 source.n487 9.3005
R468 source.n471 source.n470 9.3005
R469 source.n410 source.n409 9.3005
R470 source.n465 source.n464 9.3005
R471 source.n463 source.n462 9.3005
R472 source.n414 source.n413 9.3005
R473 source.n457 source.n456 9.3005
R474 source.n455 source.n454 9.3005
R475 source.n431 source.n430 9.3005
R476 source.n426 source.n425 9.3005
R477 source.n437 source.n436 9.3005
R478 source.n439 source.n438 9.3005
R479 source.n422 source.n421 9.3005
R480 source.n445 source.n444 9.3005
R481 source.n447 source.n446 9.3005
R482 source.n448 source.n417 9.3005
R483 source.n405 source.n404 9.3005
R484 source.n344 source.n343 9.3005
R485 source.n399 source.n398 9.3005
R486 source.n397 source.n396 9.3005
R487 source.n348 source.n347 9.3005
R488 source.n391 source.n390 9.3005
R489 source.n389 source.n388 9.3005
R490 source.n365 source.n364 9.3005
R491 source.n360 source.n359 9.3005
R492 source.n371 source.n370 9.3005
R493 source.n373 source.n372 9.3005
R494 source.n356 source.n355 9.3005
R495 source.n379 source.n378 9.3005
R496 source.n381 source.n380 9.3005
R497 source.n382 source.n351 9.3005
R498 source.n335 source.n334 9.3005
R499 source.n274 source.n273 9.3005
R500 source.n329 source.n328 9.3005
R501 source.n327 source.n326 9.3005
R502 source.n278 source.n277 9.3005
R503 source.n321 source.n320 9.3005
R504 source.n319 source.n318 9.3005
R505 source.n295 source.n294 9.3005
R506 source.n290 source.n289 9.3005
R507 source.n301 source.n300 9.3005
R508 source.n303 source.n302 9.3005
R509 source.n286 source.n285 9.3005
R510 source.n309 source.n308 9.3005
R511 source.n311 source.n310 9.3005
R512 source.n312 source.n281 9.3005
R513 source.n24 source.n23 9.3005
R514 source.n19 source.n18 9.3005
R515 source.n30 source.n29 9.3005
R516 source.n32 source.n31 9.3005
R517 source.n15 source.n14 9.3005
R518 source.n38 source.n37 9.3005
R519 source.n40 source.n39 9.3005
R520 source.n12 source.n9 9.3005
R521 source.n63 source.n62 9.3005
R522 source.n2 source.n1 9.3005
R523 source.n57 source.n56 9.3005
R524 source.n55 source.n54 9.3005
R525 source.n6 source.n5 9.3005
R526 source.n49 source.n48 9.3005
R527 source.n47 source.n46 9.3005
R528 source.n94 source.n93 9.3005
R529 source.n89 source.n88 9.3005
R530 source.n100 source.n99 9.3005
R531 source.n102 source.n101 9.3005
R532 source.n85 source.n84 9.3005
R533 source.n108 source.n107 9.3005
R534 source.n110 source.n109 9.3005
R535 source.n82 source.n79 9.3005
R536 source.n133 source.n132 9.3005
R537 source.n72 source.n71 9.3005
R538 source.n127 source.n126 9.3005
R539 source.n125 source.n124 9.3005
R540 source.n76 source.n75 9.3005
R541 source.n119 source.n118 9.3005
R542 source.n117 source.n116 9.3005
R543 source.n160 source.n159 9.3005
R544 source.n155 source.n154 9.3005
R545 source.n166 source.n165 9.3005
R546 source.n168 source.n167 9.3005
R547 source.n151 source.n150 9.3005
R548 source.n174 source.n173 9.3005
R549 source.n176 source.n175 9.3005
R550 source.n148 source.n145 9.3005
R551 source.n199 source.n198 9.3005
R552 source.n138 source.n137 9.3005
R553 source.n193 source.n192 9.3005
R554 source.n191 source.n190 9.3005
R555 source.n142 source.n141 9.3005
R556 source.n185 source.n184 9.3005
R557 source.n183 source.n182 9.3005
R558 source.n230 source.n229 9.3005
R559 source.n225 source.n224 9.3005
R560 source.n236 source.n235 9.3005
R561 source.n238 source.n237 9.3005
R562 source.n221 source.n220 9.3005
R563 source.n244 source.n243 9.3005
R564 source.n246 source.n245 9.3005
R565 source.n218 source.n215 9.3005
R566 source.n269 source.n268 9.3005
R567 source.n208 source.n207 9.3005
R568 source.n263 source.n262 9.3005
R569 source.n261 source.n260 9.3005
R570 source.n212 source.n211 9.3005
R571 source.n255 source.n254 9.3005
R572 source.n253 source.n252 9.3005
R573 source.n506 source.n505 8.92171
R574 source.n539 source.n480 8.92171
R575 source.n436 source.n435 8.92171
R576 source.n469 source.n410 8.92171
R577 source.n370 source.n369 8.92171
R578 source.n403 source.n344 8.92171
R579 source.n300 source.n299 8.92171
R580 source.n333 source.n274 8.92171
R581 source.n61 source.n2 8.92171
R582 source.n29 source.n28 8.92171
R583 source.n131 source.n72 8.92171
R584 source.n99 source.n98 8.92171
R585 source.n197 source.n138 8.92171
R586 source.n165 source.n164 8.92171
R587 source.n267 source.n208 8.92171
R588 source.n235 source.n234 8.92171
R589 source.n502 source.n496 8.14595
R590 source.n540 source.n478 8.14595
R591 source.n432 source.n426 8.14595
R592 source.n470 source.n408 8.14595
R593 source.n366 source.n360 8.14595
R594 source.n404 source.n342 8.14595
R595 source.n296 source.n290 8.14595
R596 source.n334 source.n272 8.14595
R597 source.n62 source.n0 8.14595
R598 source.n25 source.n19 8.14595
R599 source.n132 source.n70 8.14595
R600 source.n95 source.n89 8.14595
R601 source.n198 source.n136 8.14595
R602 source.n161 source.n155 8.14595
R603 source.n268 source.n206 8.14595
R604 source.n231 source.n225 8.14595
R605 source.n501 source.n498 7.3702
R606 source.n431 source.n428 7.3702
R607 source.n365 source.n362 7.3702
R608 source.n295 source.n292 7.3702
R609 source.n24 source.n21 7.3702
R610 source.n94 source.n91 7.3702
R611 source.n160 source.n157 7.3702
R612 source.n230 source.n227 7.3702
R613 source.n502 source.n501 5.81868
R614 source.n542 source.n478 5.81868
R615 source.n432 source.n431 5.81868
R616 source.n472 source.n408 5.81868
R617 source.n366 source.n365 5.81868
R618 source.n406 source.n342 5.81868
R619 source.n296 source.n295 5.81868
R620 source.n336 source.n272 5.81868
R621 source.n64 source.n0 5.81868
R622 source.n25 source.n24 5.81868
R623 source.n134 source.n70 5.81868
R624 source.n95 source.n94 5.81868
R625 source.n200 source.n136 5.81868
R626 source.n161 source.n160 5.81868
R627 source.n270 source.n206 5.81868
R628 source.n231 source.n230 5.81868
R629 source.n544 source.n543 5.7505
R630 source.n505 source.n496 5.04292
R631 source.n540 source.n539 5.04292
R632 source.n435 source.n426 5.04292
R633 source.n470 source.n469 5.04292
R634 source.n369 source.n360 5.04292
R635 source.n404 source.n403 5.04292
R636 source.n299 source.n290 5.04292
R637 source.n334 source.n333 5.04292
R638 source.n62 source.n61 5.04292
R639 source.n28 source.n19 5.04292
R640 source.n132 source.n131 5.04292
R641 source.n98 source.n89 5.04292
R642 source.n198 source.n197 5.04292
R643 source.n164 source.n155 5.04292
R644 source.n268 source.n267 5.04292
R645 source.n234 source.n225 5.04292
R646 source.n506 source.n494 4.26717
R647 source.n536 source.n480 4.26717
R648 source.n436 source.n424 4.26717
R649 source.n466 source.n410 4.26717
R650 source.n370 source.n358 4.26717
R651 source.n400 source.n344 4.26717
R652 source.n300 source.n288 4.26717
R653 source.n330 source.n274 4.26717
R654 source.n58 source.n2 4.26717
R655 source.n29 source.n17 4.26717
R656 source.n128 source.n72 4.26717
R657 source.n99 source.n87 4.26717
R658 source.n194 source.n138 4.26717
R659 source.n165 source.n153 4.26717
R660 source.n264 source.n208 4.26717
R661 source.n235 source.n223 4.26717
R662 source.n510 source.n509 3.49141
R663 source.n535 source.n482 3.49141
R664 source.n440 source.n439 3.49141
R665 source.n465 source.n412 3.49141
R666 source.n374 source.n373 3.49141
R667 source.n399 source.n346 3.49141
R668 source.n304 source.n303 3.49141
R669 source.n329 source.n276 3.49141
R670 source.n57 source.n4 3.49141
R671 source.n33 source.n32 3.49141
R672 source.n127 source.n74 3.49141
R673 source.n103 source.n102 3.49141
R674 source.n193 source.n140 3.49141
R675 source.n169 source.n168 3.49141
R676 source.n263 source.n210 3.49141
R677 source.n239 source.n238 3.49141
R678 source.n500 source.n499 2.84303
R679 source.n430 source.n429 2.84303
R680 source.n364 source.n363 2.84303
R681 source.n294 source.n293 2.84303
R682 source.n23 source.n22 2.84303
R683 source.n93 source.n92 2.84303
R684 source.n159 source.n158 2.84303
R685 source.n229 source.n228 2.84303
R686 source.n513 source.n492 2.71565
R687 source.n532 source.n531 2.71565
R688 source.n443 source.n422 2.71565
R689 source.n462 source.n461 2.71565
R690 source.n377 source.n356 2.71565
R691 source.n396 source.n395 2.71565
R692 source.n307 source.n286 2.71565
R693 source.n326 source.n325 2.71565
R694 source.n54 source.n53 2.71565
R695 source.n36 source.n15 2.71565
R696 source.n124 source.n123 2.71565
R697 source.n106 source.n85 2.71565
R698 source.n190 source.n189 2.71565
R699 source.n172 source.n151 2.71565
R700 source.n260 source.n259 2.71565
R701 source.n242 source.n221 2.71565
R702 source.n514 source.n490 1.93989
R703 source.n528 source.n484 1.93989
R704 source.n444 source.n420 1.93989
R705 source.n458 source.n414 1.93989
R706 source.n378 source.n354 1.93989
R707 source.n392 source.n348 1.93989
R708 source.n308 source.n284 1.93989
R709 source.n322 source.n278 1.93989
R710 source.n50 source.n6 1.93989
R711 source.n37 source.n13 1.93989
R712 source.n120 source.n76 1.93989
R713 source.n107 source.n83 1.93989
R714 source.n186 source.n142 1.93989
R715 source.n173 source.n149 1.93989
R716 source.n256 source.n212 1.93989
R717 source.n243 source.n219 1.93989
R718 source.n476 source.t10 1.6505
R719 source.n476 source.t11 1.6505
R720 source.n474 source.t20 1.6505
R721 source.n474 source.t19 1.6505
R722 source.n340 source.t9 1.6505
R723 source.n340 source.t8 1.6505
R724 source.n338 source.t5 1.6505
R725 source.n338 source.t23 1.6505
R726 source.n66 source.t22 1.6505
R727 source.n66 source.t0 1.6505
R728 source.n68 source.t2 1.6505
R729 source.n68 source.t6 1.6505
R730 source.n202 source.t12 1.6505
R731 source.n202 source.t16 1.6505
R732 source.n204 source.t13 1.6505
R733 source.n204 source.t14 1.6505
R734 source.n519 source.n517 1.16414
R735 source.n527 source.n486 1.16414
R736 source.n449 source.n447 1.16414
R737 source.n457 source.n416 1.16414
R738 source.n383 source.n381 1.16414
R739 source.n391 source.n350 1.16414
R740 source.n313 source.n311 1.16414
R741 source.n321 source.n280 1.16414
R742 source.n49 source.n8 1.16414
R743 source.n41 source.n40 1.16414
R744 source.n119 source.n78 1.16414
R745 source.n111 source.n110 1.16414
R746 source.n185 source.n144 1.16414
R747 source.n177 source.n176 1.16414
R748 source.n255 source.n214 1.16414
R749 source.n247 source.n246 1.16414
R750 source.n271 source.n205 0.974638
R751 source.n205 source.n203 0.974638
R752 source.n203 source.n201 0.974638
R753 source.n135 source.n69 0.974638
R754 source.n69 source.n67 0.974638
R755 source.n67 source.n65 0.974638
R756 source.n339 source.n337 0.974638
R757 source.n341 source.n339 0.974638
R758 source.n407 source.n341 0.974638
R759 source.n475 source.n473 0.974638
R760 source.n477 source.n475 0.974638
R761 source.n543 source.n477 0.974638
R762 source.n201 source.n135 0.470328
R763 source.n473 source.n407 0.470328
R764 source.n518 source.n488 0.388379
R765 source.n524 source.n523 0.388379
R766 source.n448 source.n418 0.388379
R767 source.n454 source.n453 0.388379
R768 source.n382 source.n352 0.388379
R769 source.n388 source.n387 0.388379
R770 source.n312 source.n282 0.388379
R771 source.n318 source.n317 0.388379
R772 source.n46 source.n45 0.388379
R773 source.n12 source.n10 0.388379
R774 source.n116 source.n115 0.388379
R775 source.n82 source.n80 0.388379
R776 source.n182 source.n181 0.388379
R777 source.n148 source.n146 0.388379
R778 source.n252 source.n251 0.388379
R779 source.n218 source.n216 0.388379
R780 source source.n544 0.188
R781 source.n500 source.n495 0.155672
R782 source.n507 source.n495 0.155672
R783 source.n508 source.n507 0.155672
R784 source.n508 source.n491 0.155672
R785 source.n515 source.n491 0.155672
R786 source.n516 source.n515 0.155672
R787 source.n516 source.n487 0.155672
R788 source.n525 source.n487 0.155672
R789 source.n526 source.n525 0.155672
R790 source.n526 source.n483 0.155672
R791 source.n533 source.n483 0.155672
R792 source.n534 source.n533 0.155672
R793 source.n534 source.n479 0.155672
R794 source.n541 source.n479 0.155672
R795 source.n430 source.n425 0.155672
R796 source.n437 source.n425 0.155672
R797 source.n438 source.n437 0.155672
R798 source.n438 source.n421 0.155672
R799 source.n445 source.n421 0.155672
R800 source.n446 source.n445 0.155672
R801 source.n446 source.n417 0.155672
R802 source.n455 source.n417 0.155672
R803 source.n456 source.n455 0.155672
R804 source.n456 source.n413 0.155672
R805 source.n463 source.n413 0.155672
R806 source.n464 source.n463 0.155672
R807 source.n464 source.n409 0.155672
R808 source.n471 source.n409 0.155672
R809 source.n364 source.n359 0.155672
R810 source.n371 source.n359 0.155672
R811 source.n372 source.n371 0.155672
R812 source.n372 source.n355 0.155672
R813 source.n379 source.n355 0.155672
R814 source.n380 source.n379 0.155672
R815 source.n380 source.n351 0.155672
R816 source.n389 source.n351 0.155672
R817 source.n390 source.n389 0.155672
R818 source.n390 source.n347 0.155672
R819 source.n397 source.n347 0.155672
R820 source.n398 source.n397 0.155672
R821 source.n398 source.n343 0.155672
R822 source.n405 source.n343 0.155672
R823 source.n294 source.n289 0.155672
R824 source.n301 source.n289 0.155672
R825 source.n302 source.n301 0.155672
R826 source.n302 source.n285 0.155672
R827 source.n309 source.n285 0.155672
R828 source.n310 source.n309 0.155672
R829 source.n310 source.n281 0.155672
R830 source.n319 source.n281 0.155672
R831 source.n320 source.n319 0.155672
R832 source.n320 source.n277 0.155672
R833 source.n327 source.n277 0.155672
R834 source.n328 source.n327 0.155672
R835 source.n328 source.n273 0.155672
R836 source.n335 source.n273 0.155672
R837 source.n63 source.n1 0.155672
R838 source.n56 source.n1 0.155672
R839 source.n56 source.n55 0.155672
R840 source.n55 source.n5 0.155672
R841 source.n48 source.n5 0.155672
R842 source.n48 source.n47 0.155672
R843 source.n47 source.n9 0.155672
R844 source.n39 source.n9 0.155672
R845 source.n39 source.n38 0.155672
R846 source.n38 source.n14 0.155672
R847 source.n31 source.n14 0.155672
R848 source.n31 source.n30 0.155672
R849 source.n30 source.n18 0.155672
R850 source.n23 source.n18 0.155672
R851 source.n133 source.n71 0.155672
R852 source.n126 source.n71 0.155672
R853 source.n126 source.n125 0.155672
R854 source.n125 source.n75 0.155672
R855 source.n118 source.n75 0.155672
R856 source.n118 source.n117 0.155672
R857 source.n117 source.n79 0.155672
R858 source.n109 source.n79 0.155672
R859 source.n109 source.n108 0.155672
R860 source.n108 source.n84 0.155672
R861 source.n101 source.n84 0.155672
R862 source.n101 source.n100 0.155672
R863 source.n100 source.n88 0.155672
R864 source.n93 source.n88 0.155672
R865 source.n199 source.n137 0.155672
R866 source.n192 source.n137 0.155672
R867 source.n192 source.n191 0.155672
R868 source.n191 source.n141 0.155672
R869 source.n184 source.n141 0.155672
R870 source.n184 source.n183 0.155672
R871 source.n183 source.n145 0.155672
R872 source.n175 source.n145 0.155672
R873 source.n175 source.n174 0.155672
R874 source.n174 source.n150 0.155672
R875 source.n167 source.n150 0.155672
R876 source.n167 source.n166 0.155672
R877 source.n166 source.n154 0.155672
R878 source.n159 source.n154 0.155672
R879 source.n269 source.n207 0.155672
R880 source.n262 source.n207 0.155672
R881 source.n262 source.n261 0.155672
R882 source.n261 source.n211 0.155672
R883 source.n254 source.n211 0.155672
R884 source.n254 source.n253 0.155672
R885 source.n253 source.n215 0.155672
R886 source.n245 source.n215 0.155672
R887 source.n245 source.n244 0.155672
R888 source.n244 source.n220 0.155672
R889 source.n237 source.n220 0.155672
R890 source.n237 source.n236 0.155672
R891 source.n236 source.n224 0.155672
R892 source.n229 source.n224 0.155672
R893 drain_right.n6 drain_right.n4 60.5266
R894 drain_right.n3 drain_right.n2 60.4713
R895 drain_right.n3 drain_right.n0 60.4713
R896 drain_right.n6 drain_right.n5 59.5527
R897 drain_right.n8 drain_right.n7 59.5527
R898 drain_right.n3 drain_right.n1 59.5525
R899 drain_right drain_right.n3 31.6845
R900 drain_right drain_right.n8 6.62735
R901 drain_right.n1 drain_right.t2 1.6505
R902 drain_right.n1 drain_right.t10 1.6505
R903 drain_right.n2 drain_right.t1 1.6505
R904 drain_right.n2 drain_right.t11 1.6505
R905 drain_right.n0 drain_right.t0 1.6505
R906 drain_right.n0 drain_right.t9 1.6505
R907 drain_right.n4 drain_right.t7 1.6505
R908 drain_right.n4 drain_right.t6 1.6505
R909 drain_right.n5 drain_right.t4 1.6505
R910 drain_right.n5 drain_right.t8 1.6505
R911 drain_right.n7 drain_right.t5 1.6505
R912 drain_right.n7 drain_right.t3 1.6505
R913 drain_right.n8 drain_right.n6 0.974638
R914 plus.n4 plus.t10 432
R915 plus.n20 plus.t7 432
R916 plus.n14 plus.t4 410.604
R917 plus.n12 plus.t8 410.604
R918 plus.n2 plus.t5 410.604
R919 plus.n7 plus.t6 410.604
R920 plus.n5 plus.t9 410.604
R921 plus.n30 plus.t11 410.604
R922 plus.n28 plus.t2 410.604
R923 plus.n18 plus.t0 410.604
R924 plus.n23 plus.t3 410.604
R925 plus.n21 plus.t1 410.604
R926 plus.n6 plus.n3 161.3
R927 plus.n11 plus.n10 161.3
R928 plus.n12 plus.n1 161.3
R929 plus.n13 plus.n0 161.3
R930 plus.n15 plus.n14 161.3
R931 plus.n22 plus.n19 161.3
R932 plus.n27 plus.n26 161.3
R933 plus.n28 plus.n17 161.3
R934 plus.n29 plus.n16 161.3
R935 plus.n31 plus.n30 161.3
R936 plus.n8 plus.n7 80.6037
R937 plus.n9 plus.n2 80.6037
R938 plus.n24 plus.n23 80.6037
R939 plus.n25 plus.n18 80.6037
R940 plus.n7 plus.n2 48.2005
R941 plus.n23 plus.n18 48.2005
R942 plus.n4 plus.n3 44.853
R943 plus.n20 plus.n19 44.853
R944 plus.n11 plus.n2 41.6278
R945 plus.n7 plus.n6 41.6278
R946 plus.n27 plus.n18 41.6278
R947 plus.n23 plus.n22 41.6278
R948 plus plus.n31 31.9081
R949 plus.n14 plus.n13 25.5611
R950 plus.n30 plus.n29 25.5611
R951 plus.n13 plus.n12 22.6399
R952 plus.n29 plus.n28 22.6399
R953 plus.n5 plus.n4 20.5405
R954 plus.n21 plus.n20 20.5405
R955 plus plus.n15 12.3452
R956 plus.n12 plus.n11 6.57323
R957 plus.n6 plus.n5 6.57323
R958 plus.n28 plus.n27 6.57323
R959 plus.n22 plus.n21 6.57323
R960 plus.n9 plus.n8 0.380177
R961 plus.n25 plus.n24 0.380177
R962 plus.n8 plus.n3 0.285035
R963 plus.n10 plus.n9 0.285035
R964 plus.n26 plus.n25 0.285035
R965 plus.n24 plus.n19 0.285035
R966 plus.n10 plus.n1 0.189894
R967 plus.n1 plus.n0 0.189894
R968 plus.n15 plus.n0 0.189894
R969 plus.n31 plus.n16 0.189894
R970 plus.n17 plus.n16 0.189894
R971 plus.n26 plus.n17 0.189894
R972 drain_left.n6 drain_left.n4 60.5268
R973 drain_left.n3 drain_left.n2 60.4713
R974 drain_left.n3 drain_left.n0 60.4713
R975 drain_left.n6 drain_left.n5 59.5527
R976 drain_left.n3 drain_left.n1 59.5525
R977 drain_left.n8 drain_left.n7 59.5525
R978 drain_left drain_left.n3 32.2378
R979 drain_left drain_left.n8 6.62735
R980 drain_left.n1 drain_left.t11 1.6505
R981 drain_left.n1 drain_left.t8 1.6505
R982 drain_left.n2 drain_left.t10 1.6505
R983 drain_left.n2 drain_left.t4 1.6505
R984 drain_left.n0 drain_left.t0 1.6505
R985 drain_left.n0 drain_left.t9 1.6505
R986 drain_left.n7 drain_left.t3 1.6505
R987 drain_left.n7 drain_left.t7 1.6505
R988 drain_left.n5 drain_left.t5 1.6505
R989 drain_left.n5 drain_left.t6 1.6505
R990 drain_left.n4 drain_left.t1 1.6505
R991 drain_left.n4 drain_left.t2 1.6505
R992 drain_left.n8 drain_left.n6 0.974638
C0 drain_left plus 8.678901f
C1 plus minus 6.00554f
C2 source drain_right 14.565901f
C3 drain_left drain_right 1.16185f
C4 drain_left source 14.5633f
C5 drain_right minus 8.452579f
C6 source minus 8.3985f
C7 plus drain_right 0.381869f
C8 plus source 8.412539f
C9 drain_left minus 0.17224f
C10 drain_right a_n2298_n3288# 6.31989f
C11 drain_left a_n2298_n3288# 6.64481f
C12 source a_n2298_n3288# 9.216989f
C13 minus a_n2298_n3288# 9.076711f
C14 plus a_n2298_n3288# 10.72991f
C15 drain_left.t0 a_n2298_n3288# 0.252971f
C16 drain_left.t9 a_n2298_n3288# 0.252971f
C17 drain_left.n0 a_n2298_n3288# 2.2571f
C18 drain_left.t11 a_n2298_n3288# 0.252971f
C19 drain_left.t8 a_n2298_n3288# 0.252971f
C20 drain_left.n1 a_n2298_n3288# 2.25105f
C21 drain_left.t10 a_n2298_n3288# 0.252971f
C22 drain_left.t4 a_n2298_n3288# 0.252971f
C23 drain_left.n2 a_n2298_n3288# 2.2571f
C24 drain_left.n3 a_n2298_n3288# 2.55552f
C25 drain_left.t1 a_n2298_n3288# 0.252971f
C26 drain_left.t2 a_n2298_n3288# 0.252971f
C27 drain_left.n4 a_n2298_n3288# 2.25753f
C28 drain_left.t5 a_n2298_n3288# 0.252971f
C29 drain_left.t6 a_n2298_n3288# 0.252971f
C30 drain_left.n5 a_n2298_n3288# 2.25106f
C31 drain_left.n6 a_n2298_n3288# 0.786974f
C32 drain_left.t3 a_n2298_n3288# 0.252971f
C33 drain_left.t7 a_n2298_n3288# 0.252971f
C34 drain_left.n7 a_n2298_n3288# 2.25105f
C35 drain_left.n8 a_n2298_n3288# 0.63057f
C36 plus.n0 a_n2298_n3288# 0.040251f
C37 plus.t4 a_n2298_n3288# 1.10185f
C38 plus.t8 a_n2298_n3288# 1.10185f
C39 plus.n1 a_n2298_n3288# 0.040251f
C40 plus.t5 a_n2298_n3288# 1.10185f
C41 plus.n2 a_n2298_n3288# 0.447003f
C42 plus.n3 a_n2298_n3288# 0.184783f
C43 plus.t6 a_n2298_n3288# 1.10185f
C44 plus.t9 a_n2298_n3288# 1.10185f
C45 plus.t10 a_n2298_n3288# 1.12355f
C46 plus.n4 a_n2298_n3288# 0.420292f
C47 plus.n5 a_n2298_n3288# 0.438895f
C48 plus.n6 a_n2298_n3288# 0.009134f
C49 plus.n7 a_n2298_n3288# 0.447003f
C50 plus.n8 a_n2298_n3288# 0.067043f
C51 plus.n9 a_n2298_n3288# 0.067043f
C52 plus.n10 a_n2298_n3288# 0.05371f
C53 plus.n11 a_n2298_n3288# 0.009134f
C54 plus.n12 a_n2298_n3288# 0.43576f
C55 plus.n13 a_n2298_n3288# 0.009134f
C56 plus.n14 a_n2298_n3288# 0.435139f
C57 plus.n15 a_n2298_n3288# 0.469616f
C58 plus.n16 a_n2298_n3288# 0.040251f
C59 plus.t11 a_n2298_n3288# 1.10185f
C60 plus.n17 a_n2298_n3288# 0.040251f
C61 plus.t2 a_n2298_n3288# 1.10185f
C62 plus.t0 a_n2298_n3288# 1.10185f
C63 plus.n18 a_n2298_n3288# 0.447003f
C64 plus.n19 a_n2298_n3288# 0.184783f
C65 plus.t3 a_n2298_n3288# 1.10185f
C66 plus.t7 a_n2298_n3288# 1.12355f
C67 plus.n20 a_n2298_n3288# 0.420292f
C68 plus.t1 a_n2298_n3288# 1.10185f
C69 plus.n21 a_n2298_n3288# 0.438895f
C70 plus.n22 a_n2298_n3288# 0.009134f
C71 plus.n23 a_n2298_n3288# 0.447003f
C72 plus.n24 a_n2298_n3288# 0.067043f
C73 plus.n25 a_n2298_n3288# 0.067043f
C74 plus.n26 a_n2298_n3288# 0.05371f
C75 plus.n27 a_n2298_n3288# 0.009134f
C76 plus.n28 a_n2298_n3288# 0.43576f
C77 plus.n29 a_n2298_n3288# 0.009134f
C78 plus.n30 a_n2298_n3288# 0.435139f
C79 plus.n31 a_n2298_n3288# 1.31137f
C80 drain_right.t0 a_n2298_n3288# 0.251928f
C81 drain_right.t9 a_n2298_n3288# 0.251928f
C82 drain_right.n0 a_n2298_n3288# 2.24779f
C83 drain_right.t2 a_n2298_n3288# 0.251928f
C84 drain_right.t10 a_n2298_n3288# 0.251928f
C85 drain_right.n1 a_n2298_n3288# 2.24177f
C86 drain_right.t1 a_n2298_n3288# 0.251928f
C87 drain_right.t11 a_n2298_n3288# 0.251928f
C88 drain_right.n2 a_n2298_n3288# 2.24779f
C89 drain_right.n3 a_n2298_n3288# 2.49029f
C90 drain_right.t7 a_n2298_n3288# 0.251928f
C91 drain_right.t6 a_n2298_n3288# 0.251928f
C92 drain_right.n4 a_n2298_n3288# 2.24821f
C93 drain_right.t4 a_n2298_n3288# 0.251928f
C94 drain_right.t8 a_n2298_n3288# 0.251928f
C95 drain_right.n5 a_n2298_n3288# 2.24178f
C96 drain_right.n6 a_n2298_n3288# 0.783738f
C97 drain_right.t5 a_n2298_n3288# 0.251928f
C98 drain_right.t3 a_n2298_n3288# 0.251928f
C99 drain_right.n7 a_n2298_n3288# 2.24178f
C100 drain_right.n8 a_n2298_n3288# 0.62796f
C101 source.n0 a_n2298_n3288# 0.028682f
C102 source.n1 a_n2298_n3288# 0.021653f
C103 source.n2 a_n2298_n3288# 0.011635f
C104 source.n3 a_n2298_n3288# 0.027502f
C105 source.n4 a_n2298_n3288# 0.01232f
C106 source.n5 a_n2298_n3288# 0.021653f
C107 source.n6 a_n2298_n3288# 0.011635f
C108 source.n7 a_n2298_n3288# 0.027502f
C109 source.n8 a_n2298_n3288# 0.01232f
C110 source.n9 a_n2298_n3288# 0.021653f
C111 source.n10 a_n2298_n3288# 0.011978f
C112 source.n11 a_n2298_n3288# 0.027502f
C113 source.n12 a_n2298_n3288# 0.011635f
C114 source.n13 a_n2298_n3288# 0.01232f
C115 source.n14 a_n2298_n3288# 0.021653f
C116 source.n15 a_n2298_n3288# 0.011635f
C117 source.n16 a_n2298_n3288# 0.027502f
C118 source.n17 a_n2298_n3288# 0.01232f
C119 source.n18 a_n2298_n3288# 0.021653f
C120 source.n19 a_n2298_n3288# 0.011635f
C121 source.n20 a_n2298_n3288# 0.020626f
C122 source.n21 a_n2298_n3288# 0.019441f
C123 source.t4 a_n2298_n3288# 0.046448f
C124 source.n22 a_n2298_n3288# 0.156114f
C125 source.n23 a_n2298_n3288# 1.09235f
C126 source.n24 a_n2298_n3288# 0.011635f
C127 source.n25 a_n2298_n3288# 0.01232f
C128 source.n26 a_n2298_n3288# 0.027502f
C129 source.n27 a_n2298_n3288# 0.027502f
C130 source.n28 a_n2298_n3288# 0.01232f
C131 source.n29 a_n2298_n3288# 0.011635f
C132 source.n30 a_n2298_n3288# 0.021653f
C133 source.n31 a_n2298_n3288# 0.021653f
C134 source.n32 a_n2298_n3288# 0.011635f
C135 source.n33 a_n2298_n3288# 0.01232f
C136 source.n34 a_n2298_n3288# 0.027502f
C137 source.n35 a_n2298_n3288# 0.027502f
C138 source.n36 a_n2298_n3288# 0.01232f
C139 source.n37 a_n2298_n3288# 0.011635f
C140 source.n38 a_n2298_n3288# 0.021653f
C141 source.n39 a_n2298_n3288# 0.021653f
C142 source.n40 a_n2298_n3288# 0.011635f
C143 source.n41 a_n2298_n3288# 0.01232f
C144 source.n42 a_n2298_n3288# 0.027502f
C145 source.n43 a_n2298_n3288# 0.027502f
C146 source.n44 a_n2298_n3288# 0.027502f
C147 source.n45 a_n2298_n3288# 0.011978f
C148 source.n46 a_n2298_n3288# 0.011635f
C149 source.n47 a_n2298_n3288# 0.021653f
C150 source.n48 a_n2298_n3288# 0.021653f
C151 source.n49 a_n2298_n3288# 0.011635f
C152 source.n50 a_n2298_n3288# 0.01232f
C153 source.n51 a_n2298_n3288# 0.027502f
C154 source.n52 a_n2298_n3288# 0.027502f
C155 source.n53 a_n2298_n3288# 0.01232f
C156 source.n54 a_n2298_n3288# 0.011635f
C157 source.n55 a_n2298_n3288# 0.021653f
C158 source.n56 a_n2298_n3288# 0.021653f
C159 source.n57 a_n2298_n3288# 0.011635f
C160 source.n58 a_n2298_n3288# 0.01232f
C161 source.n59 a_n2298_n3288# 0.027502f
C162 source.n60 a_n2298_n3288# 0.056436f
C163 source.n61 a_n2298_n3288# 0.01232f
C164 source.n62 a_n2298_n3288# 0.011635f
C165 source.n63 a_n2298_n3288# 0.0465f
C166 source.n64 a_n2298_n3288# 0.031147f
C167 source.n65 a_n2298_n3288# 0.920704f
C168 source.t22 a_n2298_n3288# 0.205329f
C169 source.t0 a_n2298_n3288# 0.205329f
C170 source.n66 a_n2298_n3288# 1.75803f
C171 source.n67 a_n2298_n3288# 0.357304f
C172 source.t2 a_n2298_n3288# 0.205329f
C173 source.t6 a_n2298_n3288# 0.205329f
C174 source.n68 a_n2298_n3288# 1.75803f
C175 source.n69 a_n2298_n3288# 0.357304f
C176 source.n70 a_n2298_n3288# 0.028682f
C177 source.n71 a_n2298_n3288# 0.021653f
C178 source.n72 a_n2298_n3288# 0.011635f
C179 source.n73 a_n2298_n3288# 0.027502f
C180 source.n74 a_n2298_n3288# 0.01232f
C181 source.n75 a_n2298_n3288# 0.021653f
C182 source.n76 a_n2298_n3288# 0.011635f
C183 source.n77 a_n2298_n3288# 0.027502f
C184 source.n78 a_n2298_n3288# 0.01232f
C185 source.n79 a_n2298_n3288# 0.021653f
C186 source.n80 a_n2298_n3288# 0.011978f
C187 source.n81 a_n2298_n3288# 0.027502f
C188 source.n82 a_n2298_n3288# 0.011635f
C189 source.n83 a_n2298_n3288# 0.01232f
C190 source.n84 a_n2298_n3288# 0.021653f
C191 source.n85 a_n2298_n3288# 0.011635f
C192 source.n86 a_n2298_n3288# 0.027502f
C193 source.n87 a_n2298_n3288# 0.01232f
C194 source.n88 a_n2298_n3288# 0.021653f
C195 source.n89 a_n2298_n3288# 0.011635f
C196 source.n90 a_n2298_n3288# 0.020626f
C197 source.n91 a_n2298_n3288# 0.019441f
C198 source.t1 a_n2298_n3288# 0.046448f
C199 source.n92 a_n2298_n3288# 0.156114f
C200 source.n93 a_n2298_n3288# 1.09235f
C201 source.n94 a_n2298_n3288# 0.011635f
C202 source.n95 a_n2298_n3288# 0.01232f
C203 source.n96 a_n2298_n3288# 0.027502f
C204 source.n97 a_n2298_n3288# 0.027502f
C205 source.n98 a_n2298_n3288# 0.01232f
C206 source.n99 a_n2298_n3288# 0.011635f
C207 source.n100 a_n2298_n3288# 0.021653f
C208 source.n101 a_n2298_n3288# 0.021653f
C209 source.n102 a_n2298_n3288# 0.011635f
C210 source.n103 a_n2298_n3288# 0.01232f
C211 source.n104 a_n2298_n3288# 0.027502f
C212 source.n105 a_n2298_n3288# 0.027502f
C213 source.n106 a_n2298_n3288# 0.01232f
C214 source.n107 a_n2298_n3288# 0.011635f
C215 source.n108 a_n2298_n3288# 0.021653f
C216 source.n109 a_n2298_n3288# 0.021653f
C217 source.n110 a_n2298_n3288# 0.011635f
C218 source.n111 a_n2298_n3288# 0.01232f
C219 source.n112 a_n2298_n3288# 0.027502f
C220 source.n113 a_n2298_n3288# 0.027502f
C221 source.n114 a_n2298_n3288# 0.027502f
C222 source.n115 a_n2298_n3288# 0.011978f
C223 source.n116 a_n2298_n3288# 0.011635f
C224 source.n117 a_n2298_n3288# 0.021653f
C225 source.n118 a_n2298_n3288# 0.021653f
C226 source.n119 a_n2298_n3288# 0.011635f
C227 source.n120 a_n2298_n3288# 0.01232f
C228 source.n121 a_n2298_n3288# 0.027502f
C229 source.n122 a_n2298_n3288# 0.027502f
C230 source.n123 a_n2298_n3288# 0.01232f
C231 source.n124 a_n2298_n3288# 0.011635f
C232 source.n125 a_n2298_n3288# 0.021653f
C233 source.n126 a_n2298_n3288# 0.021653f
C234 source.n127 a_n2298_n3288# 0.011635f
C235 source.n128 a_n2298_n3288# 0.01232f
C236 source.n129 a_n2298_n3288# 0.027502f
C237 source.n130 a_n2298_n3288# 0.056436f
C238 source.n131 a_n2298_n3288# 0.01232f
C239 source.n132 a_n2298_n3288# 0.011635f
C240 source.n133 a_n2298_n3288# 0.0465f
C241 source.n134 a_n2298_n3288# 0.031147f
C242 source.n135 a_n2298_n3288# 0.117239f
C243 source.n136 a_n2298_n3288# 0.028682f
C244 source.n137 a_n2298_n3288# 0.021653f
C245 source.n138 a_n2298_n3288# 0.011635f
C246 source.n139 a_n2298_n3288# 0.027502f
C247 source.n140 a_n2298_n3288# 0.01232f
C248 source.n141 a_n2298_n3288# 0.021653f
C249 source.n142 a_n2298_n3288# 0.011635f
C250 source.n143 a_n2298_n3288# 0.027502f
C251 source.n144 a_n2298_n3288# 0.01232f
C252 source.n145 a_n2298_n3288# 0.021653f
C253 source.n146 a_n2298_n3288# 0.011978f
C254 source.n147 a_n2298_n3288# 0.027502f
C255 source.n148 a_n2298_n3288# 0.011635f
C256 source.n149 a_n2298_n3288# 0.01232f
C257 source.n150 a_n2298_n3288# 0.021653f
C258 source.n151 a_n2298_n3288# 0.011635f
C259 source.n152 a_n2298_n3288# 0.027502f
C260 source.n153 a_n2298_n3288# 0.01232f
C261 source.n154 a_n2298_n3288# 0.021653f
C262 source.n155 a_n2298_n3288# 0.011635f
C263 source.n156 a_n2298_n3288# 0.020626f
C264 source.n157 a_n2298_n3288# 0.019441f
C265 source.t17 a_n2298_n3288# 0.046448f
C266 source.n158 a_n2298_n3288# 0.156114f
C267 source.n159 a_n2298_n3288# 1.09235f
C268 source.n160 a_n2298_n3288# 0.011635f
C269 source.n161 a_n2298_n3288# 0.01232f
C270 source.n162 a_n2298_n3288# 0.027502f
C271 source.n163 a_n2298_n3288# 0.027502f
C272 source.n164 a_n2298_n3288# 0.01232f
C273 source.n165 a_n2298_n3288# 0.011635f
C274 source.n166 a_n2298_n3288# 0.021653f
C275 source.n167 a_n2298_n3288# 0.021653f
C276 source.n168 a_n2298_n3288# 0.011635f
C277 source.n169 a_n2298_n3288# 0.01232f
C278 source.n170 a_n2298_n3288# 0.027502f
C279 source.n171 a_n2298_n3288# 0.027502f
C280 source.n172 a_n2298_n3288# 0.01232f
C281 source.n173 a_n2298_n3288# 0.011635f
C282 source.n174 a_n2298_n3288# 0.021653f
C283 source.n175 a_n2298_n3288# 0.021653f
C284 source.n176 a_n2298_n3288# 0.011635f
C285 source.n177 a_n2298_n3288# 0.01232f
C286 source.n178 a_n2298_n3288# 0.027502f
C287 source.n179 a_n2298_n3288# 0.027502f
C288 source.n180 a_n2298_n3288# 0.027502f
C289 source.n181 a_n2298_n3288# 0.011978f
C290 source.n182 a_n2298_n3288# 0.011635f
C291 source.n183 a_n2298_n3288# 0.021653f
C292 source.n184 a_n2298_n3288# 0.021653f
C293 source.n185 a_n2298_n3288# 0.011635f
C294 source.n186 a_n2298_n3288# 0.01232f
C295 source.n187 a_n2298_n3288# 0.027502f
C296 source.n188 a_n2298_n3288# 0.027502f
C297 source.n189 a_n2298_n3288# 0.01232f
C298 source.n190 a_n2298_n3288# 0.011635f
C299 source.n191 a_n2298_n3288# 0.021653f
C300 source.n192 a_n2298_n3288# 0.021653f
C301 source.n193 a_n2298_n3288# 0.011635f
C302 source.n194 a_n2298_n3288# 0.01232f
C303 source.n195 a_n2298_n3288# 0.027502f
C304 source.n196 a_n2298_n3288# 0.056436f
C305 source.n197 a_n2298_n3288# 0.01232f
C306 source.n198 a_n2298_n3288# 0.011635f
C307 source.n199 a_n2298_n3288# 0.0465f
C308 source.n200 a_n2298_n3288# 0.031147f
C309 source.n201 a_n2298_n3288# 0.117239f
C310 source.t12 a_n2298_n3288# 0.205329f
C311 source.t16 a_n2298_n3288# 0.205329f
C312 source.n202 a_n2298_n3288# 1.75803f
C313 source.n203 a_n2298_n3288# 0.357304f
C314 source.t13 a_n2298_n3288# 0.205329f
C315 source.t14 a_n2298_n3288# 0.205329f
C316 source.n204 a_n2298_n3288# 1.75803f
C317 source.n205 a_n2298_n3288# 0.357304f
C318 source.n206 a_n2298_n3288# 0.028682f
C319 source.n207 a_n2298_n3288# 0.021653f
C320 source.n208 a_n2298_n3288# 0.011635f
C321 source.n209 a_n2298_n3288# 0.027502f
C322 source.n210 a_n2298_n3288# 0.01232f
C323 source.n211 a_n2298_n3288# 0.021653f
C324 source.n212 a_n2298_n3288# 0.011635f
C325 source.n213 a_n2298_n3288# 0.027502f
C326 source.n214 a_n2298_n3288# 0.01232f
C327 source.n215 a_n2298_n3288# 0.021653f
C328 source.n216 a_n2298_n3288# 0.011978f
C329 source.n217 a_n2298_n3288# 0.027502f
C330 source.n218 a_n2298_n3288# 0.011635f
C331 source.n219 a_n2298_n3288# 0.01232f
C332 source.n220 a_n2298_n3288# 0.021653f
C333 source.n221 a_n2298_n3288# 0.011635f
C334 source.n222 a_n2298_n3288# 0.027502f
C335 source.n223 a_n2298_n3288# 0.01232f
C336 source.n224 a_n2298_n3288# 0.021653f
C337 source.n225 a_n2298_n3288# 0.011635f
C338 source.n226 a_n2298_n3288# 0.020626f
C339 source.n227 a_n2298_n3288# 0.019441f
C340 source.t15 a_n2298_n3288# 0.046448f
C341 source.n228 a_n2298_n3288# 0.156114f
C342 source.n229 a_n2298_n3288# 1.09235f
C343 source.n230 a_n2298_n3288# 0.011635f
C344 source.n231 a_n2298_n3288# 0.01232f
C345 source.n232 a_n2298_n3288# 0.027502f
C346 source.n233 a_n2298_n3288# 0.027502f
C347 source.n234 a_n2298_n3288# 0.01232f
C348 source.n235 a_n2298_n3288# 0.011635f
C349 source.n236 a_n2298_n3288# 0.021653f
C350 source.n237 a_n2298_n3288# 0.021653f
C351 source.n238 a_n2298_n3288# 0.011635f
C352 source.n239 a_n2298_n3288# 0.01232f
C353 source.n240 a_n2298_n3288# 0.027502f
C354 source.n241 a_n2298_n3288# 0.027502f
C355 source.n242 a_n2298_n3288# 0.01232f
C356 source.n243 a_n2298_n3288# 0.011635f
C357 source.n244 a_n2298_n3288# 0.021653f
C358 source.n245 a_n2298_n3288# 0.021653f
C359 source.n246 a_n2298_n3288# 0.011635f
C360 source.n247 a_n2298_n3288# 0.01232f
C361 source.n248 a_n2298_n3288# 0.027502f
C362 source.n249 a_n2298_n3288# 0.027502f
C363 source.n250 a_n2298_n3288# 0.027502f
C364 source.n251 a_n2298_n3288# 0.011978f
C365 source.n252 a_n2298_n3288# 0.011635f
C366 source.n253 a_n2298_n3288# 0.021653f
C367 source.n254 a_n2298_n3288# 0.021653f
C368 source.n255 a_n2298_n3288# 0.011635f
C369 source.n256 a_n2298_n3288# 0.01232f
C370 source.n257 a_n2298_n3288# 0.027502f
C371 source.n258 a_n2298_n3288# 0.027502f
C372 source.n259 a_n2298_n3288# 0.01232f
C373 source.n260 a_n2298_n3288# 0.011635f
C374 source.n261 a_n2298_n3288# 0.021653f
C375 source.n262 a_n2298_n3288# 0.021653f
C376 source.n263 a_n2298_n3288# 0.011635f
C377 source.n264 a_n2298_n3288# 0.01232f
C378 source.n265 a_n2298_n3288# 0.027502f
C379 source.n266 a_n2298_n3288# 0.056436f
C380 source.n267 a_n2298_n3288# 0.01232f
C381 source.n268 a_n2298_n3288# 0.011635f
C382 source.n269 a_n2298_n3288# 0.0465f
C383 source.n270 a_n2298_n3288# 0.031147f
C384 source.n271 a_n2298_n3288# 1.27204f
C385 source.n272 a_n2298_n3288# 0.028682f
C386 source.n273 a_n2298_n3288# 0.021653f
C387 source.n274 a_n2298_n3288# 0.011635f
C388 source.n275 a_n2298_n3288# 0.027502f
C389 source.n276 a_n2298_n3288# 0.01232f
C390 source.n277 a_n2298_n3288# 0.021653f
C391 source.n278 a_n2298_n3288# 0.011635f
C392 source.n279 a_n2298_n3288# 0.027502f
C393 source.n280 a_n2298_n3288# 0.01232f
C394 source.n281 a_n2298_n3288# 0.021653f
C395 source.n282 a_n2298_n3288# 0.011978f
C396 source.n283 a_n2298_n3288# 0.027502f
C397 source.n284 a_n2298_n3288# 0.01232f
C398 source.n285 a_n2298_n3288# 0.021653f
C399 source.n286 a_n2298_n3288# 0.011635f
C400 source.n287 a_n2298_n3288# 0.027502f
C401 source.n288 a_n2298_n3288# 0.01232f
C402 source.n289 a_n2298_n3288# 0.021653f
C403 source.n290 a_n2298_n3288# 0.011635f
C404 source.n291 a_n2298_n3288# 0.020626f
C405 source.n292 a_n2298_n3288# 0.019441f
C406 source.t3 a_n2298_n3288# 0.046448f
C407 source.n293 a_n2298_n3288# 0.156114f
C408 source.n294 a_n2298_n3288# 1.09235f
C409 source.n295 a_n2298_n3288# 0.011635f
C410 source.n296 a_n2298_n3288# 0.01232f
C411 source.n297 a_n2298_n3288# 0.027502f
C412 source.n298 a_n2298_n3288# 0.027502f
C413 source.n299 a_n2298_n3288# 0.01232f
C414 source.n300 a_n2298_n3288# 0.011635f
C415 source.n301 a_n2298_n3288# 0.021653f
C416 source.n302 a_n2298_n3288# 0.021653f
C417 source.n303 a_n2298_n3288# 0.011635f
C418 source.n304 a_n2298_n3288# 0.01232f
C419 source.n305 a_n2298_n3288# 0.027502f
C420 source.n306 a_n2298_n3288# 0.027502f
C421 source.n307 a_n2298_n3288# 0.01232f
C422 source.n308 a_n2298_n3288# 0.011635f
C423 source.n309 a_n2298_n3288# 0.021653f
C424 source.n310 a_n2298_n3288# 0.021653f
C425 source.n311 a_n2298_n3288# 0.011635f
C426 source.n312 a_n2298_n3288# 0.011635f
C427 source.n313 a_n2298_n3288# 0.01232f
C428 source.n314 a_n2298_n3288# 0.027502f
C429 source.n315 a_n2298_n3288# 0.027502f
C430 source.n316 a_n2298_n3288# 0.027502f
C431 source.n317 a_n2298_n3288# 0.011978f
C432 source.n318 a_n2298_n3288# 0.011635f
C433 source.n319 a_n2298_n3288# 0.021653f
C434 source.n320 a_n2298_n3288# 0.021653f
C435 source.n321 a_n2298_n3288# 0.011635f
C436 source.n322 a_n2298_n3288# 0.01232f
C437 source.n323 a_n2298_n3288# 0.027502f
C438 source.n324 a_n2298_n3288# 0.027502f
C439 source.n325 a_n2298_n3288# 0.01232f
C440 source.n326 a_n2298_n3288# 0.011635f
C441 source.n327 a_n2298_n3288# 0.021653f
C442 source.n328 a_n2298_n3288# 0.021653f
C443 source.n329 a_n2298_n3288# 0.011635f
C444 source.n330 a_n2298_n3288# 0.01232f
C445 source.n331 a_n2298_n3288# 0.027502f
C446 source.n332 a_n2298_n3288# 0.056436f
C447 source.n333 a_n2298_n3288# 0.01232f
C448 source.n334 a_n2298_n3288# 0.011635f
C449 source.n335 a_n2298_n3288# 0.0465f
C450 source.n336 a_n2298_n3288# 0.031147f
C451 source.n337 a_n2298_n3288# 1.27204f
C452 source.t5 a_n2298_n3288# 0.205329f
C453 source.t23 a_n2298_n3288# 0.205329f
C454 source.n338 a_n2298_n3288# 1.75802f
C455 source.n339 a_n2298_n3288# 0.357315f
C456 source.t9 a_n2298_n3288# 0.205329f
C457 source.t8 a_n2298_n3288# 0.205329f
C458 source.n340 a_n2298_n3288# 1.75802f
C459 source.n341 a_n2298_n3288# 0.357315f
C460 source.n342 a_n2298_n3288# 0.028682f
C461 source.n343 a_n2298_n3288# 0.021653f
C462 source.n344 a_n2298_n3288# 0.011635f
C463 source.n345 a_n2298_n3288# 0.027502f
C464 source.n346 a_n2298_n3288# 0.01232f
C465 source.n347 a_n2298_n3288# 0.021653f
C466 source.n348 a_n2298_n3288# 0.011635f
C467 source.n349 a_n2298_n3288# 0.027502f
C468 source.n350 a_n2298_n3288# 0.01232f
C469 source.n351 a_n2298_n3288# 0.021653f
C470 source.n352 a_n2298_n3288# 0.011978f
C471 source.n353 a_n2298_n3288# 0.027502f
C472 source.n354 a_n2298_n3288# 0.01232f
C473 source.n355 a_n2298_n3288# 0.021653f
C474 source.n356 a_n2298_n3288# 0.011635f
C475 source.n357 a_n2298_n3288# 0.027502f
C476 source.n358 a_n2298_n3288# 0.01232f
C477 source.n359 a_n2298_n3288# 0.021653f
C478 source.n360 a_n2298_n3288# 0.011635f
C479 source.n361 a_n2298_n3288# 0.020626f
C480 source.n362 a_n2298_n3288# 0.019441f
C481 source.t7 a_n2298_n3288# 0.046448f
C482 source.n363 a_n2298_n3288# 0.156114f
C483 source.n364 a_n2298_n3288# 1.09235f
C484 source.n365 a_n2298_n3288# 0.011635f
C485 source.n366 a_n2298_n3288# 0.01232f
C486 source.n367 a_n2298_n3288# 0.027502f
C487 source.n368 a_n2298_n3288# 0.027502f
C488 source.n369 a_n2298_n3288# 0.01232f
C489 source.n370 a_n2298_n3288# 0.011635f
C490 source.n371 a_n2298_n3288# 0.021653f
C491 source.n372 a_n2298_n3288# 0.021653f
C492 source.n373 a_n2298_n3288# 0.011635f
C493 source.n374 a_n2298_n3288# 0.01232f
C494 source.n375 a_n2298_n3288# 0.027502f
C495 source.n376 a_n2298_n3288# 0.027502f
C496 source.n377 a_n2298_n3288# 0.01232f
C497 source.n378 a_n2298_n3288# 0.011635f
C498 source.n379 a_n2298_n3288# 0.021653f
C499 source.n380 a_n2298_n3288# 0.021653f
C500 source.n381 a_n2298_n3288# 0.011635f
C501 source.n382 a_n2298_n3288# 0.011635f
C502 source.n383 a_n2298_n3288# 0.01232f
C503 source.n384 a_n2298_n3288# 0.027502f
C504 source.n385 a_n2298_n3288# 0.027502f
C505 source.n386 a_n2298_n3288# 0.027502f
C506 source.n387 a_n2298_n3288# 0.011978f
C507 source.n388 a_n2298_n3288# 0.011635f
C508 source.n389 a_n2298_n3288# 0.021653f
C509 source.n390 a_n2298_n3288# 0.021653f
C510 source.n391 a_n2298_n3288# 0.011635f
C511 source.n392 a_n2298_n3288# 0.01232f
C512 source.n393 a_n2298_n3288# 0.027502f
C513 source.n394 a_n2298_n3288# 0.027502f
C514 source.n395 a_n2298_n3288# 0.01232f
C515 source.n396 a_n2298_n3288# 0.011635f
C516 source.n397 a_n2298_n3288# 0.021653f
C517 source.n398 a_n2298_n3288# 0.021653f
C518 source.n399 a_n2298_n3288# 0.011635f
C519 source.n400 a_n2298_n3288# 0.01232f
C520 source.n401 a_n2298_n3288# 0.027502f
C521 source.n402 a_n2298_n3288# 0.056436f
C522 source.n403 a_n2298_n3288# 0.01232f
C523 source.n404 a_n2298_n3288# 0.011635f
C524 source.n405 a_n2298_n3288# 0.0465f
C525 source.n406 a_n2298_n3288# 0.031147f
C526 source.n407 a_n2298_n3288# 0.117239f
C527 source.n408 a_n2298_n3288# 0.028682f
C528 source.n409 a_n2298_n3288# 0.021653f
C529 source.n410 a_n2298_n3288# 0.011635f
C530 source.n411 a_n2298_n3288# 0.027502f
C531 source.n412 a_n2298_n3288# 0.01232f
C532 source.n413 a_n2298_n3288# 0.021653f
C533 source.n414 a_n2298_n3288# 0.011635f
C534 source.n415 a_n2298_n3288# 0.027502f
C535 source.n416 a_n2298_n3288# 0.01232f
C536 source.n417 a_n2298_n3288# 0.021653f
C537 source.n418 a_n2298_n3288# 0.011978f
C538 source.n419 a_n2298_n3288# 0.027502f
C539 source.n420 a_n2298_n3288# 0.01232f
C540 source.n421 a_n2298_n3288# 0.021653f
C541 source.n422 a_n2298_n3288# 0.011635f
C542 source.n423 a_n2298_n3288# 0.027502f
C543 source.n424 a_n2298_n3288# 0.01232f
C544 source.n425 a_n2298_n3288# 0.021653f
C545 source.n426 a_n2298_n3288# 0.011635f
C546 source.n427 a_n2298_n3288# 0.020626f
C547 source.n428 a_n2298_n3288# 0.019441f
C548 source.t21 a_n2298_n3288# 0.046448f
C549 source.n429 a_n2298_n3288# 0.156114f
C550 source.n430 a_n2298_n3288# 1.09235f
C551 source.n431 a_n2298_n3288# 0.011635f
C552 source.n432 a_n2298_n3288# 0.01232f
C553 source.n433 a_n2298_n3288# 0.027502f
C554 source.n434 a_n2298_n3288# 0.027502f
C555 source.n435 a_n2298_n3288# 0.01232f
C556 source.n436 a_n2298_n3288# 0.011635f
C557 source.n437 a_n2298_n3288# 0.021653f
C558 source.n438 a_n2298_n3288# 0.021653f
C559 source.n439 a_n2298_n3288# 0.011635f
C560 source.n440 a_n2298_n3288# 0.01232f
C561 source.n441 a_n2298_n3288# 0.027502f
C562 source.n442 a_n2298_n3288# 0.027502f
C563 source.n443 a_n2298_n3288# 0.01232f
C564 source.n444 a_n2298_n3288# 0.011635f
C565 source.n445 a_n2298_n3288# 0.021653f
C566 source.n446 a_n2298_n3288# 0.021653f
C567 source.n447 a_n2298_n3288# 0.011635f
C568 source.n448 a_n2298_n3288# 0.011635f
C569 source.n449 a_n2298_n3288# 0.01232f
C570 source.n450 a_n2298_n3288# 0.027502f
C571 source.n451 a_n2298_n3288# 0.027502f
C572 source.n452 a_n2298_n3288# 0.027502f
C573 source.n453 a_n2298_n3288# 0.011978f
C574 source.n454 a_n2298_n3288# 0.011635f
C575 source.n455 a_n2298_n3288# 0.021653f
C576 source.n456 a_n2298_n3288# 0.021653f
C577 source.n457 a_n2298_n3288# 0.011635f
C578 source.n458 a_n2298_n3288# 0.01232f
C579 source.n459 a_n2298_n3288# 0.027502f
C580 source.n460 a_n2298_n3288# 0.027502f
C581 source.n461 a_n2298_n3288# 0.01232f
C582 source.n462 a_n2298_n3288# 0.011635f
C583 source.n463 a_n2298_n3288# 0.021653f
C584 source.n464 a_n2298_n3288# 0.021653f
C585 source.n465 a_n2298_n3288# 0.011635f
C586 source.n466 a_n2298_n3288# 0.01232f
C587 source.n467 a_n2298_n3288# 0.027502f
C588 source.n468 a_n2298_n3288# 0.056436f
C589 source.n469 a_n2298_n3288# 0.01232f
C590 source.n470 a_n2298_n3288# 0.011635f
C591 source.n471 a_n2298_n3288# 0.0465f
C592 source.n472 a_n2298_n3288# 0.031147f
C593 source.n473 a_n2298_n3288# 0.117239f
C594 source.t20 a_n2298_n3288# 0.205329f
C595 source.t19 a_n2298_n3288# 0.205329f
C596 source.n474 a_n2298_n3288# 1.75802f
C597 source.n475 a_n2298_n3288# 0.357315f
C598 source.t10 a_n2298_n3288# 0.205329f
C599 source.t11 a_n2298_n3288# 0.205329f
C600 source.n476 a_n2298_n3288# 1.75802f
C601 source.n477 a_n2298_n3288# 0.357315f
C602 source.n478 a_n2298_n3288# 0.028682f
C603 source.n479 a_n2298_n3288# 0.021653f
C604 source.n480 a_n2298_n3288# 0.011635f
C605 source.n481 a_n2298_n3288# 0.027502f
C606 source.n482 a_n2298_n3288# 0.01232f
C607 source.n483 a_n2298_n3288# 0.021653f
C608 source.n484 a_n2298_n3288# 0.011635f
C609 source.n485 a_n2298_n3288# 0.027502f
C610 source.n486 a_n2298_n3288# 0.01232f
C611 source.n487 a_n2298_n3288# 0.021653f
C612 source.n488 a_n2298_n3288# 0.011978f
C613 source.n489 a_n2298_n3288# 0.027502f
C614 source.n490 a_n2298_n3288# 0.01232f
C615 source.n491 a_n2298_n3288# 0.021653f
C616 source.n492 a_n2298_n3288# 0.011635f
C617 source.n493 a_n2298_n3288# 0.027502f
C618 source.n494 a_n2298_n3288# 0.01232f
C619 source.n495 a_n2298_n3288# 0.021653f
C620 source.n496 a_n2298_n3288# 0.011635f
C621 source.n497 a_n2298_n3288# 0.020626f
C622 source.n498 a_n2298_n3288# 0.019441f
C623 source.t18 a_n2298_n3288# 0.046448f
C624 source.n499 a_n2298_n3288# 0.156114f
C625 source.n500 a_n2298_n3288# 1.09235f
C626 source.n501 a_n2298_n3288# 0.011635f
C627 source.n502 a_n2298_n3288# 0.01232f
C628 source.n503 a_n2298_n3288# 0.027502f
C629 source.n504 a_n2298_n3288# 0.027502f
C630 source.n505 a_n2298_n3288# 0.01232f
C631 source.n506 a_n2298_n3288# 0.011635f
C632 source.n507 a_n2298_n3288# 0.021653f
C633 source.n508 a_n2298_n3288# 0.021653f
C634 source.n509 a_n2298_n3288# 0.011635f
C635 source.n510 a_n2298_n3288# 0.01232f
C636 source.n511 a_n2298_n3288# 0.027502f
C637 source.n512 a_n2298_n3288# 0.027502f
C638 source.n513 a_n2298_n3288# 0.01232f
C639 source.n514 a_n2298_n3288# 0.011635f
C640 source.n515 a_n2298_n3288# 0.021653f
C641 source.n516 a_n2298_n3288# 0.021653f
C642 source.n517 a_n2298_n3288# 0.011635f
C643 source.n518 a_n2298_n3288# 0.011635f
C644 source.n519 a_n2298_n3288# 0.01232f
C645 source.n520 a_n2298_n3288# 0.027502f
C646 source.n521 a_n2298_n3288# 0.027502f
C647 source.n522 a_n2298_n3288# 0.027502f
C648 source.n523 a_n2298_n3288# 0.011978f
C649 source.n524 a_n2298_n3288# 0.011635f
C650 source.n525 a_n2298_n3288# 0.021653f
C651 source.n526 a_n2298_n3288# 0.021653f
C652 source.n527 a_n2298_n3288# 0.011635f
C653 source.n528 a_n2298_n3288# 0.01232f
C654 source.n529 a_n2298_n3288# 0.027502f
C655 source.n530 a_n2298_n3288# 0.027502f
C656 source.n531 a_n2298_n3288# 0.01232f
C657 source.n532 a_n2298_n3288# 0.011635f
C658 source.n533 a_n2298_n3288# 0.021653f
C659 source.n534 a_n2298_n3288# 0.021653f
C660 source.n535 a_n2298_n3288# 0.011635f
C661 source.n536 a_n2298_n3288# 0.01232f
C662 source.n537 a_n2298_n3288# 0.027502f
C663 source.n538 a_n2298_n3288# 0.056436f
C664 source.n539 a_n2298_n3288# 0.01232f
C665 source.n540 a_n2298_n3288# 0.011635f
C666 source.n541 a_n2298_n3288# 0.0465f
C667 source.n542 a_n2298_n3288# 0.031147f
C668 source.n543 a_n2298_n3288# 0.263169f
C669 source.n544 a_n2298_n3288# 1.3756f
C670 minus.n0 a_n2298_n3288# 0.039762f
C671 minus.n1 a_n2298_n3288# 0.009023f
C672 minus.t8 a_n2298_n3288# 1.08848f
C673 minus.n2 a_n2298_n3288# 0.066229f
C674 minus.t4 a_n2298_n3288# 1.08848f
C675 minus.n3 a_n2298_n3288# 0.433568f
C676 minus.t5 a_n2298_n3288# 1.10991f
C677 minus.n4 a_n2298_n3288# 0.41519f
C678 minus.n5 a_n2298_n3288# 0.18254f
C679 minus.n6 a_n2298_n3288# 0.009023f
C680 minus.t3 a_n2298_n3288# 1.08848f
C681 minus.n7 a_n2298_n3288# 0.441577f
C682 minus.t7 a_n2298_n3288# 1.08848f
C683 minus.n8 a_n2298_n3288# 0.441577f
C684 minus.n9 a_n2298_n3288# 0.066229f
C685 minus.n10 a_n2298_n3288# 0.053058f
C686 minus.n11 a_n2298_n3288# 0.039762f
C687 minus.n12 a_n2298_n3288# 0.43047f
C688 minus.n13 a_n2298_n3288# 0.009023f
C689 minus.t6 a_n2298_n3288# 1.08848f
C690 minus.n14 a_n2298_n3288# 0.429857f
C691 minus.n15 a_n2298_n3288# 1.52276f
C692 minus.n16 a_n2298_n3288# 0.039762f
C693 minus.n17 a_n2298_n3288# 0.009023f
C694 minus.n18 a_n2298_n3288# 0.066229f
C695 minus.t2 a_n2298_n3288# 1.08848f
C696 minus.n19 a_n2298_n3288# 0.433568f
C697 minus.t11 a_n2298_n3288# 1.10991f
C698 minus.n20 a_n2298_n3288# 0.41519f
C699 minus.n21 a_n2298_n3288# 0.18254f
C700 minus.n22 a_n2298_n3288# 0.009023f
C701 minus.t9 a_n2298_n3288# 1.08848f
C702 minus.n23 a_n2298_n3288# 0.441577f
C703 minus.t1 a_n2298_n3288# 1.08848f
C704 minus.n24 a_n2298_n3288# 0.441577f
C705 minus.n25 a_n2298_n3288# 0.066229f
C706 minus.n26 a_n2298_n3288# 0.053058f
C707 minus.n27 a_n2298_n3288# 0.039762f
C708 minus.t10 a_n2298_n3288# 1.08848f
C709 minus.n28 a_n2298_n3288# 0.43047f
C710 minus.n29 a_n2298_n3288# 0.009023f
C711 minus.t0 a_n2298_n3288# 1.08848f
C712 minus.n30 a_n2298_n3288# 0.429857f
C713 minus.n31 a_n2298_n3288# 0.278635f
C714 minus.n32 a_n2298_n3288# 1.83412f
.ends

