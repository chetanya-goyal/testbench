* NGSPICE file created from diffpair323.ext - technology: sky130A

.subckt diffpair323 minus drain_right drain_left source plus
X0 drain_left plus source a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X1 a_n1366_n2688# a_n1366_n2688# a_n1366_n2688# a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=34.2 ps=151.6 w=9 l=0.15
X2 a_n1366_n2688# a_n1366_n2688# a_n1366_n2688# a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X3 source plus drain_left a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X4 a_n1366_n2688# a_n1366_n2688# a_n1366_n2688# a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X5 drain_left plus source a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X6 drain_right minus source a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X7 a_n1366_n2688# a_n1366_n2688# a_n1366_n2688# a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X8 source minus drain_right a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X9 source plus drain_left a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X10 drain_right minus source a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X11 source minus drain_right a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X12 source minus drain_right a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X13 source plus drain_left a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X14 drain_right minus source a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X15 drain_left plus source a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X16 drain_right minus source a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X17 source plus drain_left a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X18 drain_left plus source a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X19 source minus drain_right a_n1366_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
.ends

