* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t19 plus.t0 drain_left.t5 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X1 source.t18 plus.t1 drain_left.t1 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X2 drain_right.t9 minus.t0 source.t5 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X3 source.t4 minus.t1 drain_right.t8 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X4 a_n1412_n1088# a_n1412_n1088# a_n1412_n1088# a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.25
X5 source.t1 minus.t2 drain_right.t7 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X6 drain_right.t6 minus.t3 source.t9 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X7 drain_right.t5 minus.t4 source.t8 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X8 drain_left.t7 plus.t2 source.t17 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X9 source.t16 plus.t3 drain_left.t0 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X10 drain_left.t2 plus.t4 source.t15 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X11 drain_left.t9 plus.t5 source.t14 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X12 drain_left.t8 plus.t6 source.t13 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X13 a_n1412_n1088# a_n1412_n1088# a_n1412_n1088# a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X14 a_n1412_n1088# a_n1412_n1088# a_n1412_n1088# a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X15 drain_left.t3 plus.t7 source.t12 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X16 drain_right.t4 minus.t5 source.t7 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X17 drain_right.t3 minus.t6 source.t3 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X18 drain_left.t4 plus.t8 source.t11 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X19 source.t10 plus.t9 drain_left.t6 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X20 drain_right.t2 minus.t7 source.t6 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X21 a_n1412_n1088# a_n1412_n1088# a_n1412_n1088# a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X22 source.t0 minus.t8 drain_right.t1 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X23 source.t2 minus.t9 drain_right.t0 a_n1412_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
R0 plus.n2 plus.t2 281.606
R1 plus.n8 plus.t4 281.606
R2 plus.n12 plus.t7 281.606
R3 plus.n18 plus.t6 281.606
R4 plus.n1 plus.t1 221.72
R5 plus.n5 plus.t5 221.72
R6 plus.n7 plus.t0 221.72
R7 plus.n11 plus.t3 221.72
R8 plus.n15 plus.t8 221.72
R9 plus.n17 plus.t9 221.72
R10 plus.n3 plus.n2 161.489
R11 plus.n13 plus.n12 161.489
R12 plus.n4 plus.n3 161.3
R13 plus.n6 plus.n0 161.3
R14 plus.n9 plus.n8 161.3
R15 plus.n14 plus.n13 161.3
R16 plus.n16 plus.n10 161.3
R17 plus.n19 plus.n18 161.3
R18 plus.n4 plus.n1 48.2005
R19 plus.n7 plus.n6 48.2005
R20 plus.n17 plus.n16 48.2005
R21 plus.n14 plus.n11 48.2005
R22 plus.n5 plus.n4 36.5157
R23 plus.n6 plus.n5 36.5157
R24 plus.n16 plus.n15 36.5157
R25 plus.n15 plus.n14 36.5157
R26 plus.n2 plus.n1 24.8308
R27 plus.n8 plus.n7 24.8308
R28 plus.n18 plus.n17 24.8308
R29 plus.n12 plus.n11 24.8308
R30 plus plus.n19 24.1998
R31 plus plus.n9 7.99292
R32 plus.n3 plus.n0 0.189894
R33 plus.n9 plus.n0 0.189894
R34 plus.n19 plus.n10 0.189894
R35 plus.n13 plus.n10 0.189894
R36 drain_left.n5 drain_left.t7 260.433
R37 drain_left.n1 drain_left.t8 260.432
R38 drain_left.n3 drain_left.n2 240.452
R39 drain_left.n7 drain_left.n6 240.132
R40 drain_left.n5 drain_left.n4 240.132
R41 drain_left.n1 drain_left.n0 240.131
R42 drain_left drain_left.n3 21.1587
R43 drain_left.n2 drain_left.t0 19.8005
R44 drain_left.n2 drain_left.t3 19.8005
R45 drain_left.n0 drain_left.t6 19.8005
R46 drain_left.n0 drain_left.t4 19.8005
R47 drain_left.n6 drain_left.t5 19.8005
R48 drain_left.n6 drain_left.t2 19.8005
R49 drain_left.n4 drain_left.t1 19.8005
R50 drain_left.n4 drain_left.t9 19.8005
R51 drain_left drain_left.n7 6.15322
R52 drain_left.n7 drain_left.n5 0.5005
R53 drain_left.n3 drain_left.n1 0.070154
R54 source.n0 source.t15 243.255
R55 source.n5 source.t3 243.255
R56 source.n19 source.t9 243.254
R57 source.n14 source.t12 243.254
R58 source.n2 source.n1 223.454
R59 source.n4 source.n3 223.454
R60 source.n7 source.n6 223.454
R61 source.n9 source.n8 223.454
R62 source.n18 source.n17 223.453
R63 source.n16 source.n15 223.453
R64 source.n13 source.n12 223.453
R65 source.n11 source.n10 223.453
R66 source.n17 source.t5 19.8005
R67 source.n17 source.t2 19.8005
R68 source.n15 source.t8 19.8005
R69 source.n15 source.t0 19.8005
R70 source.n12 source.t11 19.8005
R71 source.n12 source.t16 19.8005
R72 source.n10 source.t13 19.8005
R73 source.n10 source.t10 19.8005
R74 source.n1 source.t14 19.8005
R75 source.n1 source.t19 19.8005
R76 source.n3 source.t17 19.8005
R77 source.n3 source.t18 19.8005
R78 source.n6 source.t7 19.8005
R79 source.n6 source.t1 19.8005
R80 source.n8 source.t6 19.8005
R81 source.n8 source.t4 19.8005
R82 source.n11 source.n9 13.9544
R83 source.n20 source.n0 7.94146
R84 source.n20 source.n19 5.51343
R85 source.n5 source.n4 0.720328
R86 source.n16 source.n14 0.720328
R87 source.n9 source.n7 0.5005
R88 source.n7 source.n5 0.5005
R89 source.n4 source.n2 0.5005
R90 source.n2 source.n0 0.5005
R91 source.n13 source.n11 0.5005
R92 source.n14 source.n13 0.5005
R93 source.n18 source.n16 0.5005
R94 source.n19 source.n18 0.5005
R95 source source.n20 0.188
R96 minus.n8 minus.t7 281.606
R97 minus.n2 minus.t6 281.606
R98 minus.n18 minus.t3 281.606
R99 minus.n12 minus.t4 281.606
R100 minus.n7 minus.t1 221.72
R101 minus.n5 minus.t5 221.72
R102 minus.n1 minus.t2 221.72
R103 minus.n17 minus.t9 221.72
R104 minus.n15 minus.t0 221.72
R105 minus.n11 minus.t8 221.72
R106 minus.n3 minus.n2 161.489
R107 minus.n13 minus.n12 161.489
R108 minus.n9 minus.n8 161.3
R109 minus.n6 minus.n0 161.3
R110 minus.n4 minus.n3 161.3
R111 minus.n19 minus.n18 161.3
R112 minus.n16 minus.n10 161.3
R113 minus.n14 minus.n13 161.3
R114 minus.n7 minus.n6 48.2005
R115 minus.n4 minus.n1 48.2005
R116 minus.n14 minus.n11 48.2005
R117 minus.n17 minus.n16 48.2005
R118 minus.n6 minus.n5 36.5157
R119 minus.n5 minus.n4 36.5157
R120 minus.n15 minus.n14 36.5157
R121 minus.n16 minus.n15 36.5157
R122 minus.n20 minus.n9 26.152
R123 minus.n8 minus.n7 24.8308
R124 minus.n2 minus.n1 24.8308
R125 minus.n12 minus.n11 24.8308
R126 minus.n18 minus.n17 24.8308
R127 minus.n20 minus.n19 6.51565
R128 minus.n9 minus.n0 0.189894
R129 minus.n3 minus.n0 0.189894
R130 minus.n13 minus.n10 0.189894
R131 minus.n19 minus.n10 0.189894
R132 minus minus.n20 0.188
R133 drain_right.n1 drain_right.t5 260.432
R134 drain_right.n7 drain_right.t2 259.933
R135 drain_right.n6 drain_right.n4 240.632
R136 drain_right.n3 drain_right.n2 240.452
R137 drain_right.n6 drain_right.n5 240.132
R138 drain_right.n1 drain_right.n0 240.131
R139 drain_right drain_right.n3 20.6055
R140 drain_right.n2 drain_right.t0 19.8005
R141 drain_right.n2 drain_right.t6 19.8005
R142 drain_right.n0 drain_right.t1 19.8005
R143 drain_right.n0 drain_right.t9 19.8005
R144 drain_right.n4 drain_right.t7 19.8005
R145 drain_right.n4 drain_right.t3 19.8005
R146 drain_right.n5 drain_right.t8 19.8005
R147 drain_right.n5 drain_right.t4 19.8005
R148 drain_right drain_right.n7 5.90322
R149 drain_right.n7 drain_right.n6 0.5005
R150 drain_right.n3 drain_right.n1 0.070154
C0 plus source 0.838336f
C1 drain_left minus 0.178716f
C2 drain_right minus 0.650248f
C3 drain_left source 3.82711f
C4 drain_right source 3.82461f
C5 drain_left plus 0.784132f
C6 drain_right plus 0.296839f
C7 drain_left drain_right 0.689458f
C8 minus source 0.824415f
C9 plus minus 2.88231f
C10 drain_right a_n1412_n1088# 3.14982f
C11 drain_left a_n1412_n1088# 3.34789f
C12 source a_n1412_n1088# 2.005897f
C13 minus a_n1412_n1088# 4.544176f
C14 plus a_n1412_n1088# 5.264663f
C15 drain_right.t5 a_n1412_n1088# 0.11669f
C16 drain_right.t1 a_n1412_n1088# 0.018796f
C17 drain_right.t9 a_n1412_n1088# 0.018796f
C18 drain_right.n0 a_n1412_n1088# 0.073037f
C19 drain_right.n1 a_n1412_n1088# 0.439763f
C20 drain_right.t0 a_n1412_n1088# 0.018796f
C21 drain_right.t6 a_n1412_n1088# 0.018796f
C22 drain_right.n2 a_n1412_n1088# 0.073357f
C23 drain_right.n3 a_n1412_n1088# 0.727219f
C24 drain_right.t7 a_n1412_n1088# 0.018796f
C25 drain_right.t3 a_n1412_n1088# 0.018796f
C26 drain_right.n4 a_n1412_n1088# 0.073562f
C27 drain_right.t8 a_n1412_n1088# 0.018796f
C28 drain_right.t4 a_n1412_n1088# 0.018796f
C29 drain_right.n5 a_n1412_n1088# 0.073037f
C30 drain_right.n6 a_n1412_n1088# 0.495016f
C31 drain_right.t2 a_n1412_n1088# 0.116263f
C32 drain_right.n7 a_n1412_n1088# 0.418158f
C33 minus.n0 a_n1412_n1088# 0.036647f
C34 minus.t7 a_n1412_n1088# 0.0356f
C35 minus.t1 a_n1412_n1088# 0.028243f
C36 minus.t5 a_n1412_n1088# 0.028243f
C37 minus.t2 a_n1412_n1088# 0.028243f
C38 minus.n1 a_n1412_n1088# 0.030982f
C39 minus.t6 a_n1412_n1088# 0.0356f
C40 minus.n2 a_n1412_n1088# 0.041263f
C41 minus.n3 a_n1412_n1088# 0.086115f
C42 minus.n4 a_n1412_n1088# 0.013965f
C43 minus.n5 a_n1412_n1088# 0.030982f
C44 minus.n6 a_n1412_n1088# 0.013965f
C45 minus.n7 a_n1412_n1088# 0.030982f
C46 minus.n8 a_n1412_n1088# 0.041204f
C47 minus.n9 a_n1412_n1088# 0.748205f
C48 minus.n10 a_n1412_n1088# 0.036647f
C49 minus.t9 a_n1412_n1088# 0.028243f
C50 minus.t0 a_n1412_n1088# 0.028243f
C51 minus.t8 a_n1412_n1088# 0.028243f
C52 minus.n11 a_n1412_n1088# 0.030982f
C53 minus.t4 a_n1412_n1088# 0.0356f
C54 minus.n12 a_n1412_n1088# 0.041263f
C55 minus.n13 a_n1412_n1088# 0.086115f
C56 minus.n14 a_n1412_n1088# 0.013965f
C57 minus.n15 a_n1412_n1088# 0.030982f
C58 minus.n16 a_n1412_n1088# 0.013965f
C59 minus.n17 a_n1412_n1088# 0.030982f
C60 minus.t3 a_n1412_n1088# 0.0356f
C61 minus.n18 a_n1412_n1088# 0.041204f
C62 minus.n19 a_n1412_n1088# 0.24094f
C63 minus.n20 a_n1412_n1088# 0.922722f
C64 source.t15 a_n1412_n1088# 0.138941f
C65 source.n0 a_n1412_n1088# 0.588727f
C66 source.t14 a_n1412_n1088# 0.024963f
C67 source.t19 a_n1412_n1088# 0.024963f
C68 source.n1 a_n1412_n1088# 0.08096f
C69 source.n2 a_n1412_n1088# 0.295803f
C70 source.t17 a_n1412_n1088# 0.024963f
C71 source.t18 a_n1412_n1088# 0.024963f
C72 source.n3 a_n1412_n1088# 0.08096f
C73 source.n4 a_n1412_n1088# 0.318179f
C74 source.t3 a_n1412_n1088# 0.138941f
C75 source.n5 a_n1412_n1088# 0.328278f
C76 source.t7 a_n1412_n1088# 0.024963f
C77 source.t1 a_n1412_n1088# 0.024963f
C78 source.n6 a_n1412_n1088# 0.08096f
C79 source.n7 a_n1412_n1088# 0.295803f
C80 source.t6 a_n1412_n1088# 0.024963f
C81 source.t4 a_n1412_n1088# 0.024963f
C82 source.n8 a_n1412_n1088# 0.08096f
C83 source.n9 a_n1412_n1088# 0.881741f
C84 source.t13 a_n1412_n1088# 0.024963f
C85 source.t10 a_n1412_n1088# 0.024963f
C86 source.n10 a_n1412_n1088# 0.080959f
C87 source.n11 a_n1412_n1088# 0.881742f
C88 source.t11 a_n1412_n1088# 0.024963f
C89 source.t16 a_n1412_n1088# 0.024963f
C90 source.n12 a_n1412_n1088# 0.080959f
C91 source.n13 a_n1412_n1088# 0.295803f
C92 source.t12 a_n1412_n1088# 0.138941f
C93 source.n14 a_n1412_n1088# 0.328279f
C94 source.t8 a_n1412_n1088# 0.024963f
C95 source.t0 a_n1412_n1088# 0.024963f
C96 source.n15 a_n1412_n1088# 0.080959f
C97 source.n16 a_n1412_n1088# 0.318179f
C98 source.t5 a_n1412_n1088# 0.024963f
C99 source.t2 a_n1412_n1088# 0.024963f
C100 source.n17 a_n1412_n1088# 0.080959f
C101 source.n18 a_n1412_n1088# 0.295803f
C102 source.t9 a_n1412_n1088# 0.138941f
C103 source.n19 a_n1412_n1088# 0.477643f
C104 source.n20 a_n1412_n1088# 0.637992f
C105 drain_left.t8 a_n1412_n1088# 0.113901f
C106 drain_left.t6 a_n1412_n1088# 0.018347f
C107 drain_left.t4 a_n1412_n1088# 0.018347f
C108 drain_left.n0 a_n1412_n1088# 0.071291f
C109 drain_left.n1 a_n1412_n1088# 0.429252f
C110 drain_left.t0 a_n1412_n1088# 0.018347f
C111 drain_left.t3 a_n1412_n1088# 0.018347f
C112 drain_left.n2 a_n1412_n1088# 0.071603f
C113 drain_left.n3 a_n1412_n1088# 0.754839f
C114 drain_left.t7 a_n1412_n1088# 0.113901f
C115 drain_left.t1 a_n1412_n1088# 0.018347f
C116 drain_left.t9 a_n1412_n1088# 0.018347f
C117 drain_left.n4 a_n1412_n1088# 0.071291f
C118 drain_left.n5 a_n1412_n1088# 0.453719f
C119 drain_left.t5 a_n1412_n1088# 0.018347f
C120 drain_left.t2 a_n1412_n1088# 0.018347f
C121 drain_left.n6 a_n1412_n1088# 0.071291f
C122 drain_left.n7 a_n1412_n1088# 0.428816f
C123 plus.n0 a_n1412_n1088# 0.037608f
C124 plus.t0 a_n1412_n1088# 0.028984f
C125 plus.t5 a_n1412_n1088# 0.028984f
C126 plus.t1 a_n1412_n1088# 0.028984f
C127 plus.n1 a_n1412_n1088# 0.031794f
C128 plus.t2 a_n1412_n1088# 0.036534f
C129 plus.n2 a_n1412_n1088# 0.042345f
C130 plus.n3 a_n1412_n1088# 0.088373f
C131 plus.n4 a_n1412_n1088# 0.014331f
C132 plus.n5 a_n1412_n1088# 0.031794f
C133 plus.n6 a_n1412_n1088# 0.014331f
C134 plus.n7 a_n1412_n1088# 0.031794f
C135 plus.t4 a_n1412_n1088# 0.036534f
C136 plus.n8 a_n1412_n1088# 0.042285f
C137 plus.n9 a_n1412_n1088# 0.259302f
C138 plus.n10 a_n1412_n1088# 0.037608f
C139 plus.t6 a_n1412_n1088# 0.036534f
C140 plus.t9 a_n1412_n1088# 0.028984f
C141 plus.t8 a_n1412_n1088# 0.028984f
C142 plus.t3 a_n1412_n1088# 0.028984f
C143 plus.n11 a_n1412_n1088# 0.031794f
C144 plus.t7 a_n1412_n1088# 0.036534f
C145 plus.n12 a_n1412_n1088# 0.042345f
C146 plus.n13 a_n1412_n1088# 0.088373f
C147 plus.n14 a_n1412_n1088# 0.014331f
C148 plus.n15 a_n1412_n1088# 0.031794f
C149 plus.n16 a_n1412_n1088# 0.014331f
C150 plus.n17 a_n1412_n1088# 0.031794f
C151 plus.n18 a_n1412_n1088# 0.042285f
C152 plus.n19 a_n1412_n1088# 0.749244f
.ends

