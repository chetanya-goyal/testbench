* NGSPICE file created from diffpair466.ext - technology: sky130A

.subckt diffpair466 minus drain_right drain_left source plus
X0 a_n2364_n3288# a_n2364_n3288# a_n2364_n3288# a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.7
X1 source.t27 plus.t0 drain_left.t2 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X2 drain_left.t1 plus.t1 source.t26 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X3 drain_left.t0 plus.t2 source.t25 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X4 drain_right.t13 minus.t0 source.t0 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X5 drain_left.t9 plus.t3 source.t24 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X6 source.t11 minus.t1 drain_right.t12 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X7 source.t2 minus.t2 drain_right.t11 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X8 a_n2364_n3288# a_n2364_n3288# a_n2364_n3288# a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X9 drain_left.t6 plus.t4 source.t23 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X10 drain_left.t5 plus.t5 source.t22 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X11 drain_right.t10 minus.t3 source.t6 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X12 source.t21 plus.t6 drain_left.t12 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X13 drain_right.t9 minus.t4 source.t8 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X14 drain_left.t11 plus.t7 source.t20 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X15 a_n2364_n3288# a_n2364_n3288# a_n2364_n3288# a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X16 drain_right.t8 minus.t5 source.t4 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X17 source.t19 plus.t8 drain_left.t10 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X18 source.t18 plus.t9 drain_left.t13 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X19 drain_right.t7 minus.t6 source.t13 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X20 a_n2364_n3288# a_n2364_n3288# a_n2364_n3288# a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X21 source.t17 plus.t10 drain_left.t7 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X22 drain_left.t8 plus.t11 source.t16 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X23 source.t12 minus.t7 drain_right.t6 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X24 drain_right.t5 minus.t8 source.t5 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X25 drain_left.t3 plus.t12 source.t15 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X26 drain_right.t4 minus.t9 source.t7 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X27 source.t14 plus.t13 drain_left.t4 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X28 source.t9 minus.t10 drain_right.t3 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X29 source.t1 minus.t11 drain_right.t2 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X30 source.t3 minus.t12 drain_right.t1 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X31 drain_right.t0 minus.t13 source.t10 a_n2364_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
R0 plus.n5 plus.t5 493.108
R1 plus.n27 plus.t12 493.108
R2 plus.n20 plus.t2 469.262
R3 plus.n18 plus.t9 469.262
R4 plus.n2 plus.t4 469.262
R5 plus.n12 plus.t8 469.262
R6 plus.n4 plus.t3 469.262
R7 plus.n6 plus.t10 469.262
R8 plus.n42 plus.t1 469.262
R9 plus.n40 plus.t0 469.262
R10 plus.n24 plus.t7 469.262
R11 plus.n34 plus.t6 469.262
R12 plus.n26 plus.t11 469.262
R13 plus.n28 plus.t13 469.262
R14 plus.n8 plus.n7 161.3
R15 plus.n9 plus.n4 161.3
R16 plus.n11 plus.n10 161.3
R17 plus.n12 plus.n3 161.3
R18 plus.n14 plus.n13 161.3
R19 plus.n15 plus.n2 161.3
R20 plus.n17 plus.n16 161.3
R21 plus.n18 plus.n1 161.3
R22 plus.n19 plus.n0 161.3
R23 plus.n21 plus.n20 161.3
R24 plus.n30 plus.n29 161.3
R25 plus.n31 plus.n26 161.3
R26 plus.n33 plus.n32 161.3
R27 plus.n34 plus.n25 161.3
R28 plus.n36 plus.n35 161.3
R29 plus.n37 plus.n24 161.3
R30 plus.n39 plus.n38 161.3
R31 plus.n40 plus.n23 161.3
R32 plus.n41 plus.n22 161.3
R33 plus.n43 plus.n42 161.3
R34 plus.n30 plus.n27 44.9119
R35 plus.n8 plus.n5 44.9119
R36 plus.n20 plus.n19 35.055
R37 plus.n42 plus.n41 35.055
R38 plus plus.n43 32.107
R39 plus.n18 plus.n17 30.6732
R40 plus.n7 plus.n6 30.6732
R41 plus.n40 plus.n39 30.6732
R42 plus.n29 plus.n28 30.6732
R43 plus.n13 plus.n2 26.2914
R44 plus.n11 plus.n4 26.2914
R45 plus.n35 plus.n24 26.2914
R46 plus.n33 plus.n26 26.2914
R47 plus.n13 plus.n12 21.9096
R48 plus.n12 plus.n11 21.9096
R49 plus.n35 plus.n34 21.9096
R50 plus.n34 plus.n33 21.9096
R51 plus.n28 plus.n27 17.739
R52 plus.n6 plus.n5 17.739
R53 plus.n17 plus.n2 17.5278
R54 plus.n7 plus.n4 17.5278
R55 plus.n39 plus.n24 17.5278
R56 plus.n29 plus.n26 17.5278
R57 plus.n19 plus.n18 13.146
R58 plus.n41 plus.n40 13.146
R59 plus plus.n21 12.2941
R60 plus.n9 plus.n8 0.189894
R61 plus.n10 plus.n9 0.189894
R62 plus.n10 plus.n3 0.189894
R63 plus.n14 plus.n3 0.189894
R64 plus.n15 plus.n14 0.189894
R65 plus.n16 plus.n15 0.189894
R66 plus.n16 plus.n1 0.189894
R67 plus.n1 plus.n0 0.189894
R68 plus.n21 plus.n0 0.189894
R69 plus.n43 plus.n22 0.189894
R70 plus.n23 plus.n22 0.189894
R71 plus.n38 plus.n23 0.189894
R72 plus.n38 plus.n37 0.189894
R73 plus.n37 plus.n36 0.189894
R74 plus.n36 plus.n25 0.189894
R75 plus.n32 plus.n25 0.189894
R76 plus.n32 plus.n31 0.189894
R77 plus.n31 plus.n30 0.189894
R78 drain_left.n60 drain_left.n0 289.615
R79 drain_left.n131 drain_left.n71 289.615
R80 drain_left.n20 drain_left.n19 185
R81 drain_left.n25 drain_left.n24 185
R82 drain_left.n27 drain_left.n26 185
R83 drain_left.n16 drain_left.n15 185
R84 drain_left.n33 drain_left.n32 185
R85 drain_left.n35 drain_left.n34 185
R86 drain_left.n12 drain_left.n11 185
R87 drain_left.n42 drain_left.n41 185
R88 drain_left.n43 drain_left.n10 185
R89 drain_left.n45 drain_left.n44 185
R90 drain_left.n8 drain_left.n7 185
R91 drain_left.n51 drain_left.n50 185
R92 drain_left.n53 drain_left.n52 185
R93 drain_left.n4 drain_left.n3 185
R94 drain_left.n59 drain_left.n58 185
R95 drain_left.n61 drain_left.n60 185
R96 drain_left.n132 drain_left.n131 185
R97 drain_left.n130 drain_left.n129 185
R98 drain_left.n75 drain_left.n74 185
R99 drain_left.n124 drain_left.n123 185
R100 drain_left.n122 drain_left.n121 185
R101 drain_left.n79 drain_left.n78 185
R102 drain_left.n116 drain_left.n115 185
R103 drain_left.n114 drain_left.n81 185
R104 drain_left.n113 drain_left.n112 185
R105 drain_left.n84 drain_left.n82 185
R106 drain_left.n107 drain_left.n106 185
R107 drain_left.n105 drain_left.n104 185
R108 drain_left.n88 drain_left.n87 185
R109 drain_left.n99 drain_left.n98 185
R110 drain_left.n97 drain_left.n96 185
R111 drain_left.n92 drain_left.n91 185
R112 drain_left.n21 drain_left.t1 149.524
R113 drain_left.n93 drain_left.t5 149.524
R114 drain_left.n25 drain_left.n19 104.615
R115 drain_left.n26 drain_left.n25 104.615
R116 drain_left.n26 drain_left.n15 104.615
R117 drain_left.n33 drain_left.n15 104.615
R118 drain_left.n34 drain_left.n33 104.615
R119 drain_left.n34 drain_left.n11 104.615
R120 drain_left.n42 drain_left.n11 104.615
R121 drain_left.n43 drain_left.n42 104.615
R122 drain_left.n44 drain_left.n43 104.615
R123 drain_left.n44 drain_left.n7 104.615
R124 drain_left.n51 drain_left.n7 104.615
R125 drain_left.n52 drain_left.n51 104.615
R126 drain_left.n52 drain_left.n3 104.615
R127 drain_left.n59 drain_left.n3 104.615
R128 drain_left.n60 drain_left.n59 104.615
R129 drain_left.n131 drain_left.n130 104.615
R130 drain_left.n130 drain_left.n74 104.615
R131 drain_left.n123 drain_left.n74 104.615
R132 drain_left.n123 drain_left.n122 104.615
R133 drain_left.n122 drain_left.n78 104.615
R134 drain_left.n115 drain_left.n78 104.615
R135 drain_left.n115 drain_left.n114 104.615
R136 drain_left.n114 drain_left.n113 104.615
R137 drain_left.n113 drain_left.n82 104.615
R138 drain_left.n106 drain_left.n82 104.615
R139 drain_left.n106 drain_left.n105 104.615
R140 drain_left.n105 drain_left.n87 104.615
R141 drain_left.n98 drain_left.n87 104.615
R142 drain_left.n98 drain_left.n97 104.615
R143 drain_left.n97 drain_left.n91 104.615
R144 drain_left.n69 drain_left.n67 60.4404
R145 drain_left.n139 drain_left.n138 59.5527
R146 drain_left.n137 drain_left.n136 59.5527
R147 drain_left.n69 drain_left.n68 59.5525
R148 drain_left.n66 drain_left.n65 59.5525
R149 drain_left.n141 drain_left.n140 59.5525
R150 drain_left.t1 drain_left.n19 52.3082
R151 drain_left.t5 drain_left.n91 52.3082
R152 drain_left.n66 drain_left.n64 47.4248
R153 drain_left.n137 drain_left.n135 47.4248
R154 drain_left drain_left.n70 32.4727
R155 drain_left.n45 drain_left.n10 13.1884
R156 drain_left.n116 drain_left.n81 13.1884
R157 drain_left.n41 drain_left.n40 12.8005
R158 drain_left.n46 drain_left.n8 12.8005
R159 drain_left.n117 drain_left.n79 12.8005
R160 drain_left.n112 drain_left.n83 12.8005
R161 drain_left.n39 drain_left.n12 12.0247
R162 drain_left.n50 drain_left.n49 12.0247
R163 drain_left.n121 drain_left.n120 12.0247
R164 drain_left.n111 drain_left.n84 12.0247
R165 drain_left.n36 drain_left.n35 11.249
R166 drain_left.n53 drain_left.n6 11.249
R167 drain_left.n124 drain_left.n77 11.249
R168 drain_left.n108 drain_left.n107 11.249
R169 drain_left.n32 drain_left.n14 10.4732
R170 drain_left.n54 drain_left.n4 10.4732
R171 drain_left.n125 drain_left.n75 10.4732
R172 drain_left.n104 drain_left.n86 10.4732
R173 drain_left.n21 drain_left.n20 10.2747
R174 drain_left.n93 drain_left.n92 10.2747
R175 drain_left.n31 drain_left.n16 9.69747
R176 drain_left.n58 drain_left.n57 9.69747
R177 drain_left.n129 drain_left.n128 9.69747
R178 drain_left.n103 drain_left.n88 9.69747
R179 drain_left.n64 drain_left.n63 9.45567
R180 drain_left.n135 drain_left.n134 9.45567
R181 drain_left.n63 drain_left.n62 9.3005
R182 drain_left.n2 drain_left.n1 9.3005
R183 drain_left.n57 drain_left.n56 9.3005
R184 drain_left.n55 drain_left.n54 9.3005
R185 drain_left.n6 drain_left.n5 9.3005
R186 drain_left.n49 drain_left.n48 9.3005
R187 drain_left.n47 drain_left.n46 9.3005
R188 drain_left.n23 drain_left.n22 9.3005
R189 drain_left.n18 drain_left.n17 9.3005
R190 drain_left.n29 drain_left.n28 9.3005
R191 drain_left.n31 drain_left.n30 9.3005
R192 drain_left.n14 drain_left.n13 9.3005
R193 drain_left.n37 drain_left.n36 9.3005
R194 drain_left.n39 drain_left.n38 9.3005
R195 drain_left.n40 drain_left.n9 9.3005
R196 drain_left.n95 drain_left.n94 9.3005
R197 drain_left.n90 drain_left.n89 9.3005
R198 drain_left.n101 drain_left.n100 9.3005
R199 drain_left.n103 drain_left.n102 9.3005
R200 drain_left.n86 drain_left.n85 9.3005
R201 drain_left.n109 drain_left.n108 9.3005
R202 drain_left.n111 drain_left.n110 9.3005
R203 drain_left.n83 drain_left.n80 9.3005
R204 drain_left.n134 drain_left.n133 9.3005
R205 drain_left.n73 drain_left.n72 9.3005
R206 drain_left.n128 drain_left.n127 9.3005
R207 drain_left.n126 drain_left.n125 9.3005
R208 drain_left.n77 drain_left.n76 9.3005
R209 drain_left.n120 drain_left.n119 9.3005
R210 drain_left.n118 drain_left.n117 9.3005
R211 drain_left.n28 drain_left.n27 8.92171
R212 drain_left.n61 drain_left.n2 8.92171
R213 drain_left.n132 drain_left.n73 8.92171
R214 drain_left.n100 drain_left.n99 8.92171
R215 drain_left.n24 drain_left.n18 8.14595
R216 drain_left.n62 drain_left.n0 8.14595
R217 drain_left.n133 drain_left.n71 8.14595
R218 drain_left.n96 drain_left.n90 8.14595
R219 drain_left.n23 drain_left.n20 7.3702
R220 drain_left.n95 drain_left.n92 7.3702
R221 drain_left drain_left.n141 6.54115
R222 drain_left.n24 drain_left.n23 5.81868
R223 drain_left.n64 drain_left.n0 5.81868
R224 drain_left.n135 drain_left.n71 5.81868
R225 drain_left.n96 drain_left.n95 5.81868
R226 drain_left.n27 drain_left.n18 5.04292
R227 drain_left.n62 drain_left.n61 5.04292
R228 drain_left.n133 drain_left.n132 5.04292
R229 drain_left.n99 drain_left.n90 5.04292
R230 drain_left.n28 drain_left.n16 4.26717
R231 drain_left.n58 drain_left.n2 4.26717
R232 drain_left.n129 drain_left.n73 4.26717
R233 drain_left.n100 drain_left.n88 4.26717
R234 drain_left.n32 drain_left.n31 3.49141
R235 drain_left.n57 drain_left.n4 3.49141
R236 drain_left.n128 drain_left.n75 3.49141
R237 drain_left.n104 drain_left.n103 3.49141
R238 drain_left.n22 drain_left.n21 2.84303
R239 drain_left.n94 drain_left.n93 2.84303
R240 drain_left.n35 drain_left.n14 2.71565
R241 drain_left.n54 drain_left.n53 2.71565
R242 drain_left.n125 drain_left.n124 2.71565
R243 drain_left.n107 drain_left.n86 2.71565
R244 drain_left.n36 drain_left.n12 1.93989
R245 drain_left.n50 drain_left.n6 1.93989
R246 drain_left.n121 drain_left.n77 1.93989
R247 drain_left.n108 drain_left.n84 1.93989
R248 drain_left.n67 drain_left.t4 1.6505
R249 drain_left.n67 drain_left.t3 1.6505
R250 drain_left.n68 drain_left.t12 1.6505
R251 drain_left.n68 drain_left.t8 1.6505
R252 drain_left.n65 drain_left.t2 1.6505
R253 drain_left.n65 drain_left.t11 1.6505
R254 drain_left.n140 drain_left.t13 1.6505
R255 drain_left.n140 drain_left.t0 1.6505
R256 drain_left.n138 drain_left.t10 1.6505
R257 drain_left.n138 drain_left.t6 1.6505
R258 drain_left.n136 drain_left.t7 1.6505
R259 drain_left.n136 drain_left.t9 1.6505
R260 drain_left.n41 drain_left.n39 1.16414
R261 drain_left.n49 drain_left.n8 1.16414
R262 drain_left.n120 drain_left.n79 1.16414
R263 drain_left.n112 drain_left.n111 1.16414
R264 drain_left.n139 drain_left.n137 0.888431
R265 drain_left.n141 drain_left.n139 0.888431
R266 drain_left.n70 drain_left.n66 0.611102
R267 drain_left.n40 drain_left.n10 0.388379
R268 drain_left.n46 drain_left.n45 0.388379
R269 drain_left.n117 drain_left.n116 0.388379
R270 drain_left.n83 drain_left.n81 0.388379
R271 drain_left.n70 drain_left.n69 0.167137
R272 drain_left.n22 drain_left.n17 0.155672
R273 drain_left.n29 drain_left.n17 0.155672
R274 drain_left.n30 drain_left.n29 0.155672
R275 drain_left.n30 drain_left.n13 0.155672
R276 drain_left.n37 drain_left.n13 0.155672
R277 drain_left.n38 drain_left.n37 0.155672
R278 drain_left.n38 drain_left.n9 0.155672
R279 drain_left.n47 drain_left.n9 0.155672
R280 drain_left.n48 drain_left.n47 0.155672
R281 drain_left.n48 drain_left.n5 0.155672
R282 drain_left.n55 drain_left.n5 0.155672
R283 drain_left.n56 drain_left.n55 0.155672
R284 drain_left.n56 drain_left.n1 0.155672
R285 drain_left.n63 drain_left.n1 0.155672
R286 drain_left.n134 drain_left.n72 0.155672
R287 drain_left.n127 drain_left.n72 0.155672
R288 drain_left.n127 drain_left.n126 0.155672
R289 drain_left.n126 drain_left.n76 0.155672
R290 drain_left.n119 drain_left.n76 0.155672
R291 drain_left.n119 drain_left.n118 0.155672
R292 drain_left.n118 drain_left.n80 0.155672
R293 drain_left.n110 drain_left.n80 0.155672
R294 drain_left.n110 drain_left.n109 0.155672
R295 drain_left.n109 drain_left.n85 0.155672
R296 drain_left.n102 drain_left.n85 0.155672
R297 drain_left.n102 drain_left.n101 0.155672
R298 drain_left.n101 drain_left.n89 0.155672
R299 drain_left.n94 drain_left.n89 0.155672
R300 source.n282 source.n222 289.615
R301 source.n210 source.n150 289.615
R302 source.n60 source.n0 289.615
R303 source.n132 source.n72 289.615
R304 source.n242 source.n241 185
R305 source.n247 source.n246 185
R306 source.n249 source.n248 185
R307 source.n238 source.n237 185
R308 source.n255 source.n254 185
R309 source.n257 source.n256 185
R310 source.n234 source.n233 185
R311 source.n264 source.n263 185
R312 source.n265 source.n232 185
R313 source.n267 source.n266 185
R314 source.n230 source.n229 185
R315 source.n273 source.n272 185
R316 source.n275 source.n274 185
R317 source.n226 source.n225 185
R318 source.n281 source.n280 185
R319 source.n283 source.n282 185
R320 source.n170 source.n169 185
R321 source.n175 source.n174 185
R322 source.n177 source.n176 185
R323 source.n166 source.n165 185
R324 source.n183 source.n182 185
R325 source.n185 source.n184 185
R326 source.n162 source.n161 185
R327 source.n192 source.n191 185
R328 source.n193 source.n160 185
R329 source.n195 source.n194 185
R330 source.n158 source.n157 185
R331 source.n201 source.n200 185
R332 source.n203 source.n202 185
R333 source.n154 source.n153 185
R334 source.n209 source.n208 185
R335 source.n211 source.n210 185
R336 source.n61 source.n60 185
R337 source.n59 source.n58 185
R338 source.n4 source.n3 185
R339 source.n53 source.n52 185
R340 source.n51 source.n50 185
R341 source.n8 source.n7 185
R342 source.n45 source.n44 185
R343 source.n43 source.n10 185
R344 source.n42 source.n41 185
R345 source.n13 source.n11 185
R346 source.n36 source.n35 185
R347 source.n34 source.n33 185
R348 source.n17 source.n16 185
R349 source.n28 source.n27 185
R350 source.n26 source.n25 185
R351 source.n21 source.n20 185
R352 source.n133 source.n132 185
R353 source.n131 source.n130 185
R354 source.n76 source.n75 185
R355 source.n125 source.n124 185
R356 source.n123 source.n122 185
R357 source.n80 source.n79 185
R358 source.n117 source.n116 185
R359 source.n115 source.n82 185
R360 source.n114 source.n113 185
R361 source.n85 source.n83 185
R362 source.n108 source.n107 185
R363 source.n106 source.n105 185
R364 source.n89 source.n88 185
R365 source.n100 source.n99 185
R366 source.n98 source.n97 185
R367 source.n93 source.n92 185
R368 source.n243 source.t5 149.524
R369 source.n171 source.t15 149.524
R370 source.n22 source.t25 149.524
R371 source.n94 source.t13 149.524
R372 source.n247 source.n241 104.615
R373 source.n248 source.n247 104.615
R374 source.n248 source.n237 104.615
R375 source.n255 source.n237 104.615
R376 source.n256 source.n255 104.615
R377 source.n256 source.n233 104.615
R378 source.n264 source.n233 104.615
R379 source.n265 source.n264 104.615
R380 source.n266 source.n265 104.615
R381 source.n266 source.n229 104.615
R382 source.n273 source.n229 104.615
R383 source.n274 source.n273 104.615
R384 source.n274 source.n225 104.615
R385 source.n281 source.n225 104.615
R386 source.n282 source.n281 104.615
R387 source.n175 source.n169 104.615
R388 source.n176 source.n175 104.615
R389 source.n176 source.n165 104.615
R390 source.n183 source.n165 104.615
R391 source.n184 source.n183 104.615
R392 source.n184 source.n161 104.615
R393 source.n192 source.n161 104.615
R394 source.n193 source.n192 104.615
R395 source.n194 source.n193 104.615
R396 source.n194 source.n157 104.615
R397 source.n201 source.n157 104.615
R398 source.n202 source.n201 104.615
R399 source.n202 source.n153 104.615
R400 source.n209 source.n153 104.615
R401 source.n210 source.n209 104.615
R402 source.n60 source.n59 104.615
R403 source.n59 source.n3 104.615
R404 source.n52 source.n3 104.615
R405 source.n52 source.n51 104.615
R406 source.n51 source.n7 104.615
R407 source.n44 source.n7 104.615
R408 source.n44 source.n43 104.615
R409 source.n43 source.n42 104.615
R410 source.n42 source.n11 104.615
R411 source.n35 source.n11 104.615
R412 source.n35 source.n34 104.615
R413 source.n34 source.n16 104.615
R414 source.n27 source.n16 104.615
R415 source.n27 source.n26 104.615
R416 source.n26 source.n20 104.615
R417 source.n132 source.n131 104.615
R418 source.n131 source.n75 104.615
R419 source.n124 source.n75 104.615
R420 source.n124 source.n123 104.615
R421 source.n123 source.n79 104.615
R422 source.n116 source.n79 104.615
R423 source.n116 source.n115 104.615
R424 source.n115 source.n114 104.615
R425 source.n114 source.n83 104.615
R426 source.n107 source.n83 104.615
R427 source.n107 source.n106 104.615
R428 source.n106 source.n88 104.615
R429 source.n99 source.n88 104.615
R430 source.n99 source.n98 104.615
R431 source.n98 source.n92 104.615
R432 source.t5 source.n241 52.3082
R433 source.t15 source.n169 52.3082
R434 source.t25 source.n20 52.3082
R435 source.t13 source.n92 52.3082
R436 source.n67 source.n66 42.8739
R437 source.n69 source.n68 42.8739
R438 source.n71 source.n70 42.8739
R439 source.n139 source.n138 42.8739
R440 source.n141 source.n140 42.8739
R441 source.n143 source.n142 42.8739
R442 source.n221 source.n220 42.8737
R443 source.n219 source.n218 42.8737
R444 source.n217 source.n216 42.8737
R445 source.n149 source.n148 42.8737
R446 source.n147 source.n146 42.8737
R447 source.n145 source.n144 42.8737
R448 source.n287 source.n286 29.8581
R449 source.n215 source.n214 29.8581
R450 source.n65 source.n64 29.8581
R451 source.n137 source.n136 29.8581
R452 source.n145 source.n143 23.0636
R453 source.n288 source.n65 16.4688
R454 source.n267 source.n232 13.1884
R455 source.n195 source.n160 13.1884
R456 source.n45 source.n10 13.1884
R457 source.n117 source.n82 13.1884
R458 source.n263 source.n262 12.8005
R459 source.n268 source.n230 12.8005
R460 source.n191 source.n190 12.8005
R461 source.n196 source.n158 12.8005
R462 source.n46 source.n8 12.8005
R463 source.n41 source.n12 12.8005
R464 source.n118 source.n80 12.8005
R465 source.n113 source.n84 12.8005
R466 source.n261 source.n234 12.0247
R467 source.n272 source.n271 12.0247
R468 source.n189 source.n162 12.0247
R469 source.n200 source.n199 12.0247
R470 source.n50 source.n49 12.0247
R471 source.n40 source.n13 12.0247
R472 source.n122 source.n121 12.0247
R473 source.n112 source.n85 12.0247
R474 source.n258 source.n257 11.249
R475 source.n275 source.n228 11.249
R476 source.n186 source.n185 11.249
R477 source.n203 source.n156 11.249
R478 source.n53 source.n6 11.249
R479 source.n37 source.n36 11.249
R480 source.n125 source.n78 11.249
R481 source.n109 source.n108 11.249
R482 source.n254 source.n236 10.4732
R483 source.n276 source.n226 10.4732
R484 source.n182 source.n164 10.4732
R485 source.n204 source.n154 10.4732
R486 source.n54 source.n4 10.4732
R487 source.n33 source.n15 10.4732
R488 source.n126 source.n76 10.4732
R489 source.n105 source.n87 10.4732
R490 source.n243 source.n242 10.2747
R491 source.n171 source.n170 10.2747
R492 source.n22 source.n21 10.2747
R493 source.n94 source.n93 10.2747
R494 source.n253 source.n238 9.69747
R495 source.n280 source.n279 9.69747
R496 source.n181 source.n166 9.69747
R497 source.n208 source.n207 9.69747
R498 source.n58 source.n57 9.69747
R499 source.n32 source.n17 9.69747
R500 source.n130 source.n129 9.69747
R501 source.n104 source.n89 9.69747
R502 source.n286 source.n285 9.45567
R503 source.n214 source.n213 9.45567
R504 source.n64 source.n63 9.45567
R505 source.n136 source.n135 9.45567
R506 source.n285 source.n284 9.3005
R507 source.n224 source.n223 9.3005
R508 source.n279 source.n278 9.3005
R509 source.n277 source.n276 9.3005
R510 source.n228 source.n227 9.3005
R511 source.n271 source.n270 9.3005
R512 source.n269 source.n268 9.3005
R513 source.n245 source.n244 9.3005
R514 source.n240 source.n239 9.3005
R515 source.n251 source.n250 9.3005
R516 source.n253 source.n252 9.3005
R517 source.n236 source.n235 9.3005
R518 source.n259 source.n258 9.3005
R519 source.n261 source.n260 9.3005
R520 source.n262 source.n231 9.3005
R521 source.n213 source.n212 9.3005
R522 source.n152 source.n151 9.3005
R523 source.n207 source.n206 9.3005
R524 source.n205 source.n204 9.3005
R525 source.n156 source.n155 9.3005
R526 source.n199 source.n198 9.3005
R527 source.n197 source.n196 9.3005
R528 source.n173 source.n172 9.3005
R529 source.n168 source.n167 9.3005
R530 source.n179 source.n178 9.3005
R531 source.n181 source.n180 9.3005
R532 source.n164 source.n163 9.3005
R533 source.n187 source.n186 9.3005
R534 source.n189 source.n188 9.3005
R535 source.n190 source.n159 9.3005
R536 source.n24 source.n23 9.3005
R537 source.n19 source.n18 9.3005
R538 source.n30 source.n29 9.3005
R539 source.n32 source.n31 9.3005
R540 source.n15 source.n14 9.3005
R541 source.n38 source.n37 9.3005
R542 source.n40 source.n39 9.3005
R543 source.n12 source.n9 9.3005
R544 source.n63 source.n62 9.3005
R545 source.n2 source.n1 9.3005
R546 source.n57 source.n56 9.3005
R547 source.n55 source.n54 9.3005
R548 source.n6 source.n5 9.3005
R549 source.n49 source.n48 9.3005
R550 source.n47 source.n46 9.3005
R551 source.n96 source.n95 9.3005
R552 source.n91 source.n90 9.3005
R553 source.n102 source.n101 9.3005
R554 source.n104 source.n103 9.3005
R555 source.n87 source.n86 9.3005
R556 source.n110 source.n109 9.3005
R557 source.n112 source.n111 9.3005
R558 source.n84 source.n81 9.3005
R559 source.n135 source.n134 9.3005
R560 source.n74 source.n73 9.3005
R561 source.n129 source.n128 9.3005
R562 source.n127 source.n126 9.3005
R563 source.n78 source.n77 9.3005
R564 source.n121 source.n120 9.3005
R565 source.n119 source.n118 9.3005
R566 source.n250 source.n249 8.92171
R567 source.n283 source.n224 8.92171
R568 source.n178 source.n177 8.92171
R569 source.n211 source.n152 8.92171
R570 source.n61 source.n2 8.92171
R571 source.n29 source.n28 8.92171
R572 source.n133 source.n74 8.92171
R573 source.n101 source.n100 8.92171
R574 source.n246 source.n240 8.14595
R575 source.n284 source.n222 8.14595
R576 source.n174 source.n168 8.14595
R577 source.n212 source.n150 8.14595
R578 source.n62 source.n0 8.14595
R579 source.n25 source.n19 8.14595
R580 source.n134 source.n72 8.14595
R581 source.n97 source.n91 8.14595
R582 source.n245 source.n242 7.3702
R583 source.n173 source.n170 7.3702
R584 source.n24 source.n21 7.3702
R585 source.n96 source.n93 7.3702
R586 source.n246 source.n245 5.81868
R587 source.n286 source.n222 5.81868
R588 source.n174 source.n173 5.81868
R589 source.n214 source.n150 5.81868
R590 source.n64 source.n0 5.81868
R591 source.n25 source.n24 5.81868
R592 source.n136 source.n72 5.81868
R593 source.n97 source.n96 5.81868
R594 source.n288 source.n287 5.7074
R595 source.n249 source.n240 5.04292
R596 source.n284 source.n283 5.04292
R597 source.n177 source.n168 5.04292
R598 source.n212 source.n211 5.04292
R599 source.n62 source.n61 5.04292
R600 source.n28 source.n19 5.04292
R601 source.n134 source.n133 5.04292
R602 source.n100 source.n91 5.04292
R603 source.n250 source.n238 4.26717
R604 source.n280 source.n224 4.26717
R605 source.n178 source.n166 4.26717
R606 source.n208 source.n152 4.26717
R607 source.n58 source.n2 4.26717
R608 source.n29 source.n17 4.26717
R609 source.n130 source.n74 4.26717
R610 source.n101 source.n89 4.26717
R611 source.n254 source.n253 3.49141
R612 source.n279 source.n226 3.49141
R613 source.n182 source.n181 3.49141
R614 source.n207 source.n154 3.49141
R615 source.n57 source.n4 3.49141
R616 source.n33 source.n32 3.49141
R617 source.n129 source.n76 3.49141
R618 source.n105 source.n104 3.49141
R619 source.n244 source.n243 2.84303
R620 source.n172 source.n171 2.84303
R621 source.n23 source.n22 2.84303
R622 source.n95 source.n94 2.84303
R623 source.n257 source.n236 2.71565
R624 source.n276 source.n275 2.71565
R625 source.n185 source.n164 2.71565
R626 source.n204 source.n203 2.71565
R627 source.n54 source.n53 2.71565
R628 source.n36 source.n15 2.71565
R629 source.n126 source.n125 2.71565
R630 source.n108 source.n87 2.71565
R631 source.n258 source.n234 1.93989
R632 source.n272 source.n228 1.93989
R633 source.n186 source.n162 1.93989
R634 source.n200 source.n156 1.93989
R635 source.n50 source.n6 1.93989
R636 source.n37 source.n13 1.93989
R637 source.n122 source.n78 1.93989
R638 source.n109 source.n85 1.93989
R639 source.n220 source.t10 1.6505
R640 source.n220 source.t12 1.6505
R641 source.n218 source.t7 1.6505
R642 source.n218 source.t9 1.6505
R643 source.n216 source.t0 1.6505
R644 source.n216 source.t2 1.6505
R645 source.n148 source.t16 1.6505
R646 source.n148 source.t14 1.6505
R647 source.n146 source.t20 1.6505
R648 source.n146 source.t21 1.6505
R649 source.n144 source.t26 1.6505
R650 source.n144 source.t27 1.6505
R651 source.n66 source.t23 1.6505
R652 source.n66 source.t18 1.6505
R653 source.n68 source.t24 1.6505
R654 source.n68 source.t19 1.6505
R655 source.n70 source.t22 1.6505
R656 source.n70 source.t17 1.6505
R657 source.n138 source.t4 1.6505
R658 source.n138 source.t11 1.6505
R659 source.n140 source.t8 1.6505
R660 source.n140 source.t1 1.6505
R661 source.n142 source.t6 1.6505
R662 source.n142 source.t3 1.6505
R663 source.n263 source.n261 1.16414
R664 source.n271 source.n230 1.16414
R665 source.n191 source.n189 1.16414
R666 source.n199 source.n158 1.16414
R667 source.n49 source.n8 1.16414
R668 source.n41 source.n40 1.16414
R669 source.n121 source.n80 1.16414
R670 source.n113 source.n112 1.16414
R671 source.n137 source.n71 0.914293
R672 source.n217 source.n215 0.914293
R673 source.n143 source.n141 0.888431
R674 source.n141 source.n139 0.888431
R675 source.n139 source.n137 0.888431
R676 source.n71 source.n69 0.888431
R677 source.n69 source.n67 0.888431
R678 source.n67 source.n65 0.888431
R679 source.n147 source.n145 0.888431
R680 source.n149 source.n147 0.888431
R681 source.n215 source.n149 0.888431
R682 source.n219 source.n217 0.888431
R683 source.n221 source.n219 0.888431
R684 source.n287 source.n221 0.888431
R685 source.n262 source.n232 0.388379
R686 source.n268 source.n267 0.388379
R687 source.n190 source.n160 0.388379
R688 source.n196 source.n195 0.388379
R689 source.n46 source.n45 0.388379
R690 source.n12 source.n10 0.388379
R691 source.n118 source.n117 0.388379
R692 source.n84 source.n82 0.388379
R693 source source.n288 0.188
R694 source.n244 source.n239 0.155672
R695 source.n251 source.n239 0.155672
R696 source.n252 source.n251 0.155672
R697 source.n252 source.n235 0.155672
R698 source.n259 source.n235 0.155672
R699 source.n260 source.n259 0.155672
R700 source.n260 source.n231 0.155672
R701 source.n269 source.n231 0.155672
R702 source.n270 source.n269 0.155672
R703 source.n270 source.n227 0.155672
R704 source.n277 source.n227 0.155672
R705 source.n278 source.n277 0.155672
R706 source.n278 source.n223 0.155672
R707 source.n285 source.n223 0.155672
R708 source.n172 source.n167 0.155672
R709 source.n179 source.n167 0.155672
R710 source.n180 source.n179 0.155672
R711 source.n180 source.n163 0.155672
R712 source.n187 source.n163 0.155672
R713 source.n188 source.n187 0.155672
R714 source.n188 source.n159 0.155672
R715 source.n197 source.n159 0.155672
R716 source.n198 source.n197 0.155672
R717 source.n198 source.n155 0.155672
R718 source.n205 source.n155 0.155672
R719 source.n206 source.n205 0.155672
R720 source.n206 source.n151 0.155672
R721 source.n213 source.n151 0.155672
R722 source.n63 source.n1 0.155672
R723 source.n56 source.n1 0.155672
R724 source.n56 source.n55 0.155672
R725 source.n55 source.n5 0.155672
R726 source.n48 source.n5 0.155672
R727 source.n48 source.n47 0.155672
R728 source.n47 source.n9 0.155672
R729 source.n39 source.n9 0.155672
R730 source.n39 source.n38 0.155672
R731 source.n38 source.n14 0.155672
R732 source.n31 source.n14 0.155672
R733 source.n31 source.n30 0.155672
R734 source.n30 source.n18 0.155672
R735 source.n23 source.n18 0.155672
R736 source.n135 source.n73 0.155672
R737 source.n128 source.n73 0.155672
R738 source.n128 source.n127 0.155672
R739 source.n127 source.n77 0.155672
R740 source.n120 source.n77 0.155672
R741 source.n120 source.n119 0.155672
R742 source.n119 source.n81 0.155672
R743 source.n111 source.n81 0.155672
R744 source.n111 source.n110 0.155672
R745 source.n110 source.n86 0.155672
R746 source.n103 source.n86 0.155672
R747 source.n103 source.n102 0.155672
R748 source.n102 source.n90 0.155672
R749 source.n95 source.n90 0.155672
R750 minus.n5 minus.t6 493.108
R751 minus.n27 minus.t0 493.108
R752 minus.n6 minus.t1 469.262
R753 minus.n8 minus.t5 469.262
R754 minus.n12 minus.t11 469.262
R755 minus.n14 minus.t4 469.262
R756 minus.n18 minus.t12 469.262
R757 minus.n20 minus.t3 469.262
R758 minus.n28 minus.t2 469.262
R759 minus.n30 minus.t9 469.262
R760 minus.n34 minus.t10 469.262
R761 minus.n36 minus.t13 469.262
R762 minus.n40 minus.t7 469.262
R763 minus.n42 minus.t8 469.262
R764 minus.n21 minus.n20 161.3
R765 minus.n19 minus.n0 161.3
R766 minus.n18 minus.n17 161.3
R767 minus.n16 minus.n1 161.3
R768 minus.n15 minus.n14 161.3
R769 minus.n13 minus.n2 161.3
R770 minus.n12 minus.n11 161.3
R771 minus.n10 minus.n3 161.3
R772 minus.n9 minus.n8 161.3
R773 minus.n7 minus.n4 161.3
R774 minus.n43 minus.n42 161.3
R775 minus.n41 minus.n22 161.3
R776 minus.n40 minus.n39 161.3
R777 minus.n38 minus.n23 161.3
R778 minus.n37 minus.n36 161.3
R779 minus.n35 minus.n24 161.3
R780 minus.n34 minus.n33 161.3
R781 minus.n32 minus.n25 161.3
R782 minus.n31 minus.n30 161.3
R783 minus.n29 minus.n26 161.3
R784 minus.n5 minus.n4 44.9119
R785 minus.n27 minus.n26 44.9119
R786 minus.n44 minus.n21 38.2259
R787 minus.n20 minus.n19 35.055
R788 minus.n42 minus.n41 35.055
R789 minus.n7 minus.n6 30.6732
R790 minus.n18 minus.n1 30.6732
R791 minus.n29 minus.n28 30.6732
R792 minus.n40 minus.n23 30.6732
R793 minus.n8 minus.n3 26.2914
R794 minus.n14 minus.n13 26.2914
R795 minus.n30 minus.n25 26.2914
R796 minus.n36 minus.n35 26.2914
R797 minus.n12 minus.n3 21.9096
R798 minus.n13 minus.n12 21.9096
R799 minus.n34 minus.n25 21.9096
R800 minus.n35 minus.n34 21.9096
R801 minus.n6 minus.n5 17.739
R802 minus.n28 minus.n27 17.739
R803 minus.n8 minus.n7 17.5278
R804 minus.n14 minus.n1 17.5278
R805 minus.n30 minus.n29 17.5278
R806 minus.n36 minus.n23 17.5278
R807 minus.n19 minus.n18 13.146
R808 minus.n41 minus.n40 13.146
R809 minus.n44 minus.n43 6.65012
R810 minus.n21 minus.n0 0.189894
R811 minus.n17 minus.n0 0.189894
R812 minus.n17 minus.n16 0.189894
R813 minus.n16 minus.n15 0.189894
R814 minus.n15 minus.n2 0.189894
R815 minus.n11 minus.n2 0.189894
R816 minus.n11 minus.n10 0.189894
R817 minus.n10 minus.n9 0.189894
R818 minus.n9 minus.n4 0.189894
R819 minus.n31 minus.n26 0.189894
R820 minus.n32 minus.n31 0.189894
R821 minus.n33 minus.n32 0.189894
R822 minus.n33 minus.n24 0.189894
R823 minus.n37 minus.n24 0.189894
R824 minus.n38 minus.n37 0.189894
R825 minus.n39 minus.n38 0.189894
R826 minus.n39 minus.n22 0.189894
R827 minus.n43 minus.n22 0.189894
R828 minus minus.n44 0.188
R829 drain_right.n60 drain_right.n0 289.615
R830 drain_right.n136 drain_right.n76 289.615
R831 drain_right.n20 drain_right.n19 185
R832 drain_right.n25 drain_right.n24 185
R833 drain_right.n27 drain_right.n26 185
R834 drain_right.n16 drain_right.n15 185
R835 drain_right.n33 drain_right.n32 185
R836 drain_right.n35 drain_right.n34 185
R837 drain_right.n12 drain_right.n11 185
R838 drain_right.n42 drain_right.n41 185
R839 drain_right.n43 drain_right.n10 185
R840 drain_right.n45 drain_right.n44 185
R841 drain_right.n8 drain_right.n7 185
R842 drain_right.n51 drain_right.n50 185
R843 drain_right.n53 drain_right.n52 185
R844 drain_right.n4 drain_right.n3 185
R845 drain_right.n59 drain_right.n58 185
R846 drain_right.n61 drain_right.n60 185
R847 drain_right.n137 drain_right.n136 185
R848 drain_right.n135 drain_right.n134 185
R849 drain_right.n80 drain_right.n79 185
R850 drain_right.n129 drain_right.n128 185
R851 drain_right.n127 drain_right.n126 185
R852 drain_right.n84 drain_right.n83 185
R853 drain_right.n121 drain_right.n120 185
R854 drain_right.n119 drain_right.n86 185
R855 drain_right.n118 drain_right.n117 185
R856 drain_right.n89 drain_right.n87 185
R857 drain_right.n112 drain_right.n111 185
R858 drain_right.n110 drain_right.n109 185
R859 drain_right.n93 drain_right.n92 185
R860 drain_right.n104 drain_right.n103 185
R861 drain_right.n102 drain_right.n101 185
R862 drain_right.n97 drain_right.n96 185
R863 drain_right.n21 drain_right.t13 149.524
R864 drain_right.n98 drain_right.t10 149.524
R865 drain_right.n25 drain_right.n19 104.615
R866 drain_right.n26 drain_right.n25 104.615
R867 drain_right.n26 drain_right.n15 104.615
R868 drain_right.n33 drain_right.n15 104.615
R869 drain_right.n34 drain_right.n33 104.615
R870 drain_right.n34 drain_right.n11 104.615
R871 drain_right.n42 drain_right.n11 104.615
R872 drain_right.n43 drain_right.n42 104.615
R873 drain_right.n44 drain_right.n43 104.615
R874 drain_right.n44 drain_right.n7 104.615
R875 drain_right.n51 drain_right.n7 104.615
R876 drain_right.n52 drain_right.n51 104.615
R877 drain_right.n52 drain_right.n3 104.615
R878 drain_right.n59 drain_right.n3 104.615
R879 drain_right.n60 drain_right.n59 104.615
R880 drain_right.n136 drain_right.n135 104.615
R881 drain_right.n135 drain_right.n79 104.615
R882 drain_right.n128 drain_right.n79 104.615
R883 drain_right.n128 drain_right.n127 104.615
R884 drain_right.n127 drain_right.n83 104.615
R885 drain_right.n120 drain_right.n83 104.615
R886 drain_right.n120 drain_right.n119 104.615
R887 drain_right.n119 drain_right.n118 104.615
R888 drain_right.n118 drain_right.n87 104.615
R889 drain_right.n111 drain_right.n87 104.615
R890 drain_right.n111 drain_right.n110 104.615
R891 drain_right.n110 drain_right.n92 104.615
R892 drain_right.n103 drain_right.n92 104.615
R893 drain_right.n103 drain_right.n102 104.615
R894 drain_right.n102 drain_right.n96 104.615
R895 drain_right.n69 drain_right.n67 60.4404
R896 drain_right.n73 drain_right.n71 60.4404
R897 drain_right.n73 drain_right.n72 59.5527
R898 drain_right.n75 drain_right.n74 59.5527
R899 drain_right.n69 drain_right.n68 59.5525
R900 drain_right.n66 drain_right.n65 59.5525
R901 drain_right.t13 drain_right.n19 52.3082
R902 drain_right.t10 drain_right.n96 52.3082
R903 drain_right.n66 drain_right.n64 47.4248
R904 drain_right.n141 drain_right.n140 46.5369
R905 drain_right drain_right.n70 31.9194
R906 drain_right.n45 drain_right.n10 13.1884
R907 drain_right.n121 drain_right.n86 13.1884
R908 drain_right.n41 drain_right.n40 12.8005
R909 drain_right.n46 drain_right.n8 12.8005
R910 drain_right.n122 drain_right.n84 12.8005
R911 drain_right.n117 drain_right.n88 12.8005
R912 drain_right.n39 drain_right.n12 12.0247
R913 drain_right.n50 drain_right.n49 12.0247
R914 drain_right.n126 drain_right.n125 12.0247
R915 drain_right.n116 drain_right.n89 12.0247
R916 drain_right.n36 drain_right.n35 11.249
R917 drain_right.n53 drain_right.n6 11.249
R918 drain_right.n129 drain_right.n82 11.249
R919 drain_right.n113 drain_right.n112 11.249
R920 drain_right.n32 drain_right.n14 10.4732
R921 drain_right.n54 drain_right.n4 10.4732
R922 drain_right.n130 drain_right.n80 10.4732
R923 drain_right.n109 drain_right.n91 10.4732
R924 drain_right.n21 drain_right.n20 10.2747
R925 drain_right.n98 drain_right.n97 10.2747
R926 drain_right.n31 drain_right.n16 9.69747
R927 drain_right.n58 drain_right.n57 9.69747
R928 drain_right.n134 drain_right.n133 9.69747
R929 drain_right.n108 drain_right.n93 9.69747
R930 drain_right.n64 drain_right.n63 9.45567
R931 drain_right.n140 drain_right.n139 9.45567
R932 drain_right.n63 drain_right.n62 9.3005
R933 drain_right.n2 drain_right.n1 9.3005
R934 drain_right.n57 drain_right.n56 9.3005
R935 drain_right.n55 drain_right.n54 9.3005
R936 drain_right.n6 drain_right.n5 9.3005
R937 drain_right.n49 drain_right.n48 9.3005
R938 drain_right.n47 drain_right.n46 9.3005
R939 drain_right.n23 drain_right.n22 9.3005
R940 drain_right.n18 drain_right.n17 9.3005
R941 drain_right.n29 drain_right.n28 9.3005
R942 drain_right.n31 drain_right.n30 9.3005
R943 drain_right.n14 drain_right.n13 9.3005
R944 drain_right.n37 drain_right.n36 9.3005
R945 drain_right.n39 drain_right.n38 9.3005
R946 drain_right.n40 drain_right.n9 9.3005
R947 drain_right.n100 drain_right.n99 9.3005
R948 drain_right.n95 drain_right.n94 9.3005
R949 drain_right.n106 drain_right.n105 9.3005
R950 drain_right.n108 drain_right.n107 9.3005
R951 drain_right.n91 drain_right.n90 9.3005
R952 drain_right.n114 drain_right.n113 9.3005
R953 drain_right.n116 drain_right.n115 9.3005
R954 drain_right.n88 drain_right.n85 9.3005
R955 drain_right.n139 drain_right.n138 9.3005
R956 drain_right.n78 drain_right.n77 9.3005
R957 drain_right.n133 drain_right.n132 9.3005
R958 drain_right.n131 drain_right.n130 9.3005
R959 drain_right.n82 drain_right.n81 9.3005
R960 drain_right.n125 drain_right.n124 9.3005
R961 drain_right.n123 drain_right.n122 9.3005
R962 drain_right.n28 drain_right.n27 8.92171
R963 drain_right.n61 drain_right.n2 8.92171
R964 drain_right.n137 drain_right.n78 8.92171
R965 drain_right.n105 drain_right.n104 8.92171
R966 drain_right.n24 drain_right.n18 8.14595
R967 drain_right.n62 drain_right.n0 8.14595
R968 drain_right.n138 drain_right.n76 8.14595
R969 drain_right.n101 drain_right.n95 8.14595
R970 drain_right.n23 drain_right.n20 7.3702
R971 drain_right.n100 drain_right.n97 7.3702
R972 drain_right drain_right.n141 6.09718
R973 drain_right.n24 drain_right.n23 5.81868
R974 drain_right.n64 drain_right.n0 5.81868
R975 drain_right.n140 drain_right.n76 5.81868
R976 drain_right.n101 drain_right.n100 5.81868
R977 drain_right.n27 drain_right.n18 5.04292
R978 drain_right.n62 drain_right.n61 5.04292
R979 drain_right.n138 drain_right.n137 5.04292
R980 drain_right.n104 drain_right.n95 5.04292
R981 drain_right.n28 drain_right.n16 4.26717
R982 drain_right.n58 drain_right.n2 4.26717
R983 drain_right.n134 drain_right.n78 4.26717
R984 drain_right.n105 drain_right.n93 4.26717
R985 drain_right.n32 drain_right.n31 3.49141
R986 drain_right.n57 drain_right.n4 3.49141
R987 drain_right.n133 drain_right.n80 3.49141
R988 drain_right.n109 drain_right.n108 3.49141
R989 drain_right.n22 drain_right.n21 2.84303
R990 drain_right.n99 drain_right.n98 2.84303
R991 drain_right.n35 drain_right.n14 2.71565
R992 drain_right.n54 drain_right.n53 2.71565
R993 drain_right.n130 drain_right.n129 2.71565
R994 drain_right.n112 drain_right.n91 2.71565
R995 drain_right.n36 drain_right.n12 1.93989
R996 drain_right.n50 drain_right.n6 1.93989
R997 drain_right.n126 drain_right.n82 1.93989
R998 drain_right.n113 drain_right.n89 1.93989
R999 drain_right.n67 drain_right.t6 1.6505
R1000 drain_right.n67 drain_right.t5 1.6505
R1001 drain_right.n68 drain_right.t3 1.6505
R1002 drain_right.n68 drain_right.t0 1.6505
R1003 drain_right.n65 drain_right.t11 1.6505
R1004 drain_right.n65 drain_right.t4 1.6505
R1005 drain_right.n71 drain_right.t12 1.6505
R1006 drain_right.n71 drain_right.t7 1.6505
R1007 drain_right.n72 drain_right.t2 1.6505
R1008 drain_right.n72 drain_right.t8 1.6505
R1009 drain_right.n74 drain_right.t1 1.6505
R1010 drain_right.n74 drain_right.t9 1.6505
R1011 drain_right.n41 drain_right.n39 1.16414
R1012 drain_right.n49 drain_right.n8 1.16414
R1013 drain_right.n125 drain_right.n84 1.16414
R1014 drain_right.n117 drain_right.n116 1.16414
R1015 drain_right.n141 drain_right.n75 0.888431
R1016 drain_right.n75 drain_right.n73 0.888431
R1017 drain_right.n70 drain_right.n66 0.611102
R1018 drain_right.n40 drain_right.n10 0.388379
R1019 drain_right.n46 drain_right.n45 0.388379
R1020 drain_right.n122 drain_right.n121 0.388379
R1021 drain_right.n88 drain_right.n86 0.388379
R1022 drain_right.n70 drain_right.n69 0.167137
R1023 drain_right.n22 drain_right.n17 0.155672
R1024 drain_right.n29 drain_right.n17 0.155672
R1025 drain_right.n30 drain_right.n29 0.155672
R1026 drain_right.n30 drain_right.n13 0.155672
R1027 drain_right.n37 drain_right.n13 0.155672
R1028 drain_right.n38 drain_right.n37 0.155672
R1029 drain_right.n38 drain_right.n9 0.155672
R1030 drain_right.n47 drain_right.n9 0.155672
R1031 drain_right.n48 drain_right.n47 0.155672
R1032 drain_right.n48 drain_right.n5 0.155672
R1033 drain_right.n55 drain_right.n5 0.155672
R1034 drain_right.n56 drain_right.n55 0.155672
R1035 drain_right.n56 drain_right.n1 0.155672
R1036 drain_right.n63 drain_right.n1 0.155672
R1037 drain_right.n139 drain_right.n77 0.155672
R1038 drain_right.n132 drain_right.n77 0.155672
R1039 drain_right.n132 drain_right.n131 0.155672
R1040 drain_right.n131 drain_right.n81 0.155672
R1041 drain_right.n124 drain_right.n81 0.155672
R1042 drain_right.n124 drain_right.n123 0.155672
R1043 drain_right.n123 drain_right.n85 0.155672
R1044 drain_right.n115 drain_right.n85 0.155672
R1045 drain_right.n115 drain_right.n114 0.155672
R1046 drain_right.n114 drain_right.n90 0.155672
R1047 drain_right.n107 drain_right.n90 0.155672
R1048 drain_right.n107 drain_right.n106 0.155672
R1049 drain_right.n106 drain_right.n94 0.155672
R1050 drain_right.n99 drain_right.n94 0.155672
C0 drain_right drain_left 1.23389f
C1 drain_right source 18.639198f
C2 drain_left minus 0.172675f
C3 drain_right plus 0.39102f
C4 minus source 9.0289f
C5 minus plus 6.09248f
C6 drain_right minus 9.06606f
C7 drain_left source 18.6455f
C8 drain_left plus 9.296901f
C9 plus source 9.043441f
C10 drain_right a_n2364_n3288# 7.55399f
C11 drain_left a_n2364_n3288# 7.904f
C12 source a_n2364_n3288# 6.674157f
C13 minus a_n2364_n3288# 9.382834f
C14 plus a_n2364_n3288# 11.10981f
C15 drain_right.n0 a_n2364_n3288# 0.033044f
C16 drain_right.n1 a_n2364_n3288# 0.024946f
C17 drain_right.n2 a_n2364_n3288# 0.013405f
C18 drain_right.n3 a_n2364_n3288# 0.031684f
C19 drain_right.n4 a_n2364_n3288# 0.014193f
C20 drain_right.n5 a_n2364_n3288# 0.024946f
C21 drain_right.n6 a_n2364_n3288# 0.013405f
C22 drain_right.n7 a_n2364_n3288# 0.031684f
C23 drain_right.n8 a_n2364_n3288# 0.014193f
C24 drain_right.n9 a_n2364_n3288# 0.024946f
C25 drain_right.n10 a_n2364_n3288# 0.013799f
C26 drain_right.n11 a_n2364_n3288# 0.031684f
C27 drain_right.n12 a_n2364_n3288# 0.014193f
C28 drain_right.n13 a_n2364_n3288# 0.024946f
C29 drain_right.n14 a_n2364_n3288# 0.013405f
C30 drain_right.n15 a_n2364_n3288# 0.031684f
C31 drain_right.n16 a_n2364_n3288# 0.014193f
C32 drain_right.n17 a_n2364_n3288# 0.024946f
C33 drain_right.n18 a_n2364_n3288# 0.013405f
C34 drain_right.n19 a_n2364_n3288# 0.023763f
C35 drain_right.n20 a_n2364_n3288# 0.022398f
C36 drain_right.t13 a_n2364_n3288# 0.053513f
C37 drain_right.n21 a_n2364_n3288# 0.179857f
C38 drain_right.n22 a_n2364_n3288# 1.25848f
C39 drain_right.n23 a_n2364_n3288# 0.013405f
C40 drain_right.n24 a_n2364_n3288# 0.014193f
C41 drain_right.n25 a_n2364_n3288# 0.031684f
C42 drain_right.n26 a_n2364_n3288# 0.031684f
C43 drain_right.n27 a_n2364_n3288# 0.014193f
C44 drain_right.n28 a_n2364_n3288# 0.013405f
C45 drain_right.n29 a_n2364_n3288# 0.024946f
C46 drain_right.n30 a_n2364_n3288# 0.024946f
C47 drain_right.n31 a_n2364_n3288# 0.013405f
C48 drain_right.n32 a_n2364_n3288# 0.014193f
C49 drain_right.n33 a_n2364_n3288# 0.031684f
C50 drain_right.n34 a_n2364_n3288# 0.031684f
C51 drain_right.n35 a_n2364_n3288# 0.014193f
C52 drain_right.n36 a_n2364_n3288# 0.013405f
C53 drain_right.n37 a_n2364_n3288# 0.024946f
C54 drain_right.n38 a_n2364_n3288# 0.024946f
C55 drain_right.n39 a_n2364_n3288# 0.013405f
C56 drain_right.n40 a_n2364_n3288# 0.013405f
C57 drain_right.n41 a_n2364_n3288# 0.014193f
C58 drain_right.n42 a_n2364_n3288# 0.031684f
C59 drain_right.n43 a_n2364_n3288# 0.031684f
C60 drain_right.n44 a_n2364_n3288# 0.031684f
C61 drain_right.n45 a_n2364_n3288# 0.013799f
C62 drain_right.n46 a_n2364_n3288# 0.013405f
C63 drain_right.n47 a_n2364_n3288# 0.024946f
C64 drain_right.n48 a_n2364_n3288# 0.024946f
C65 drain_right.n49 a_n2364_n3288# 0.013405f
C66 drain_right.n50 a_n2364_n3288# 0.014193f
C67 drain_right.n51 a_n2364_n3288# 0.031684f
C68 drain_right.n52 a_n2364_n3288# 0.031684f
C69 drain_right.n53 a_n2364_n3288# 0.014193f
C70 drain_right.n54 a_n2364_n3288# 0.013405f
C71 drain_right.n55 a_n2364_n3288# 0.024946f
C72 drain_right.n56 a_n2364_n3288# 0.024946f
C73 drain_right.n57 a_n2364_n3288# 0.013405f
C74 drain_right.n58 a_n2364_n3288# 0.014193f
C75 drain_right.n59 a_n2364_n3288# 0.031684f
C76 drain_right.n60 a_n2364_n3288# 0.065019f
C77 drain_right.n61 a_n2364_n3288# 0.014193f
C78 drain_right.n62 a_n2364_n3288# 0.013405f
C79 drain_right.n63 a_n2364_n3288# 0.053572f
C80 drain_right.n64 a_n2364_n3288# 0.055336f
C81 drain_right.t11 a_n2364_n3288# 0.236557f
C82 drain_right.t4 a_n2364_n3288# 0.236557f
C83 drain_right.n65 a_n2364_n3288# 2.10499f
C84 drain_right.n66 a_n2364_n3288# 0.445639f
C85 drain_right.t6 a_n2364_n3288# 0.236557f
C86 drain_right.t5 a_n2364_n3288# 0.236557f
C87 drain_right.n67 a_n2364_n3288# 2.11031f
C88 drain_right.t3 a_n2364_n3288# 0.236557f
C89 drain_right.t0 a_n2364_n3288# 0.236557f
C90 drain_right.n68 a_n2364_n3288# 2.10499f
C91 drain_right.n69 a_n2364_n3288# 0.654432f
C92 drain_right.n70 a_n2364_n3288# 1.32641f
C93 drain_right.t12 a_n2364_n3288# 0.236557f
C94 drain_right.t7 a_n2364_n3288# 0.236557f
C95 drain_right.n71 a_n2364_n3288# 2.11031f
C96 drain_right.t2 a_n2364_n3288# 0.236557f
C97 drain_right.t8 a_n2364_n3288# 0.236557f
C98 drain_right.n72 a_n2364_n3288# 2.105f
C99 drain_right.n73 a_n2364_n3288# 0.708932f
C100 drain_right.t1 a_n2364_n3288# 0.236557f
C101 drain_right.t9 a_n2364_n3288# 0.236557f
C102 drain_right.n74 a_n2364_n3288# 2.105f
C103 drain_right.n75 a_n2364_n3288# 0.352098f
C104 drain_right.n76 a_n2364_n3288# 0.033044f
C105 drain_right.n77 a_n2364_n3288# 0.024946f
C106 drain_right.n78 a_n2364_n3288# 0.013405f
C107 drain_right.n79 a_n2364_n3288# 0.031684f
C108 drain_right.n80 a_n2364_n3288# 0.014193f
C109 drain_right.n81 a_n2364_n3288# 0.024946f
C110 drain_right.n82 a_n2364_n3288# 0.013405f
C111 drain_right.n83 a_n2364_n3288# 0.031684f
C112 drain_right.n84 a_n2364_n3288# 0.014193f
C113 drain_right.n85 a_n2364_n3288# 0.024946f
C114 drain_right.n86 a_n2364_n3288# 0.013799f
C115 drain_right.n87 a_n2364_n3288# 0.031684f
C116 drain_right.n88 a_n2364_n3288# 0.013405f
C117 drain_right.n89 a_n2364_n3288# 0.014193f
C118 drain_right.n90 a_n2364_n3288# 0.024946f
C119 drain_right.n91 a_n2364_n3288# 0.013405f
C120 drain_right.n92 a_n2364_n3288# 0.031684f
C121 drain_right.n93 a_n2364_n3288# 0.014193f
C122 drain_right.n94 a_n2364_n3288# 0.024946f
C123 drain_right.n95 a_n2364_n3288# 0.013405f
C124 drain_right.n96 a_n2364_n3288# 0.023763f
C125 drain_right.n97 a_n2364_n3288# 0.022398f
C126 drain_right.t10 a_n2364_n3288# 0.053513f
C127 drain_right.n98 a_n2364_n3288# 0.179857f
C128 drain_right.n99 a_n2364_n3288# 1.25848f
C129 drain_right.n100 a_n2364_n3288# 0.013405f
C130 drain_right.n101 a_n2364_n3288# 0.014193f
C131 drain_right.n102 a_n2364_n3288# 0.031684f
C132 drain_right.n103 a_n2364_n3288# 0.031684f
C133 drain_right.n104 a_n2364_n3288# 0.014193f
C134 drain_right.n105 a_n2364_n3288# 0.013405f
C135 drain_right.n106 a_n2364_n3288# 0.024946f
C136 drain_right.n107 a_n2364_n3288# 0.024946f
C137 drain_right.n108 a_n2364_n3288# 0.013405f
C138 drain_right.n109 a_n2364_n3288# 0.014193f
C139 drain_right.n110 a_n2364_n3288# 0.031684f
C140 drain_right.n111 a_n2364_n3288# 0.031684f
C141 drain_right.n112 a_n2364_n3288# 0.014193f
C142 drain_right.n113 a_n2364_n3288# 0.013405f
C143 drain_right.n114 a_n2364_n3288# 0.024946f
C144 drain_right.n115 a_n2364_n3288# 0.024946f
C145 drain_right.n116 a_n2364_n3288# 0.013405f
C146 drain_right.n117 a_n2364_n3288# 0.014193f
C147 drain_right.n118 a_n2364_n3288# 0.031684f
C148 drain_right.n119 a_n2364_n3288# 0.031684f
C149 drain_right.n120 a_n2364_n3288# 0.031684f
C150 drain_right.n121 a_n2364_n3288# 0.013799f
C151 drain_right.n122 a_n2364_n3288# 0.013405f
C152 drain_right.n123 a_n2364_n3288# 0.024946f
C153 drain_right.n124 a_n2364_n3288# 0.024946f
C154 drain_right.n125 a_n2364_n3288# 0.013405f
C155 drain_right.n126 a_n2364_n3288# 0.014193f
C156 drain_right.n127 a_n2364_n3288# 0.031684f
C157 drain_right.n128 a_n2364_n3288# 0.031684f
C158 drain_right.n129 a_n2364_n3288# 0.014193f
C159 drain_right.n130 a_n2364_n3288# 0.013405f
C160 drain_right.n131 a_n2364_n3288# 0.024946f
C161 drain_right.n132 a_n2364_n3288# 0.024946f
C162 drain_right.n133 a_n2364_n3288# 0.013405f
C163 drain_right.n134 a_n2364_n3288# 0.014193f
C164 drain_right.n135 a_n2364_n3288# 0.031684f
C165 drain_right.n136 a_n2364_n3288# 0.065019f
C166 drain_right.n137 a_n2364_n3288# 0.014193f
C167 drain_right.n138 a_n2364_n3288# 0.013405f
C168 drain_right.n139 a_n2364_n3288# 0.053572f
C169 drain_right.n140 a_n2364_n3288# 0.053144f
C170 drain_right.n141 a_n2364_n3288# 0.346336f
C171 minus.n0 a_n2364_n3288# 0.041108f
C172 minus.n1 a_n2364_n3288# 0.009328f
C173 minus.t12 a_n2364_n3288# 0.984654f
C174 minus.n2 a_n2364_n3288# 0.041108f
C175 minus.n3 a_n2364_n3288# 0.009328f
C176 minus.t11 a_n2364_n3288# 0.984654f
C177 minus.n4 a_n2364_n3288# 0.173207f
C178 minus.t6 a_n2364_n3288# 1.00365f
C179 minus.n5 a_n2364_n3288# 0.377279f
C180 minus.t1 a_n2364_n3288# 0.984654f
C181 minus.n6 a_n2364_n3288# 0.397791f
C182 minus.n7 a_n2364_n3288# 0.009328f
C183 minus.t5 a_n2364_n3288# 0.984654f
C184 minus.n8 a_n2364_n3288# 0.392699f
C185 minus.n9 a_n2364_n3288# 0.041108f
C186 minus.n10 a_n2364_n3288# 0.041108f
C187 minus.n11 a_n2364_n3288# 0.041108f
C188 minus.n12 a_n2364_n3288# 0.392699f
C189 minus.n13 a_n2364_n3288# 0.009328f
C190 minus.t4 a_n2364_n3288# 0.984654f
C191 minus.n14 a_n2364_n3288# 0.392699f
C192 minus.n15 a_n2364_n3288# 0.041108f
C193 minus.n16 a_n2364_n3288# 0.041108f
C194 minus.n17 a_n2364_n3288# 0.041108f
C195 minus.n18 a_n2364_n3288# 0.392699f
C196 minus.n19 a_n2364_n3288# 0.009328f
C197 minus.t3 a_n2364_n3288# 0.984654f
C198 minus.n20 a_n2364_n3288# 0.391178f
C199 minus.n21 a_n2364_n3288# 1.5853f
C200 minus.n22 a_n2364_n3288# 0.041108f
C201 minus.n23 a_n2364_n3288# 0.009328f
C202 minus.n24 a_n2364_n3288# 0.041108f
C203 minus.n25 a_n2364_n3288# 0.009328f
C204 minus.n26 a_n2364_n3288# 0.173207f
C205 minus.t0 a_n2364_n3288# 1.00365f
C206 minus.n27 a_n2364_n3288# 0.377279f
C207 minus.t2 a_n2364_n3288# 0.984654f
C208 minus.n28 a_n2364_n3288# 0.397791f
C209 minus.n29 a_n2364_n3288# 0.009328f
C210 minus.t9 a_n2364_n3288# 0.984654f
C211 minus.n30 a_n2364_n3288# 0.392699f
C212 minus.n31 a_n2364_n3288# 0.041108f
C213 minus.n32 a_n2364_n3288# 0.041108f
C214 minus.n33 a_n2364_n3288# 0.041108f
C215 minus.t10 a_n2364_n3288# 0.984654f
C216 minus.n34 a_n2364_n3288# 0.392699f
C217 minus.n35 a_n2364_n3288# 0.009328f
C218 minus.t13 a_n2364_n3288# 0.984654f
C219 minus.n36 a_n2364_n3288# 0.392699f
C220 minus.n37 a_n2364_n3288# 0.041108f
C221 minus.n38 a_n2364_n3288# 0.041108f
C222 minus.n39 a_n2364_n3288# 0.041108f
C223 minus.t7 a_n2364_n3288# 0.984654f
C224 minus.n40 a_n2364_n3288# 0.392699f
C225 minus.n41 a_n2364_n3288# 0.009328f
C226 minus.t8 a_n2364_n3288# 0.984654f
C227 minus.n42 a_n2364_n3288# 0.391178f
C228 minus.n43 a_n2364_n3288# 0.283193f
C229 minus.n44 a_n2364_n3288# 1.90985f
C230 source.n0 a_n2364_n3288# 0.03481f
C231 source.n1 a_n2364_n3288# 0.026279f
C232 source.n2 a_n2364_n3288# 0.014121f
C233 source.n3 a_n2364_n3288# 0.033378f
C234 source.n4 a_n2364_n3288# 0.014952f
C235 source.n5 a_n2364_n3288# 0.026279f
C236 source.n6 a_n2364_n3288# 0.014121f
C237 source.n7 a_n2364_n3288# 0.033378f
C238 source.n8 a_n2364_n3288# 0.014952f
C239 source.n9 a_n2364_n3288# 0.026279f
C240 source.n10 a_n2364_n3288# 0.014537f
C241 source.n11 a_n2364_n3288# 0.033378f
C242 source.n12 a_n2364_n3288# 0.014121f
C243 source.n13 a_n2364_n3288# 0.014952f
C244 source.n14 a_n2364_n3288# 0.026279f
C245 source.n15 a_n2364_n3288# 0.014121f
C246 source.n16 a_n2364_n3288# 0.033378f
C247 source.n17 a_n2364_n3288# 0.014952f
C248 source.n18 a_n2364_n3288# 0.026279f
C249 source.n19 a_n2364_n3288# 0.014121f
C250 source.n20 a_n2364_n3288# 0.025033f
C251 source.n21 a_n2364_n3288# 0.023596f
C252 source.t25 a_n2364_n3288# 0.056373f
C253 source.n22 a_n2364_n3288# 0.18947f
C254 source.n23 a_n2364_n3288# 1.32574f
C255 source.n24 a_n2364_n3288# 0.014121f
C256 source.n25 a_n2364_n3288# 0.014952f
C257 source.n26 a_n2364_n3288# 0.033378f
C258 source.n27 a_n2364_n3288# 0.033378f
C259 source.n28 a_n2364_n3288# 0.014952f
C260 source.n29 a_n2364_n3288# 0.014121f
C261 source.n30 a_n2364_n3288# 0.026279f
C262 source.n31 a_n2364_n3288# 0.026279f
C263 source.n32 a_n2364_n3288# 0.014121f
C264 source.n33 a_n2364_n3288# 0.014952f
C265 source.n34 a_n2364_n3288# 0.033378f
C266 source.n35 a_n2364_n3288# 0.033378f
C267 source.n36 a_n2364_n3288# 0.014952f
C268 source.n37 a_n2364_n3288# 0.014121f
C269 source.n38 a_n2364_n3288# 0.026279f
C270 source.n39 a_n2364_n3288# 0.026279f
C271 source.n40 a_n2364_n3288# 0.014121f
C272 source.n41 a_n2364_n3288# 0.014952f
C273 source.n42 a_n2364_n3288# 0.033378f
C274 source.n43 a_n2364_n3288# 0.033378f
C275 source.n44 a_n2364_n3288# 0.033378f
C276 source.n45 a_n2364_n3288# 0.014537f
C277 source.n46 a_n2364_n3288# 0.014121f
C278 source.n47 a_n2364_n3288# 0.026279f
C279 source.n48 a_n2364_n3288# 0.026279f
C280 source.n49 a_n2364_n3288# 0.014121f
C281 source.n50 a_n2364_n3288# 0.014952f
C282 source.n51 a_n2364_n3288# 0.033378f
C283 source.n52 a_n2364_n3288# 0.033378f
C284 source.n53 a_n2364_n3288# 0.014952f
C285 source.n54 a_n2364_n3288# 0.014121f
C286 source.n55 a_n2364_n3288# 0.026279f
C287 source.n56 a_n2364_n3288# 0.026279f
C288 source.n57 a_n2364_n3288# 0.014121f
C289 source.n58 a_n2364_n3288# 0.014952f
C290 source.n59 a_n2364_n3288# 0.033378f
C291 source.n60 a_n2364_n3288# 0.068495f
C292 source.n61 a_n2364_n3288# 0.014952f
C293 source.n62 a_n2364_n3288# 0.014121f
C294 source.n63 a_n2364_n3288# 0.056435f
C295 source.n64 a_n2364_n3288# 0.037802f
C296 source.n65 a_n2364_n3288# 1.10547f
C297 source.t23 a_n2364_n3288# 0.2492f
C298 source.t18 a_n2364_n3288# 0.2492f
C299 source.n66 a_n2364_n3288# 2.13366f
C300 source.n67 a_n2364_n3288# 0.419048f
C301 source.t24 a_n2364_n3288# 0.2492f
C302 source.t19 a_n2364_n3288# 0.2492f
C303 source.n68 a_n2364_n3288# 2.13366f
C304 source.n69 a_n2364_n3288# 0.419048f
C305 source.t22 a_n2364_n3288# 0.2492f
C306 source.t17 a_n2364_n3288# 0.2492f
C307 source.n70 a_n2364_n3288# 2.13366f
C308 source.n71 a_n2364_n3288# 0.421238f
C309 source.n72 a_n2364_n3288# 0.03481f
C310 source.n73 a_n2364_n3288# 0.026279f
C311 source.n74 a_n2364_n3288# 0.014121f
C312 source.n75 a_n2364_n3288# 0.033378f
C313 source.n76 a_n2364_n3288# 0.014952f
C314 source.n77 a_n2364_n3288# 0.026279f
C315 source.n78 a_n2364_n3288# 0.014121f
C316 source.n79 a_n2364_n3288# 0.033378f
C317 source.n80 a_n2364_n3288# 0.014952f
C318 source.n81 a_n2364_n3288# 0.026279f
C319 source.n82 a_n2364_n3288# 0.014537f
C320 source.n83 a_n2364_n3288# 0.033378f
C321 source.n84 a_n2364_n3288# 0.014121f
C322 source.n85 a_n2364_n3288# 0.014952f
C323 source.n86 a_n2364_n3288# 0.026279f
C324 source.n87 a_n2364_n3288# 0.014121f
C325 source.n88 a_n2364_n3288# 0.033378f
C326 source.n89 a_n2364_n3288# 0.014952f
C327 source.n90 a_n2364_n3288# 0.026279f
C328 source.n91 a_n2364_n3288# 0.014121f
C329 source.n92 a_n2364_n3288# 0.025033f
C330 source.n93 a_n2364_n3288# 0.023596f
C331 source.t13 a_n2364_n3288# 0.056373f
C332 source.n94 a_n2364_n3288# 0.18947f
C333 source.n95 a_n2364_n3288# 1.32574f
C334 source.n96 a_n2364_n3288# 0.014121f
C335 source.n97 a_n2364_n3288# 0.014952f
C336 source.n98 a_n2364_n3288# 0.033378f
C337 source.n99 a_n2364_n3288# 0.033378f
C338 source.n100 a_n2364_n3288# 0.014952f
C339 source.n101 a_n2364_n3288# 0.014121f
C340 source.n102 a_n2364_n3288# 0.026279f
C341 source.n103 a_n2364_n3288# 0.026279f
C342 source.n104 a_n2364_n3288# 0.014121f
C343 source.n105 a_n2364_n3288# 0.014952f
C344 source.n106 a_n2364_n3288# 0.033378f
C345 source.n107 a_n2364_n3288# 0.033378f
C346 source.n108 a_n2364_n3288# 0.014952f
C347 source.n109 a_n2364_n3288# 0.014121f
C348 source.n110 a_n2364_n3288# 0.026279f
C349 source.n111 a_n2364_n3288# 0.026279f
C350 source.n112 a_n2364_n3288# 0.014121f
C351 source.n113 a_n2364_n3288# 0.014952f
C352 source.n114 a_n2364_n3288# 0.033378f
C353 source.n115 a_n2364_n3288# 0.033378f
C354 source.n116 a_n2364_n3288# 0.033378f
C355 source.n117 a_n2364_n3288# 0.014537f
C356 source.n118 a_n2364_n3288# 0.014121f
C357 source.n119 a_n2364_n3288# 0.026279f
C358 source.n120 a_n2364_n3288# 0.026279f
C359 source.n121 a_n2364_n3288# 0.014121f
C360 source.n122 a_n2364_n3288# 0.014952f
C361 source.n123 a_n2364_n3288# 0.033378f
C362 source.n124 a_n2364_n3288# 0.033378f
C363 source.n125 a_n2364_n3288# 0.014952f
C364 source.n126 a_n2364_n3288# 0.014121f
C365 source.n127 a_n2364_n3288# 0.026279f
C366 source.n128 a_n2364_n3288# 0.026279f
C367 source.n129 a_n2364_n3288# 0.014121f
C368 source.n130 a_n2364_n3288# 0.014952f
C369 source.n131 a_n2364_n3288# 0.033378f
C370 source.n132 a_n2364_n3288# 0.068495f
C371 source.n133 a_n2364_n3288# 0.014952f
C372 source.n134 a_n2364_n3288# 0.014121f
C373 source.n135 a_n2364_n3288# 0.056435f
C374 source.n136 a_n2364_n3288# 0.037802f
C375 source.n137 a_n2364_n3288# 0.172583f
C376 source.t4 a_n2364_n3288# 0.2492f
C377 source.t11 a_n2364_n3288# 0.2492f
C378 source.n138 a_n2364_n3288# 2.13366f
C379 source.n139 a_n2364_n3288# 0.419048f
C380 source.t8 a_n2364_n3288# 0.2492f
C381 source.t1 a_n2364_n3288# 0.2492f
C382 source.n140 a_n2364_n3288# 2.13366f
C383 source.n141 a_n2364_n3288# 0.419048f
C384 source.t6 a_n2364_n3288# 0.2492f
C385 source.t3 a_n2364_n3288# 0.2492f
C386 source.n142 a_n2364_n3288# 2.13366f
C387 source.n143 a_n2364_n3288# 1.85307f
C388 source.t26 a_n2364_n3288# 0.2492f
C389 source.t27 a_n2364_n3288# 0.2492f
C390 source.n144 a_n2364_n3288# 2.13364f
C391 source.n145 a_n2364_n3288# 1.85308f
C392 source.t20 a_n2364_n3288# 0.2492f
C393 source.t21 a_n2364_n3288# 0.2492f
C394 source.n146 a_n2364_n3288# 2.13364f
C395 source.n147 a_n2364_n3288# 0.419061f
C396 source.t16 a_n2364_n3288# 0.2492f
C397 source.t14 a_n2364_n3288# 0.2492f
C398 source.n148 a_n2364_n3288# 2.13364f
C399 source.n149 a_n2364_n3288# 0.419061f
C400 source.n150 a_n2364_n3288# 0.03481f
C401 source.n151 a_n2364_n3288# 0.026279f
C402 source.n152 a_n2364_n3288# 0.014121f
C403 source.n153 a_n2364_n3288# 0.033378f
C404 source.n154 a_n2364_n3288# 0.014952f
C405 source.n155 a_n2364_n3288# 0.026279f
C406 source.n156 a_n2364_n3288# 0.014121f
C407 source.n157 a_n2364_n3288# 0.033378f
C408 source.n158 a_n2364_n3288# 0.014952f
C409 source.n159 a_n2364_n3288# 0.026279f
C410 source.n160 a_n2364_n3288# 0.014537f
C411 source.n161 a_n2364_n3288# 0.033378f
C412 source.n162 a_n2364_n3288# 0.014952f
C413 source.n163 a_n2364_n3288# 0.026279f
C414 source.n164 a_n2364_n3288# 0.014121f
C415 source.n165 a_n2364_n3288# 0.033378f
C416 source.n166 a_n2364_n3288# 0.014952f
C417 source.n167 a_n2364_n3288# 0.026279f
C418 source.n168 a_n2364_n3288# 0.014121f
C419 source.n169 a_n2364_n3288# 0.025033f
C420 source.n170 a_n2364_n3288# 0.023596f
C421 source.t15 a_n2364_n3288# 0.056373f
C422 source.n171 a_n2364_n3288# 0.18947f
C423 source.n172 a_n2364_n3288# 1.32574f
C424 source.n173 a_n2364_n3288# 0.014121f
C425 source.n174 a_n2364_n3288# 0.014952f
C426 source.n175 a_n2364_n3288# 0.033378f
C427 source.n176 a_n2364_n3288# 0.033378f
C428 source.n177 a_n2364_n3288# 0.014952f
C429 source.n178 a_n2364_n3288# 0.014121f
C430 source.n179 a_n2364_n3288# 0.026279f
C431 source.n180 a_n2364_n3288# 0.026279f
C432 source.n181 a_n2364_n3288# 0.014121f
C433 source.n182 a_n2364_n3288# 0.014952f
C434 source.n183 a_n2364_n3288# 0.033378f
C435 source.n184 a_n2364_n3288# 0.033378f
C436 source.n185 a_n2364_n3288# 0.014952f
C437 source.n186 a_n2364_n3288# 0.014121f
C438 source.n187 a_n2364_n3288# 0.026279f
C439 source.n188 a_n2364_n3288# 0.026279f
C440 source.n189 a_n2364_n3288# 0.014121f
C441 source.n190 a_n2364_n3288# 0.014121f
C442 source.n191 a_n2364_n3288# 0.014952f
C443 source.n192 a_n2364_n3288# 0.033378f
C444 source.n193 a_n2364_n3288# 0.033378f
C445 source.n194 a_n2364_n3288# 0.033378f
C446 source.n195 a_n2364_n3288# 0.014537f
C447 source.n196 a_n2364_n3288# 0.014121f
C448 source.n197 a_n2364_n3288# 0.026279f
C449 source.n198 a_n2364_n3288# 0.026279f
C450 source.n199 a_n2364_n3288# 0.014121f
C451 source.n200 a_n2364_n3288# 0.014952f
C452 source.n201 a_n2364_n3288# 0.033378f
C453 source.n202 a_n2364_n3288# 0.033378f
C454 source.n203 a_n2364_n3288# 0.014952f
C455 source.n204 a_n2364_n3288# 0.014121f
C456 source.n205 a_n2364_n3288# 0.026279f
C457 source.n206 a_n2364_n3288# 0.026279f
C458 source.n207 a_n2364_n3288# 0.014121f
C459 source.n208 a_n2364_n3288# 0.014952f
C460 source.n209 a_n2364_n3288# 0.033378f
C461 source.n210 a_n2364_n3288# 0.068495f
C462 source.n211 a_n2364_n3288# 0.014952f
C463 source.n212 a_n2364_n3288# 0.014121f
C464 source.n213 a_n2364_n3288# 0.056435f
C465 source.n214 a_n2364_n3288# 0.037802f
C466 source.n215 a_n2364_n3288# 0.172583f
C467 source.t0 a_n2364_n3288# 0.2492f
C468 source.t2 a_n2364_n3288# 0.2492f
C469 source.n216 a_n2364_n3288# 2.13364f
C470 source.n217 a_n2364_n3288# 0.421251f
C471 source.t7 a_n2364_n3288# 0.2492f
C472 source.t9 a_n2364_n3288# 0.2492f
C473 source.n218 a_n2364_n3288# 2.13364f
C474 source.n219 a_n2364_n3288# 0.419061f
C475 source.t10 a_n2364_n3288# 0.2492f
C476 source.t12 a_n2364_n3288# 0.2492f
C477 source.n220 a_n2364_n3288# 2.13364f
C478 source.n221 a_n2364_n3288# 0.419061f
C479 source.n222 a_n2364_n3288# 0.03481f
C480 source.n223 a_n2364_n3288# 0.026279f
C481 source.n224 a_n2364_n3288# 0.014121f
C482 source.n225 a_n2364_n3288# 0.033378f
C483 source.n226 a_n2364_n3288# 0.014952f
C484 source.n227 a_n2364_n3288# 0.026279f
C485 source.n228 a_n2364_n3288# 0.014121f
C486 source.n229 a_n2364_n3288# 0.033378f
C487 source.n230 a_n2364_n3288# 0.014952f
C488 source.n231 a_n2364_n3288# 0.026279f
C489 source.n232 a_n2364_n3288# 0.014537f
C490 source.n233 a_n2364_n3288# 0.033378f
C491 source.n234 a_n2364_n3288# 0.014952f
C492 source.n235 a_n2364_n3288# 0.026279f
C493 source.n236 a_n2364_n3288# 0.014121f
C494 source.n237 a_n2364_n3288# 0.033378f
C495 source.n238 a_n2364_n3288# 0.014952f
C496 source.n239 a_n2364_n3288# 0.026279f
C497 source.n240 a_n2364_n3288# 0.014121f
C498 source.n241 a_n2364_n3288# 0.025033f
C499 source.n242 a_n2364_n3288# 0.023596f
C500 source.t5 a_n2364_n3288# 0.056373f
C501 source.n243 a_n2364_n3288# 0.18947f
C502 source.n244 a_n2364_n3288# 1.32574f
C503 source.n245 a_n2364_n3288# 0.014121f
C504 source.n246 a_n2364_n3288# 0.014952f
C505 source.n247 a_n2364_n3288# 0.033378f
C506 source.n248 a_n2364_n3288# 0.033378f
C507 source.n249 a_n2364_n3288# 0.014952f
C508 source.n250 a_n2364_n3288# 0.014121f
C509 source.n251 a_n2364_n3288# 0.026279f
C510 source.n252 a_n2364_n3288# 0.026279f
C511 source.n253 a_n2364_n3288# 0.014121f
C512 source.n254 a_n2364_n3288# 0.014952f
C513 source.n255 a_n2364_n3288# 0.033378f
C514 source.n256 a_n2364_n3288# 0.033378f
C515 source.n257 a_n2364_n3288# 0.014952f
C516 source.n258 a_n2364_n3288# 0.014121f
C517 source.n259 a_n2364_n3288# 0.026279f
C518 source.n260 a_n2364_n3288# 0.026279f
C519 source.n261 a_n2364_n3288# 0.014121f
C520 source.n262 a_n2364_n3288# 0.014121f
C521 source.n263 a_n2364_n3288# 0.014952f
C522 source.n264 a_n2364_n3288# 0.033378f
C523 source.n265 a_n2364_n3288# 0.033378f
C524 source.n266 a_n2364_n3288# 0.033378f
C525 source.n267 a_n2364_n3288# 0.014537f
C526 source.n268 a_n2364_n3288# 0.014121f
C527 source.n269 a_n2364_n3288# 0.026279f
C528 source.n270 a_n2364_n3288# 0.026279f
C529 source.n271 a_n2364_n3288# 0.014121f
C530 source.n272 a_n2364_n3288# 0.014952f
C531 source.n273 a_n2364_n3288# 0.033378f
C532 source.n274 a_n2364_n3288# 0.033378f
C533 source.n275 a_n2364_n3288# 0.014952f
C534 source.n276 a_n2364_n3288# 0.014121f
C535 source.n277 a_n2364_n3288# 0.026279f
C536 source.n278 a_n2364_n3288# 0.026279f
C537 source.n279 a_n2364_n3288# 0.014121f
C538 source.n280 a_n2364_n3288# 0.014952f
C539 source.n281 a_n2364_n3288# 0.033378f
C540 source.n282 a_n2364_n3288# 0.068495f
C541 source.n283 a_n2364_n3288# 0.014952f
C542 source.n284 a_n2364_n3288# 0.014121f
C543 source.n285 a_n2364_n3288# 0.056435f
C544 source.n286 a_n2364_n3288# 0.037802f
C545 source.n287 a_n2364_n3288# 0.30641f
C546 source.n288 a_n2364_n3288# 1.66526f
C547 drain_left.n0 a_n2364_n3288# 0.033166f
C548 drain_left.n1 a_n2364_n3288# 0.025038f
C549 drain_left.n2 a_n2364_n3288# 0.013454f
C550 drain_left.n3 a_n2364_n3288# 0.031801f
C551 drain_left.n4 a_n2364_n3288# 0.014246f
C552 drain_left.n5 a_n2364_n3288# 0.025038f
C553 drain_left.n6 a_n2364_n3288# 0.013454f
C554 drain_left.n7 a_n2364_n3288# 0.031801f
C555 drain_left.n8 a_n2364_n3288# 0.014246f
C556 drain_left.n9 a_n2364_n3288# 0.025038f
C557 drain_left.n10 a_n2364_n3288# 0.01385f
C558 drain_left.n11 a_n2364_n3288# 0.031801f
C559 drain_left.n12 a_n2364_n3288# 0.014246f
C560 drain_left.n13 a_n2364_n3288# 0.025038f
C561 drain_left.n14 a_n2364_n3288# 0.013454f
C562 drain_left.n15 a_n2364_n3288# 0.031801f
C563 drain_left.n16 a_n2364_n3288# 0.014246f
C564 drain_left.n17 a_n2364_n3288# 0.025038f
C565 drain_left.n18 a_n2364_n3288# 0.013454f
C566 drain_left.n19 a_n2364_n3288# 0.023851f
C567 drain_left.n20 a_n2364_n3288# 0.022481f
C568 drain_left.t1 a_n2364_n3288# 0.05371f
C569 drain_left.n21 a_n2364_n3288# 0.18052f
C570 drain_left.n22 a_n2364_n3288# 1.26312f
C571 drain_left.n23 a_n2364_n3288# 0.013454f
C572 drain_left.n24 a_n2364_n3288# 0.014246f
C573 drain_left.n25 a_n2364_n3288# 0.031801f
C574 drain_left.n26 a_n2364_n3288# 0.031801f
C575 drain_left.n27 a_n2364_n3288# 0.014246f
C576 drain_left.n28 a_n2364_n3288# 0.013454f
C577 drain_left.n29 a_n2364_n3288# 0.025038f
C578 drain_left.n30 a_n2364_n3288# 0.025038f
C579 drain_left.n31 a_n2364_n3288# 0.013454f
C580 drain_left.n32 a_n2364_n3288# 0.014246f
C581 drain_left.n33 a_n2364_n3288# 0.031801f
C582 drain_left.n34 a_n2364_n3288# 0.031801f
C583 drain_left.n35 a_n2364_n3288# 0.014246f
C584 drain_left.n36 a_n2364_n3288# 0.013454f
C585 drain_left.n37 a_n2364_n3288# 0.025038f
C586 drain_left.n38 a_n2364_n3288# 0.025038f
C587 drain_left.n39 a_n2364_n3288# 0.013454f
C588 drain_left.n40 a_n2364_n3288# 0.013454f
C589 drain_left.n41 a_n2364_n3288# 0.014246f
C590 drain_left.n42 a_n2364_n3288# 0.031801f
C591 drain_left.n43 a_n2364_n3288# 0.031801f
C592 drain_left.n44 a_n2364_n3288# 0.031801f
C593 drain_left.n45 a_n2364_n3288# 0.01385f
C594 drain_left.n46 a_n2364_n3288# 0.013454f
C595 drain_left.n47 a_n2364_n3288# 0.025038f
C596 drain_left.n48 a_n2364_n3288# 0.025038f
C597 drain_left.n49 a_n2364_n3288# 0.013454f
C598 drain_left.n50 a_n2364_n3288# 0.014246f
C599 drain_left.n51 a_n2364_n3288# 0.031801f
C600 drain_left.n52 a_n2364_n3288# 0.031801f
C601 drain_left.n53 a_n2364_n3288# 0.014246f
C602 drain_left.n54 a_n2364_n3288# 0.013454f
C603 drain_left.n55 a_n2364_n3288# 0.025038f
C604 drain_left.n56 a_n2364_n3288# 0.025038f
C605 drain_left.n57 a_n2364_n3288# 0.013454f
C606 drain_left.n58 a_n2364_n3288# 0.014246f
C607 drain_left.n59 a_n2364_n3288# 0.031801f
C608 drain_left.n60 a_n2364_n3288# 0.065259f
C609 drain_left.n61 a_n2364_n3288# 0.014246f
C610 drain_left.n62 a_n2364_n3288# 0.013454f
C611 drain_left.n63 a_n2364_n3288# 0.053769f
C612 drain_left.n64 a_n2364_n3288# 0.05554f
C613 drain_left.t2 a_n2364_n3288# 0.237428f
C614 drain_left.t11 a_n2364_n3288# 0.237428f
C615 drain_left.n65 a_n2364_n3288# 2.11274f
C616 drain_left.n66 a_n2364_n3288# 0.447281f
C617 drain_left.t4 a_n2364_n3288# 0.237428f
C618 drain_left.t3 a_n2364_n3288# 0.237428f
C619 drain_left.n67 a_n2364_n3288# 2.11808f
C620 drain_left.t12 a_n2364_n3288# 0.237428f
C621 drain_left.t8 a_n2364_n3288# 0.237428f
C622 drain_left.n68 a_n2364_n3288# 2.11274f
C623 drain_left.n69 a_n2364_n3288# 0.656844f
C624 drain_left.n70 a_n2364_n3288# 1.38279f
C625 drain_left.n71 a_n2364_n3288# 0.033166f
C626 drain_left.n72 a_n2364_n3288# 0.025038f
C627 drain_left.n73 a_n2364_n3288# 0.013454f
C628 drain_left.n74 a_n2364_n3288# 0.031801f
C629 drain_left.n75 a_n2364_n3288# 0.014246f
C630 drain_left.n76 a_n2364_n3288# 0.025038f
C631 drain_left.n77 a_n2364_n3288# 0.013454f
C632 drain_left.n78 a_n2364_n3288# 0.031801f
C633 drain_left.n79 a_n2364_n3288# 0.014246f
C634 drain_left.n80 a_n2364_n3288# 0.025038f
C635 drain_left.n81 a_n2364_n3288# 0.01385f
C636 drain_left.n82 a_n2364_n3288# 0.031801f
C637 drain_left.n83 a_n2364_n3288# 0.013454f
C638 drain_left.n84 a_n2364_n3288# 0.014246f
C639 drain_left.n85 a_n2364_n3288# 0.025038f
C640 drain_left.n86 a_n2364_n3288# 0.013454f
C641 drain_left.n87 a_n2364_n3288# 0.031801f
C642 drain_left.n88 a_n2364_n3288# 0.014246f
C643 drain_left.n89 a_n2364_n3288# 0.025038f
C644 drain_left.n90 a_n2364_n3288# 0.013454f
C645 drain_left.n91 a_n2364_n3288# 0.023851f
C646 drain_left.n92 a_n2364_n3288# 0.022481f
C647 drain_left.t5 a_n2364_n3288# 0.05371f
C648 drain_left.n93 a_n2364_n3288# 0.18052f
C649 drain_left.n94 a_n2364_n3288# 1.26312f
C650 drain_left.n95 a_n2364_n3288# 0.013454f
C651 drain_left.n96 a_n2364_n3288# 0.014246f
C652 drain_left.n97 a_n2364_n3288# 0.031801f
C653 drain_left.n98 a_n2364_n3288# 0.031801f
C654 drain_left.n99 a_n2364_n3288# 0.014246f
C655 drain_left.n100 a_n2364_n3288# 0.013454f
C656 drain_left.n101 a_n2364_n3288# 0.025038f
C657 drain_left.n102 a_n2364_n3288# 0.025038f
C658 drain_left.n103 a_n2364_n3288# 0.013454f
C659 drain_left.n104 a_n2364_n3288# 0.014246f
C660 drain_left.n105 a_n2364_n3288# 0.031801f
C661 drain_left.n106 a_n2364_n3288# 0.031801f
C662 drain_left.n107 a_n2364_n3288# 0.014246f
C663 drain_left.n108 a_n2364_n3288# 0.013454f
C664 drain_left.n109 a_n2364_n3288# 0.025038f
C665 drain_left.n110 a_n2364_n3288# 0.025038f
C666 drain_left.n111 a_n2364_n3288# 0.013454f
C667 drain_left.n112 a_n2364_n3288# 0.014246f
C668 drain_left.n113 a_n2364_n3288# 0.031801f
C669 drain_left.n114 a_n2364_n3288# 0.031801f
C670 drain_left.n115 a_n2364_n3288# 0.031801f
C671 drain_left.n116 a_n2364_n3288# 0.01385f
C672 drain_left.n117 a_n2364_n3288# 0.013454f
C673 drain_left.n118 a_n2364_n3288# 0.025038f
C674 drain_left.n119 a_n2364_n3288# 0.025038f
C675 drain_left.n120 a_n2364_n3288# 0.013454f
C676 drain_left.n121 a_n2364_n3288# 0.014246f
C677 drain_left.n122 a_n2364_n3288# 0.031801f
C678 drain_left.n123 a_n2364_n3288# 0.031801f
C679 drain_left.n124 a_n2364_n3288# 0.014246f
C680 drain_left.n125 a_n2364_n3288# 0.013454f
C681 drain_left.n126 a_n2364_n3288# 0.025038f
C682 drain_left.n127 a_n2364_n3288# 0.025038f
C683 drain_left.n128 a_n2364_n3288# 0.013454f
C684 drain_left.n129 a_n2364_n3288# 0.014246f
C685 drain_left.n130 a_n2364_n3288# 0.031801f
C686 drain_left.n131 a_n2364_n3288# 0.065259f
C687 drain_left.n132 a_n2364_n3288# 0.014246f
C688 drain_left.n133 a_n2364_n3288# 0.013454f
C689 drain_left.n134 a_n2364_n3288# 0.053769f
C690 drain_left.n135 a_n2364_n3288# 0.05554f
C691 drain_left.t7 a_n2364_n3288# 0.237428f
C692 drain_left.t9 a_n2364_n3288# 0.237428f
C693 drain_left.n136 a_n2364_n3288# 2.11275f
C694 drain_left.n137 a_n2364_n3288# 0.468696f
C695 drain_left.t10 a_n2364_n3288# 0.237428f
C696 drain_left.t6 a_n2364_n3288# 0.237428f
C697 drain_left.n138 a_n2364_n3288# 2.11275f
C698 drain_left.n139 a_n2364_n3288# 0.353395f
C699 drain_left.t13 a_n2364_n3288# 0.237428f
C700 drain_left.t0 a_n2364_n3288# 0.237428f
C701 drain_left.n140 a_n2364_n3288# 2.11274f
C702 drain_left.n141 a_n2364_n3288# 0.574865f
C703 plus.n0 a_n2364_n3288# 0.041591f
C704 plus.t2 a_n2364_n3288# 0.996214f
C705 plus.t9 a_n2364_n3288# 0.996214f
C706 plus.n1 a_n2364_n3288# 0.041591f
C707 plus.t4 a_n2364_n3288# 0.996214f
C708 plus.n2 a_n2364_n3288# 0.397309f
C709 plus.n3 a_n2364_n3288# 0.041591f
C710 plus.t8 a_n2364_n3288# 0.996214f
C711 plus.t3 a_n2364_n3288# 0.996214f
C712 plus.n4 a_n2364_n3288# 0.397309f
C713 plus.t5 a_n2364_n3288# 1.01543f
C714 plus.n5 a_n2364_n3288# 0.381708f
C715 plus.t10 a_n2364_n3288# 0.996214f
C716 plus.n6 a_n2364_n3288# 0.402461f
C717 plus.n7 a_n2364_n3288# 0.009438f
C718 plus.n8 a_n2364_n3288# 0.175241f
C719 plus.n9 a_n2364_n3288# 0.041591f
C720 plus.n10 a_n2364_n3288# 0.041591f
C721 plus.n11 a_n2364_n3288# 0.009438f
C722 plus.n12 a_n2364_n3288# 0.397309f
C723 plus.n13 a_n2364_n3288# 0.009438f
C724 plus.n14 a_n2364_n3288# 0.041591f
C725 plus.n15 a_n2364_n3288# 0.041591f
C726 plus.n16 a_n2364_n3288# 0.041591f
C727 plus.n17 a_n2364_n3288# 0.009438f
C728 plus.n18 a_n2364_n3288# 0.397309f
C729 plus.n19 a_n2364_n3288# 0.009438f
C730 plus.n20 a_n2364_n3288# 0.39577f
C731 plus.n21 a_n2364_n3288# 0.480209f
C732 plus.n22 a_n2364_n3288# 0.041591f
C733 plus.t1 a_n2364_n3288# 0.996214f
C734 plus.n23 a_n2364_n3288# 0.041591f
C735 plus.t0 a_n2364_n3288# 0.996214f
C736 plus.t7 a_n2364_n3288# 0.996214f
C737 plus.n24 a_n2364_n3288# 0.397309f
C738 plus.n25 a_n2364_n3288# 0.041591f
C739 plus.t6 a_n2364_n3288# 0.996214f
C740 plus.t11 a_n2364_n3288# 0.996214f
C741 plus.n26 a_n2364_n3288# 0.397309f
C742 plus.t12 a_n2364_n3288# 1.01543f
C743 plus.n27 a_n2364_n3288# 0.381708f
C744 plus.t13 a_n2364_n3288# 0.996214f
C745 plus.n28 a_n2364_n3288# 0.402461f
C746 plus.n29 a_n2364_n3288# 0.009438f
C747 plus.n30 a_n2364_n3288# 0.175241f
C748 plus.n31 a_n2364_n3288# 0.041591f
C749 plus.n32 a_n2364_n3288# 0.041591f
C750 plus.n33 a_n2364_n3288# 0.009438f
C751 plus.n34 a_n2364_n3288# 0.397309f
C752 plus.n35 a_n2364_n3288# 0.009438f
C753 plus.n36 a_n2364_n3288# 0.041591f
C754 plus.n37 a_n2364_n3288# 0.041591f
C755 plus.n38 a_n2364_n3288# 0.041591f
C756 plus.n39 a_n2364_n3288# 0.009438f
C757 plus.n40 a_n2364_n3288# 0.397309f
C758 plus.n41 a_n2364_n3288# 0.009438f
C759 plus.n42 a_n2364_n3288# 0.39577f
C760 plus.n43 a_n2364_n3288# 1.36461f
.ends

