* NGSPICE file created from diffpair621.ext - technology: sky130A

.subckt diffpair621 minus drain_right drain_left source plus
X0 drain_left.t3 plus.t0 source.t7 a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X1 source.t5 plus.t1 drain_left.t2 a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X2 a_n1334_n4888# a_n1334_n4888# a_n1334_n4888# a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.7
X3 source.t3 minus.t0 drain_right.t3 a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X4 source.t4 plus.t2 drain_left.t1 a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X5 drain_right.t2 minus.t1 source.t2 a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X6 source.t1 minus.t2 drain_right.t1 a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X7 a_n1334_n4888# a_n1334_n4888# a_n1334_n4888# a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X8 drain_right.t0 minus.t3 source.t0 a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X9 drain_left.t0 plus.t3 source.t6 a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X10 a_n1334_n4888# a_n1334_n4888# a_n1334_n4888# a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X11 a_n1334_n4888# a_n1334_n4888# a_n1334_n4888# a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
R0 plus.n0 plus.t2 765.687
R1 plus.n1 plus.t0 765.687
R2 plus.n0 plus.t3 765.638
R3 plus.n1 plus.t1 765.638
R4 plus plus.n1 75.8689
R5 plus plus.n0 59.9575
R6 source.n0 source.t6 44.1297
R7 source.n1 source.t4 44.1296
R8 source.n2 source.t0 44.1296
R9 source.n3 source.t3 44.1296
R10 source.n7 source.t2 44.1295
R11 source.n6 source.t1 44.1295
R12 source.n5 source.t7 44.1295
R13 source.n4 source.t5 44.1295
R14 source.n4 source.n3 28.2363
R15 source.n8 source.n0 22.5294
R16 source.n8 source.n7 5.7074
R17 source.n3 source.n2 0.888431
R18 source.n1 source.n0 0.888431
R19 source.n5 source.n4 0.888431
R20 source.n7 source.n6 0.888431
R21 source.n2 source.n1 0.470328
R22 source.n6 source.n5 0.470328
R23 source source.n8 0.188
R24 drain_left drain_left.n0 95.0214
R25 drain_left drain_left.n1 66.3591
R26 drain_left.n0 drain_left.t2 0.9905
R27 drain_left.n0 drain_left.t3 0.9905
R28 drain_left.n1 drain_left.t1 0.9905
R29 drain_left.n1 drain_left.t0 0.9905
R30 minus.n0 minus.t3 765.687
R31 minus.n1 minus.t2 765.687
R32 minus.n0 minus.t0 765.638
R33 minus.n1 minus.t1 765.638
R34 minus.n2 minus.n0 85.0181
R35 minus.n2 minus.n1 51.2833
R36 minus minus.n2 0.188
R37 drain_right drain_right.n0 94.4682
R38 drain_right drain_right.n1 66.3591
R39 drain_right.n0 drain_right.t1 0.9905
R40 drain_right.n0 drain_right.t2 0.9905
R41 drain_right.n1 drain_right.t3 0.9905
R42 drain_right.n1 drain_right.t0 0.9905
C0 minus drain_right 5.10577f
C1 source minus 4.37327f
C2 plus drain_left 5.23172f
C3 plus drain_right 0.279168f
C4 plus source 4.38731f
C5 plus minus 6.28551f
C6 drain_left drain_right 0.565372f
C7 drain_left source 10.5531f
C8 drain_left minus 0.170337f
C9 source drain_right 10.5541f
C10 drain_right a_n1334_n4888# 8.40371f
C11 drain_left a_n1334_n4888# 8.61276f
C12 source a_n1334_n4888# 13.370366f
C13 minus a_n1334_n4888# 5.555969f
C14 plus a_n1334_n4888# 9.50793f
C15 drain_right.t1 a_n1334_n4888# 0.441831f
C16 drain_right.t2 a_n1334_n4888# 0.441831f
C17 drain_right.n0 a_n1334_n4888# 4.68882f
C18 drain_right.t3 a_n1334_n4888# 0.441831f
C19 drain_right.t0 a_n1334_n4888# 0.441831f
C20 drain_right.n1 a_n1334_n4888# 4.10381f
C21 minus.t3 a_n1334_n4888# 1.96809f
C22 minus.t0 a_n1334_n4888# 1.96804f
C23 minus.n0 a_n1334_n4888# 2.44181f
C24 minus.t2 a_n1334_n4888# 1.96809f
C25 minus.t1 a_n1334_n4888# 1.96804f
C26 minus.n1 a_n1334_n4888# 1.4733f
C27 minus.n2 a_n1334_n4888# 3.98037f
C28 drain_left.t2 a_n1334_n4888# 0.44157f
C29 drain_left.t3 a_n1334_n4888# 0.44157f
C30 drain_left.n0 a_n1334_n4888# 4.7143f
C31 drain_left.t1 a_n1334_n4888# 0.44157f
C32 drain_left.t0 a_n1334_n4888# 0.44157f
C33 drain_left.n1 a_n1334_n4888# 4.10139f
C34 source.t6 a_n1334_n4888# 2.83975f
C35 source.n0 a_n1334_n4888# 1.23537f
C36 source.t4 a_n1334_n4888# 2.83975f
C37 source.n1 a_n1334_n4888# 0.28969f
C38 source.t0 a_n1334_n4888# 2.83975f
C39 source.n2 a_n1334_n4888# 0.28969f
C40 source.t3 a_n1334_n4888# 2.83975f
C41 source.n3 a_n1334_n4888# 1.52139f
C42 source.t5 a_n1334_n4888# 2.83974f
C43 source.n4 a_n1334_n4888# 1.52141f
C44 source.t7 a_n1334_n4888# 2.83974f
C45 source.n5 a_n1334_n4888# 0.289705f
C46 source.t1 a_n1334_n4888# 2.83974f
C47 source.n6 a_n1334_n4888# 0.289705f
C48 source.t2 a_n1334_n4888# 2.83974f
C49 source.n7 a_n1334_n4888# 0.392261f
C50 source.n8 a_n1334_n4888# 1.42636f
C51 plus.t3 a_n1334_n4888# 1.99303f
C52 plus.t2 a_n1334_n4888# 1.99308f
C53 plus.n0 a_n1334_n4888# 1.65787f
C54 plus.t0 a_n1334_n4888# 1.99308f
C55 plus.t1 a_n1334_n4888# 1.99303f
C56 plus.n1 a_n1334_n4888# 2.15158f
.ends

