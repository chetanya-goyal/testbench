* NGSPICE file created from diffpair139.ext - technology: sky130A

.subckt diffpair139 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t22 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X1 a_n3134_n1288# a_n3134_n1288# a_n3134_n1288# a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.6
X2 a_n3134_n1288# a_n3134_n1288# a_n3134_n1288# a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X3 drain_right.t23 minus.t0 source.t9 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X4 drain_left.t22 plus.t1 source.t36 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X5 source.t24 plus.t2 drain_left.t21 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X6 drain_left.t20 plus.t3 source.t23 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X7 source.t1 minus.t1 drain_right.t22 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X8 source.t33 plus.t4 drain_left.t19 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X9 drain_right.t21 minus.t2 source.t5 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X10 source.t12 minus.t3 drain_right.t20 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X11 a_n3134_n1288# a_n3134_n1288# a_n3134_n1288# a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X12 drain_left.t18 plus.t5 source.t37 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X13 source.t15 minus.t4 drain_right.t19 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X14 source.t35 plus.t6 drain_left.t17 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X15 source.t16 minus.t5 drain_right.t18 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X16 source.t10 minus.t6 drain_right.t17 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X17 drain_right.t16 minus.t7 source.t46 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X18 drain_right.t15 minus.t8 source.t47 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X19 drain_right.t14 minus.t9 source.t3 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X20 drain_right.t13 minus.t10 source.t0 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X21 source.t2 minus.t11 drain_right.t12 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X22 source.t28 plus.t7 drain_left.t16 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X23 source.t19 minus.t12 drain_right.t11 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X24 drain_left.t15 plus.t8 source.t42 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X25 drain_left.t14 plus.t9 source.t29 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X26 source.t43 plus.t10 drain_left.t13 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X27 source.t44 plus.t11 drain_left.t12 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X28 source.t11 minus.t13 drain_right.t10 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X29 source.t7 minus.t14 drain_right.t9 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X30 drain_right.t8 minus.t15 source.t13 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X31 drain_left.t11 plus.t12 source.t39 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X32 source.t17 minus.t16 drain_right.t7 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X33 source.t40 plus.t13 drain_left.t10 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X34 drain_right.t6 minus.t17 source.t6 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X35 drain_right.t5 minus.t18 source.t8 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X36 source.t21 minus.t19 drain_right.t4 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X37 source.t27 plus.t14 drain_left.t9 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X38 source.t26 plus.t15 drain_left.t8 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X39 drain_left.t7 plus.t16 source.t45 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X40 drain_left.t6 plus.t17 source.t38 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X41 source.t41 plus.t18 drain_left.t5 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X42 source.t31 plus.t19 drain_left.t4 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X43 drain_right.t3 minus.t20 source.t20 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X44 drain_right.t2 minus.t21 source.t18 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X45 source.t14 minus.t22 drain_right.t1 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X46 source.t34 plus.t20 drain_left.t3 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X47 drain_right.t0 minus.t23 source.t4 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X48 drain_left.t2 plus.t21 source.t32 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
X49 a_n3134_n1288# a_n3134_n1288# a_n3134_n1288# a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X50 drain_left.t1 plus.t22 source.t25 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X51 drain_left.t0 plus.t23 source.t30 a_n3134_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.6
R0 plus.n9 plus.t18 172.163
R1 plus.n43 plus.t22 172.163
R2 plus.n13 plus.n8 161.3
R3 plus.n15 plus.n14 161.3
R4 plus.n16 plus.n7 161.3
R5 plus.n18 plus.n17 161.3
R6 plus.n19 plus.n6 161.3
R7 plus.n21 plus.n20 161.3
R8 plus.n22 plus.n5 161.3
R9 plus.n24 plus.n23 161.3
R10 plus.n25 plus.n4 161.3
R11 plus.n27 plus.n26 161.3
R12 plus.n28 plus.n3 161.3
R13 plus.n30 plus.n1 161.3
R14 plus.n31 plus.n0 161.3
R15 plus.n33 plus.n32 161.3
R16 plus.n47 plus.n42 161.3
R17 plus.n49 plus.n48 161.3
R18 plus.n50 plus.n41 161.3
R19 plus.n52 plus.n51 161.3
R20 plus.n53 plus.n40 161.3
R21 plus.n55 plus.n54 161.3
R22 plus.n56 plus.n39 161.3
R23 plus.n58 plus.n57 161.3
R24 plus.n59 plus.n38 161.3
R25 plus.n61 plus.n60 161.3
R26 plus.n62 plus.n37 161.3
R27 plus.n64 plus.n35 161.3
R28 plus.n65 plus.n34 161.3
R29 plus.n67 plus.n66 161.3
R30 plus.n32 plus.t16 145.805
R31 plus.n30 plus.t19 145.805
R32 plus.n29 plus.t0 145.805
R33 plus.n28 plus.t2 145.805
R34 plus.n4 plus.t3 145.805
R35 plus.n22 plus.t4 145.805
R36 plus.n6 plus.t5 145.805
R37 plus.n16 plus.t10 145.805
R38 plus.n8 plus.t12 145.805
R39 plus.n11 plus.t13 145.805
R40 plus.n10 plus.t17 145.805
R41 plus.n66 plus.t15 145.805
R42 plus.n64 plus.t21 145.805
R43 plus.n63 plus.t14 145.805
R44 plus.n62 plus.t1 145.805
R45 plus.n38 plus.t7 145.805
R46 plus.n56 plus.t9 145.805
R47 plus.n40 plus.t20 145.805
R48 plus.n50 plus.t23 145.805
R49 plus.n42 plus.t6 145.805
R50 plus.n45 plus.t8 145.805
R51 plus.n44 plus.t11 145.805
R52 plus.n12 plus.n11 80.6037
R53 plus.n29 plus.n2 80.6037
R54 plus.n46 plus.n45 80.6037
R55 plus.n63 plus.n36 80.6037
R56 plus.n30 plus.n29 48.2005
R57 plus.n29 plus.n28 48.2005
R58 plus.n11 plus.n8 48.2005
R59 plus.n11 plus.n10 48.2005
R60 plus.n64 plus.n63 48.2005
R61 plus.n63 plus.n62 48.2005
R62 plus.n45 plus.n42 48.2005
R63 plus.n45 plus.n44 48.2005
R64 plus.n32 plus.n31 46.0096
R65 plus.n66 plus.n65 46.0096
R66 plus.n12 plus.n9 45.1822
R67 plus.n46 plus.n43 45.1822
R68 plus.n27 plus.n4 44.549
R69 plus.n16 plus.n15 44.549
R70 plus.n61 plus.n38 44.549
R71 plus.n50 plus.n49 44.549
R72 plus.n23 plus.n22 34.3247
R73 plus.n17 plus.n6 34.3247
R74 plus.n57 plus.n56 34.3247
R75 plus.n51 plus.n40 34.3247
R76 plus plus.n67 31.1884
R77 plus.n21 plus.n6 24.1005
R78 plus.n22 plus.n21 24.1005
R79 plus.n56 plus.n55 24.1005
R80 plus.n55 plus.n40 24.1005
R81 plus.n10 plus.n9 14.1472
R82 plus.n44 plus.n43 14.1472
R83 plus.n23 plus.n4 13.8763
R84 plus.n17 plus.n16 13.8763
R85 plus.n57 plus.n38 13.8763
R86 plus.n51 plus.n50 13.8763
R87 plus plus.n33 8.45883
R88 plus.n28 plus.n27 3.65202
R89 plus.n15 plus.n8 3.65202
R90 plus.n62 plus.n61 3.65202
R91 plus.n49 plus.n42 3.65202
R92 plus.n31 plus.n30 2.19141
R93 plus.n65 plus.n64 2.19141
R94 plus.n13 plus.n12 0.285035
R95 plus.n3 plus.n2 0.285035
R96 plus.n2 plus.n1 0.285035
R97 plus.n36 plus.n35 0.285035
R98 plus.n37 plus.n36 0.285035
R99 plus.n47 plus.n46 0.285035
R100 plus.n14 plus.n13 0.189894
R101 plus.n14 plus.n7 0.189894
R102 plus.n18 plus.n7 0.189894
R103 plus.n19 plus.n18 0.189894
R104 plus.n20 plus.n19 0.189894
R105 plus.n20 plus.n5 0.189894
R106 plus.n24 plus.n5 0.189894
R107 plus.n25 plus.n24 0.189894
R108 plus.n26 plus.n25 0.189894
R109 plus.n26 plus.n3 0.189894
R110 plus.n1 plus.n0 0.189894
R111 plus.n33 plus.n0 0.189894
R112 plus.n67 plus.n34 0.189894
R113 plus.n35 plus.n34 0.189894
R114 plus.n60 plus.n37 0.189894
R115 plus.n60 plus.n59 0.189894
R116 plus.n59 plus.n58 0.189894
R117 plus.n58 plus.n39 0.189894
R118 plus.n54 plus.n39 0.189894
R119 plus.n54 plus.n53 0.189894
R120 plus.n53 plus.n52 0.189894
R121 plus.n52 plus.n41 0.189894
R122 plus.n48 plus.n41 0.189894
R123 plus.n48 plus.n47 0.189894
R124 source.n98 source.n96 289.615
R125 source.n80 source.n78 289.615
R126 source.n72 source.n70 289.615
R127 source.n54 source.n52 289.615
R128 source.n2 source.n0 289.615
R129 source.n20 source.n18 289.615
R130 source.n28 source.n26 289.615
R131 source.n46 source.n44 289.615
R132 source.n99 source.n98 185
R133 source.n81 source.n80 185
R134 source.n73 source.n72 185
R135 source.n55 source.n54 185
R136 source.n3 source.n2 185
R137 source.n21 source.n20 185
R138 source.n29 source.n28 185
R139 source.n47 source.n46 185
R140 source.t18 source.n97 167.117
R141 source.t2 source.n79 167.117
R142 source.t25 source.n71 167.117
R143 source.t26 source.n53 167.117
R144 source.t45 source.n1 167.117
R145 source.t41 source.n19 167.117
R146 source.t6 source.n27 167.117
R147 source.t7 source.n45 167.117
R148 source.n9 source.n8 84.1169
R149 source.n11 source.n10 84.1169
R150 source.n13 source.n12 84.1169
R151 source.n15 source.n14 84.1169
R152 source.n17 source.n16 84.1169
R153 source.n35 source.n34 84.1169
R154 source.n37 source.n36 84.1169
R155 source.n39 source.n38 84.1169
R156 source.n41 source.n40 84.1169
R157 source.n43 source.n42 84.1169
R158 source.n95 source.n94 84.1168
R159 source.n93 source.n92 84.1168
R160 source.n91 source.n90 84.1168
R161 source.n89 source.n88 84.1168
R162 source.n87 source.n86 84.1168
R163 source.n69 source.n68 84.1168
R164 source.n67 source.n66 84.1168
R165 source.n65 source.n64 84.1168
R166 source.n63 source.n62 84.1168
R167 source.n61 source.n60 84.1168
R168 source.n98 source.t18 52.3082
R169 source.n80 source.t2 52.3082
R170 source.n72 source.t25 52.3082
R171 source.n54 source.t26 52.3082
R172 source.n2 source.t45 52.3082
R173 source.n20 source.t41 52.3082
R174 source.n28 source.t6 52.3082
R175 source.n46 source.t7 52.3082
R176 source.n103 source.n102 31.4096
R177 source.n85 source.n84 31.4096
R178 source.n77 source.n76 31.4096
R179 source.n59 source.n58 31.4096
R180 source.n7 source.n6 31.4096
R181 source.n25 source.n24 31.4096
R182 source.n33 source.n32 31.4096
R183 source.n51 source.n50 31.4096
R184 source.n59 source.n51 14.5137
R185 source.n94 source.t9 9.9005
R186 source.n94 source.t16 9.9005
R187 source.n92 source.t8 9.9005
R188 source.n92 source.t10 9.9005
R189 source.n90 source.t46 9.9005
R190 source.n90 source.t14 9.9005
R191 source.n88 source.t0 9.9005
R192 source.n88 source.t12 9.9005
R193 source.n86 source.t4 9.9005
R194 source.n86 source.t21 9.9005
R195 source.n68 source.t42 9.9005
R196 source.n68 source.t44 9.9005
R197 source.n66 source.t30 9.9005
R198 source.n66 source.t35 9.9005
R199 source.n64 source.t29 9.9005
R200 source.n64 source.t34 9.9005
R201 source.n62 source.t36 9.9005
R202 source.n62 source.t28 9.9005
R203 source.n60 source.t32 9.9005
R204 source.n60 source.t27 9.9005
R205 source.n8 source.t22 9.9005
R206 source.n8 source.t31 9.9005
R207 source.n10 source.t23 9.9005
R208 source.n10 source.t24 9.9005
R209 source.n12 source.t37 9.9005
R210 source.n12 source.t33 9.9005
R211 source.n14 source.t39 9.9005
R212 source.n14 source.t43 9.9005
R213 source.n16 source.t38 9.9005
R214 source.n16 source.t40 9.9005
R215 source.n34 source.t13 9.9005
R216 source.n34 source.t17 9.9005
R217 source.n36 source.t47 9.9005
R218 source.n36 source.t11 9.9005
R219 source.n38 source.t3 9.9005
R220 source.n38 source.t19 9.9005
R221 source.n40 source.t5 9.9005
R222 source.n40 source.t15 9.9005
R223 source.n42 source.t20 9.9005
R224 source.n42 source.t1 9.9005
R225 source.n99 source.n97 9.71174
R226 source.n81 source.n79 9.71174
R227 source.n73 source.n71 9.71174
R228 source.n55 source.n53 9.71174
R229 source.n3 source.n1 9.71174
R230 source.n21 source.n19 9.71174
R231 source.n29 source.n27 9.71174
R232 source.n47 source.n45 9.71174
R233 source.n102 source.n101 9.45567
R234 source.n84 source.n83 9.45567
R235 source.n76 source.n75 9.45567
R236 source.n58 source.n57 9.45567
R237 source.n6 source.n5 9.45567
R238 source.n24 source.n23 9.45567
R239 source.n32 source.n31 9.45567
R240 source.n50 source.n49 9.45567
R241 source.n101 source.n100 9.3005
R242 source.n83 source.n82 9.3005
R243 source.n75 source.n74 9.3005
R244 source.n57 source.n56 9.3005
R245 source.n5 source.n4 9.3005
R246 source.n23 source.n22 9.3005
R247 source.n31 source.n30 9.3005
R248 source.n49 source.n48 9.3005
R249 source.n104 source.n7 8.8499
R250 source.n102 source.n96 8.14595
R251 source.n84 source.n78 8.14595
R252 source.n76 source.n70 8.14595
R253 source.n58 source.n52 8.14595
R254 source.n6 source.n0 8.14595
R255 source.n24 source.n18 8.14595
R256 source.n32 source.n26 8.14595
R257 source.n50 source.n44 8.14595
R258 source.n100 source.n99 7.3702
R259 source.n82 source.n81 7.3702
R260 source.n74 source.n73 7.3702
R261 source.n56 source.n55 7.3702
R262 source.n4 source.n3 7.3702
R263 source.n22 source.n21 7.3702
R264 source.n30 source.n29 7.3702
R265 source.n48 source.n47 7.3702
R266 source.n100 source.n96 5.81868
R267 source.n82 source.n78 5.81868
R268 source.n74 source.n70 5.81868
R269 source.n56 source.n52 5.81868
R270 source.n4 source.n0 5.81868
R271 source.n22 source.n18 5.81868
R272 source.n30 source.n26 5.81868
R273 source.n48 source.n44 5.81868
R274 source.n104 source.n103 5.66429
R275 source.n101 source.n97 3.44771
R276 source.n83 source.n79 3.44771
R277 source.n75 source.n71 3.44771
R278 source.n57 source.n53 3.44771
R279 source.n5 source.n1 3.44771
R280 source.n23 source.n19 3.44771
R281 source.n31 source.n27 3.44771
R282 source.n49 source.n45 3.44771
R283 source.n51 source.n43 0.802224
R284 source.n43 source.n41 0.802224
R285 source.n41 source.n39 0.802224
R286 source.n39 source.n37 0.802224
R287 source.n37 source.n35 0.802224
R288 source.n35 source.n33 0.802224
R289 source.n25 source.n17 0.802224
R290 source.n17 source.n15 0.802224
R291 source.n15 source.n13 0.802224
R292 source.n13 source.n11 0.802224
R293 source.n11 source.n9 0.802224
R294 source.n9 source.n7 0.802224
R295 source.n61 source.n59 0.802224
R296 source.n63 source.n61 0.802224
R297 source.n65 source.n63 0.802224
R298 source.n67 source.n65 0.802224
R299 source.n69 source.n67 0.802224
R300 source.n77 source.n69 0.802224
R301 source.n87 source.n85 0.802224
R302 source.n89 source.n87 0.802224
R303 source.n91 source.n89 0.802224
R304 source.n93 source.n91 0.802224
R305 source.n95 source.n93 0.802224
R306 source.n103 source.n95 0.802224
R307 source.n33 source.n25 0.470328
R308 source.n85 source.n77 0.470328
R309 source source.n104 0.188
R310 drain_left.n13 drain_left.n11 101.597
R311 drain_left.n7 drain_left.n5 101.597
R312 drain_left.n2 drain_left.n0 101.597
R313 drain_left.n21 drain_left.n20 100.796
R314 drain_left.n19 drain_left.n18 100.796
R315 drain_left.n17 drain_left.n16 100.796
R316 drain_left.n15 drain_left.n14 100.796
R317 drain_left.n13 drain_left.n12 100.796
R318 drain_left.n7 drain_left.n6 100.796
R319 drain_left.n9 drain_left.n8 100.796
R320 drain_left.n4 drain_left.n3 100.796
R321 drain_left.n2 drain_left.n1 100.796
R322 drain_left drain_left.n10 27.4077
R323 drain_left.n5 drain_left.t12 9.9005
R324 drain_left.n5 drain_left.t1 9.9005
R325 drain_left.n6 drain_left.t17 9.9005
R326 drain_left.n6 drain_left.t15 9.9005
R327 drain_left.n8 drain_left.t3 9.9005
R328 drain_left.n8 drain_left.t0 9.9005
R329 drain_left.n3 drain_left.t16 9.9005
R330 drain_left.n3 drain_left.t14 9.9005
R331 drain_left.n1 drain_left.t9 9.9005
R332 drain_left.n1 drain_left.t22 9.9005
R333 drain_left.n0 drain_left.t8 9.9005
R334 drain_left.n0 drain_left.t2 9.9005
R335 drain_left.n20 drain_left.t4 9.9005
R336 drain_left.n20 drain_left.t7 9.9005
R337 drain_left.n18 drain_left.t21 9.9005
R338 drain_left.n18 drain_left.t23 9.9005
R339 drain_left.n16 drain_left.t19 9.9005
R340 drain_left.n16 drain_left.t20 9.9005
R341 drain_left.n14 drain_left.t13 9.9005
R342 drain_left.n14 drain_left.t18 9.9005
R343 drain_left.n12 drain_left.t10 9.9005
R344 drain_left.n12 drain_left.t11 9.9005
R345 drain_left.n11 drain_left.t5 9.9005
R346 drain_left.n11 drain_left.t6 9.9005
R347 drain_left drain_left.n21 6.45494
R348 drain_left.n9 drain_left.n7 0.802224
R349 drain_left.n4 drain_left.n2 0.802224
R350 drain_left.n15 drain_left.n13 0.802224
R351 drain_left.n17 drain_left.n15 0.802224
R352 drain_left.n19 drain_left.n17 0.802224
R353 drain_left.n21 drain_left.n19 0.802224
R354 drain_left.n10 drain_left.n9 0.346016
R355 drain_left.n10 drain_left.n4 0.346016
R356 minus.n9 minus.t17 172.163
R357 minus.n43 minus.t11 172.163
R358 minus.n33 minus.n32 161.3
R359 minus.n31 minus.n0 161.3
R360 minus.n30 minus.n29 161.3
R361 minus.n27 minus.n26 161.3
R362 minus.n25 minus.n2 161.3
R363 minus.n24 minus.n23 161.3
R364 minus.n22 minus.n3 161.3
R365 minus.n21 minus.n20 161.3
R366 minus.n19 minus.n4 161.3
R367 minus.n18 minus.n17 161.3
R368 minus.n16 minus.n5 161.3
R369 minus.n15 minus.n14 161.3
R370 minus.n13 minus.n6 161.3
R371 minus.n12 minus.n11 161.3
R372 minus.n67 minus.n66 161.3
R373 minus.n65 minus.n34 161.3
R374 minus.n64 minus.n63 161.3
R375 minus.n61 minus.n60 161.3
R376 minus.n59 minus.n36 161.3
R377 minus.n58 minus.n57 161.3
R378 minus.n56 minus.n37 161.3
R379 minus.n55 minus.n54 161.3
R380 minus.n53 minus.n38 161.3
R381 minus.n52 minus.n51 161.3
R382 minus.n50 minus.n39 161.3
R383 minus.n49 minus.n48 161.3
R384 minus.n47 minus.n40 161.3
R385 minus.n46 minus.n45 161.3
R386 minus.n8 minus.t16 145.805
R387 minus.n7 minus.t15 145.805
R388 minus.n12 minus.t13 145.805
R389 minus.n14 minus.t8 145.805
R390 minus.n18 minus.t12 145.805
R391 minus.n20 minus.t9 145.805
R392 minus.n24 minus.t4 145.805
R393 minus.n26 minus.t2 145.805
R394 minus.n1 minus.t1 145.805
R395 minus.n30 minus.t20 145.805
R396 minus.n32 minus.t14 145.805
R397 minus.n42 minus.t23 145.805
R398 minus.n41 minus.t19 145.805
R399 minus.n46 minus.t10 145.805
R400 minus.n48 minus.t3 145.805
R401 minus.n52 minus.t7 145.805
R402 minus.n54 minus.t22 145.805
R403 minus.n58 minus.t18 145.805
R404 minus.n60 minus.t6 145.805
R405 minus.n35 minus.t0 145.805
R406 minus.n64 minus.t5 145.805
R407 minus.n66 minus.t21 145.805
R408 minus.n28 minus.n1 80.6037
R409 minus.n10 minus.n7 80.6037
R410 minus.n62 minus.n35 80.6037
R411 minus.n44 minus.n41 80.6037
R412 minus.n8 minus.n7 48.2005
R413 minus.n12 minus.n7 48.2005
R414 minus.n26 minus.n1 48.2005
R415 minus.n30 minus.n1 48.2005
R416 minus.n42 minus.n41 48.2005
R417 minus.n46 minus.n41 48.2005
R418 minus.n60 minus.n35 48.2005
R419 minus.n64 minus.n35 48.2005
R420 minus.n32 minus.n31 46.0096
R421 minus.n66 minus.n65 46.0096
R422 minus.n10 minus.n9 45.1822
R423 minus.n44 minus.n43 45.1822
R424 minus.n14 minus.n13 44.549
R425 minus.n25 minus.n24 44.549
R426 minus.n48 minus.n47 44.549
R427 minus.n59 minus.n58 44.549
R428 minus.n18 minus.n5 34.3247
R429 minus.n20 minus.n3 34.3247
R430 minus.n52 minus.n39 34.3247
R431 minus.n54 minus.n37 34.3247
R432 minus.n68 minus.n33 33.5194
R433 minus.n20 minus.n19 24.1005
R434 minus.n19 minus.n18 24.1005
R435 minus.n53 minus.n52 24.1005
R436 minus.n54 minus.n53 24.1005
R437 minus.n9 minus.n8 14.1472
R438 minus.n43 minus.n42 14.1472
R439 minus.n14 minus.n5 13.8763
R440 minus.n24 minus.n3 13.8763
R441 minus.n48 minus.n39 13.8763
R442 minus.n58 minus.n37 13.8763
R443 minus.n68 minus.n67 6.60277
R444 minus.n13 minus.n12 3.65202
R445 minus.n26 minus.n25 3.65202
R446 minus.n47 minus.n46 3.65202
R447 minus.n60 minus.n59 3.65202
R448 minus.n31 minus.n30 2.19141
R449 minus.n65 minus.n64 2.19141
R450 minus.n29 minus.n28 0.285035
R451 minus.n28 minus.n27 0.285035
R452 minus.n11 minus.n10 0.285035
R453 minus.n45 minus.n44 0.285035
R454 minus.n62 minus.n61 0.285035
R455 minus.n63 minus.n62 0.285035
R456 minus.n33 minus.n0 0.189894
R457 minus.n29 minus.n0 0.189894
R458 minus.n27 minus.n2 0.189894
R459 minus.n23 minus.n2 0.189894
R460 minus.n23 minus.n22 0.189894
R461 minus.n22 minus.n21 0.189894
R462 minus.n21 minus.n4 0.189894
R463 minus.n17 minus.n4 0.189894
R464 minus.n17 minus.n16 0.189894
R465 minus.n16 minus.n15 0.189894
R466 minus.n15 minus.n6 0.189894
R467 minus.n11 minus.n6 0.189894
R468 minus.n45 minus.n40 0.189894
R469 minus.n49 minus.n40 0.189894
R470 minus.n50 minus.n49 0.189894
R471 minus.n51 minus.n50 0.189894
R472 minus.n51 minus.n38 0.189894
R473 minus.n55 minus.n38 0.189894
R474 minus.n56 minus.n55 0.189894
R475 minus.n57 minus.n56 0.189894
R476 minus.n57 minus.n36 0.189894
R477 minus.n61 minus.n36 0.189894
R478 minus.n63 minus.n34 0.189894
R479 minus.n67 minus.n34 0.189894
R480 minus minus.n68 0.188
R481 drain_right.n13 drain_right.n11 101.597
R482 drain_right.n7 drain_right.n5 101.597
R483 drain_right.n2 drain_right.n0 101.597
R484 drain_right.n13 drain_right.n12 100.796
R485 drain_right.n15 drain_right.n14 100.796
R486 drain_right.n17 drain_right.n16 100.796
R487 drain_right.n19 drain_right.n18 100.796
R488 drain_right.n21 drain_right.n20 100.796
R489 drain_right.n7 drain_right.n6 100.796
R490 drain_right.n9 drain_right.n8 100.796
R491 drain_right.n4 drain_right.n3 100.796
R492 drain_right.n2 drain_right.n1 100.796
R493 drain_right drain_right.n10 26.8545
R494 drain_right.n5 drain_right.t18 9.9005
R495 drain_right.n5 drain_right.t2 9.9005
R496 drain_right.n6 drain_right.t17 9.9005
R497 drain_right.n6 drain_right.t23 9.9005
R498 drain_right.n8 drain_right.t1 9.9005
R499 drain_right.n8 drain_right.t5 9.9005
R500 drain_right.n3 drain_right.t20 9.9005
R501 drain_right.n3 drain_right.t16 9.9005
R502 drain_right.n1 drain_right.t4 9.9005
R503 drain_right.n1 drain_right.t13 9.9005
R504 drain_right.n0 drain_right.t12 9.9005
R505 drain_right.n0 drain_right.t0 9.9005
R506 drain_right.n11 drain_right.t7 9.9005
R507 drain_right.n11 drain_right.t6 9.9005
R508 drain_right.n12 drain_right.t10 9.9005
R509 drain_right.n12 drain_right.t8 9.9005
R510 drain_right.n14 drain_right.t11 9.9005
R511 drain_right.n14 drain_right.t15 9.9005
R512 drain_right.n16 drain_right.t19 9.9005
R513 drain_right.n16 drain_right.t14 9.9005
R514 drain_right.n18 drain_right.t22 9.9005
R515 drain_right.n18 drain_right.t21 9.9005
R516 drain_right.n20 drain_right.t9 9.9005
R517 drain_right.n20 drain_right.t3 9.9005
R518 drain_right drain_right.n21 6.45494
R519 drain_right.n9 drain_right.n7 0.802224
R520 drain_right.n4 drain_right.n2 0.802224
R521 drain_right.n21 drain_right.n19 0.802224
R522 drain_right.n19 drain_right.n17 0.802224
R523 drain_right.n17 drain_right.n15 0.802224
R524 drain_right.n15 drain_right.n13 0.802224
R525 drain_right.n10 drain_right.n9 0.346016
R526 drain_right.n10 drain_right.n4 0.346016
C0 drain_left source 8.87966f
C1 minus drain_right 2.90277f
C2 plus drain_left 3.21598f
C3 minus source 3.65886f
C4 drain_right source 8.88171f
C5 plus minus 5.21759f
C6 plus drain_right 0.478436f
C7 plus source 3.67282f
C8 minus drain_left 0.180449f
C9 drain_left drain_right 1.7173f
C10 drain_right a_n3134_n1288# 5.72051f
C11 drain_left a_n3134_n1288# 6.17981f
C12 source a_n3134_n1288# 3.603836f
C13 minus a_n3134_n1288# 11.791546f
C14 plus a_n3134_n1288# 13.229771f
C15 drain_right.t12 a_n3134_n1288# 0.043753f
C16 drain_right.t0 a_n3134_n1288# 0.043753f
C17 drain_right.n0 a_n3134_n1288# 0.27776f
C18 drain_right.t4 a_n3134_n1288# 0.043753f
C19 drain_right.t13 a_n3134_n1288# 0.043753f
C20 drain_right.n1 a_n3134_n1288# 0.274871f
C21 drain_right.n2 a_n3134_n1288# 0.718107f
C22 drain_right.t20 a_n3134_n1288# 0.043753f
C23 drain_right.t16 a_n3134_n1288# 0.043753f
C24 drain_right.n3 a_n3134_n1288# 0.274871f
C25 drain_right.n4 a_n3134_n1288# 0.316085f
C26 drain_right.t18 a_n3134_n1288# 0.043753f
C27 drain_right.t2 a_n3134_n1288# 0.043753f
C28 drain_right.n5 a_n3134_n1288# 0.27776f
C29 drain_right.t17 a_n3134_n1288# 0.043753f
C30 drain_right.t23 a_n3134_n1288# 0.043753f
C31 drain_right.n6 a_n3134_n1288# 0.274871f
C32 drain_right.n7 a_n3134_n1288# 0.718108f
C33 drain_right.t1 a_n3134_n1288# 0.043753f
C34 drain_right.t5 a_n3134_n1288# 0.043753f
C35 drain_right.n8 a_n3134_n1288# 0.274871f
C36 drain_right.n9 a_n3134_n1288# 0.316085f
C37 drain_right.n10 a_n3134_n1288# 1.10972f
C38 drain_right.t7 a_n3134_n1288# 0.043753f
C39 drain_right.t6 a_n3134_n1288# 0.043753f
C40 drain_right.n11 a_n3134_n1288# 0.277761f
C41 drain_right.t10 a_n3134_n1288# 0.043753f
C42 drain_right.t8 a_n3134_n1288# 0.043753f
C43 drain_right.n12 a_n3134_n1288# 0.274872f
C44 drain_right.n13 a_n3134_n1288# 0.718105f
C45 drain_right.t11 a_n3134_n1288# 0.043753f
C46 drain_right.t15 a_n3134_n1288# 0.043753f
C47 drain_right.n14 a_n3134_n1288# 0.274872f
C48 drain_right.n15 a_n3134_n1288# 0.354922f
C49 drain_right.t19 a_n3134_n1288# 0.043753f
C50 drain_right.t14 a_n3134_n1288# 0.043753f
C51 drain_right.n16 a_n3134_n1288# 0.274872f
C52 drain_right.n17 a_n3134_n1288# 0.354922f
C53 drain_right.t22 a_n3134_n1288# 0.043753f
C54 drain_right.t21 a_n3134_n1288# 0.043753f
C55 drain_right.n18 a_n3134_n1288# 0.274872f
C56 drain_right.n19 a_n3134_n1288# 0.354922f
C57 drain_right.t9 a_n3134_n1288# 0.043753f
C58 drain_right.t3 a_n3134_n1288# 0.043753f
C59 drain_right.n20 a_n3134_n1288# 0.274872f
C60 drain_right.n21 a_n3134_n1288# 0.596323f
C61 minus.n0 a_n3134_n1288# 0.043014f
C62 minus.t1 a_n3134_n1288# 0.159841f
C63 minus.n1 a_n3134_n1288# 0.122948f
C64 minus.t20 a_n3134_n1288# 0.159841f
C65 minus.n2 a_n3134_n1288# 0.043014f
C66 minus.n3 a_n3134_n1288# 0.009761f
C67 minus.t4 a_n3134_n1288# 0.159841f
C68 minus.n4 a_n3134_n1288# 0.043014f
C69 minus.n5 a_n3134_n1288# 0.009761f
C70 minus.t12 a_n3134_n1288# 0.159841f
C71 minus.n6 a_n3134_n1288# 0.043014f
C72 minus.t15 a_n3134_n1288# 0.159841f
C73 minus.n7 a_n3134_n1288# 0.122948f
C74 minus.t13 a_n3134_n1288# 0.159841f
C75 minus.t17 a_n3134_n1288# 0.177163f
C76 minus.t16 a_n3134_n1288# 0.159841f
C77 minus.n8 a_n3134_n1288# 0.122388f
C78 minus.n9 a_n3134_n1288# 0.097697f
C79 minus.n10 a_n3134_n1288# 0.208166f
C80 minus.n11 a_n3134_n1288# 0.057396f
C81 minus.n12 a_n3134_n1288# 0.113851f
C82 minus.n13 a_n3134_n1288# 0.009761f
C83 minus.t8 a_n3134_n1288# 0.159841f
C84 minus.n14 a_n3134_n1288# 0.115044f
C85 minus.n15 a_n3134_n1288# 0.043014f
C86 minus.n16 a_n3134_n1288# 0.043014f
C87 minus.n17 a_n3134_n1288# 0.043014f
C88 minus.n18 a_n3134_n1288# 0.115044f
C89 minus.n19 a_n3134_n1288# 0.009761f
C90 minus.t9 a_n3134_n1288# 0.159841f
C91 minus.n20 a_n3134_n1288# 0.115044f
C92 minus.n21 a_n3134_n1288# 0.043014f
C93 minus.n22 a_n3134_n1288# 0.043014f
C94 minus.n23 a_n3134_n1288# 0.043014f
C95 minus.n24 a_n3134_n1288# 0.115044f
C96 minus.n25 a_n3134_n1288# 0.009761f
C97 minus.t2 a_n3134_n1288# 0.159841f
C98 minus.n26 a_n3134_n1288# 0.113851f
C99 minus.n27 a_n3134_n1288# 0.057396f
C100 minus.n28 a_n3134_n1288# 0.057262f
C101 minus.n29 a_n3134_n1288# 0.057396f
C102 minus.n30 a_n3134_n1288# 0.113585f
C103 minus.n31 a_n3134_n1288# 0.009761f
C104 minus.t14 a_n3134_n1288# 0.159841f
C105 minus.n32 a_n3134_n1288# 0.11279f
C106 minus.n33 a_n3134_n1288# 1.34913f
C107 minus.n34 a_n3134_n1288# 0.043014f
C108 minus.t0 a_n3134_n1288# 0.159841f
C109 minus.n35 a_n3134_n1288# 0.122948f
C110 minus.n36 a_n3134_n1288# 0.043014f
C111 minus.n37 a_n3134_n1288# 0.009761f
C112 minus.n38 a_n3134_n1288# 0.043014f
C113 minus.n39 a_n3134_n1288# 0.009761f
C114 minus.n40 a_n3134_n1288# 0.043014f
C115 minus.t19 a_n3134_n1288# 0.159841f
C116 minus.n41 a_n3134_n1288# 0.122948f
C117 minus.t11 a_n3134_n1288# 0.177163f
C118 minus.t23 a_n3134_n1288# 0.159841f
C119 minus.n42 a_n3134_n1288# 0.122388f
C120 minus.n43 a_n3134_n1288# 0.097697f
C121 minus.n44 a_n3134_n1288# 0.208166f
C122 minus.n45 a_n3134_n1288# 0.057396f
C123 minus.t10 a_n3134_n1288# 0.159841f
C124 minus.n46 a_n3134_n1288# 0.113851f
C125 minus.n47 a_n3134_n1288# 0.009761f
C126 minus.t3 a_n3134_n1288# 0.159841f
C127 minus.n48 a_n3134_n1288# 0.115044f
C128 minus.n49 a_n3134_n1288# 0.043014f
C129 minus.n50 a_n3134_n1288# 0.043014f
C130 minus.n51 a_n3134_n1288# 0.043014f
C131 minus.t7 a_n3134_n1288# 0.159841f
C132 minus.n52 a_n3134_n1288# 0.115044f
C133 minus.n53 a_n3134_n1288# 0.009761f
C134 minus.t22 a_n3134_n1288# 0.159841f
C135 minus.n54 a_n3134_n1288# 0.115044f
C136 minus.n55 a_n3134_n1288# 0.043014f
C137 minus.n56 a_n3134_n1288# 0.043014f
C138 minus.n57 a_n3134_n1288# 0.043014f
C139 minus.t18 a_n3134_n1288# 0.159841f
C140 minus.n58 a_n3134_n1288# 0.115044f
C141 minus.n59 a_n3134_n1288# 0.009761f
C142 minus.t6 a_n3134_n1288# 0.159841f
C143 minus.n60 a_n3134_n1288# 0.113851f
C144 minus.n61 a_n3134_n1288# 0.057396f
C145 minus.n62 a_n3134_n1288# 0.057262f
C146 minus.n63 a_n3134_n1288# 0.057396f
C147 minus.t5 a_n3134_n1288# 0.159841f
C148 minus.n64 a_n3134_n1288# 0.113585f
C149 minus.n65 a_n3134_n1288# 0.009761f
C150 minus.t21 a_n3134_n1288# 0.159841f
C151 minus.n66 a_n3134_n1288# 0.11279f
C152 minus.n67 a_n3134_n1288# 0.291576f
C153 minus.n68 a_n3134_n1288# 1.64711f
C154 drain_left.t8 a_n3134_n1288# 0.044458f
C155 drain_left.t2 a_n3134_n1288# 0.044458f
C156 drain_left.n0 a_n3134_n1288# 0.282231f
C157 drain_left.t9 a_n3134_n1288# 0.044458f
C158 drain_left.t22 a_n3134_n1288# 0.044458f
C159 drain_left.n1 a_n3134_n1288# 0.279296f
C160 drain_left.n2 a_n3134_n1288# 0.729668f
C161 drain_left.t16 a_n3134_n1288# 0.044458f
C162 drain_left.t14 a_n3134_n1288# 0.044458f
C163 drain_left.n3 a_n3134_n1288# 0.279296f
C164 drain_left.n4 a_n3134_n1288# 0.321174f
C165 drain_left.t12 a_n3134_n1288# 0.044458f
C166 drain_left.t1 a_n3134_n1288# 0.044458f
C167 drain_left.n5 a_n3134_n1288# 0.282231f
C168 drain_left.t17 a_n3134_n1288# 0.044458f
C169 drain_left.t15 a_n3134_n1288# 0.044458f
C170 drain_left.n6 a_n3134_n1288# 0.279296f
C171 drain_left.n7 a_n3134_n1288# 0.729668f
C172 drain_left.t3 a_n3134_n1288# 0.044458f
C173 drain_left.t0 a_n3134_n1288# 0.044458f
C174 drain_left.n8 a_n3134_n1288# 0.279296f
C175 drain_left.n9 a_n3134_n1288# 0.321174f
C176 drain_left.n10 a_n3134_n1288# 1.18203f
C177 drain_left.t5 a_n3134_n1288# 0.044458f
C178 drain_left.t6 a_n3134_n1288# 0.044458f
C179 drain_left.n11 a_n3134_n1288# 0.282233f
C180 drain_left.t10 a_n3134_n1288# 0.044458f
C181 drain_left.t11 a_n3134_n1288# 0.044458f
C182 drain_left.n12 a_n3134_n1288# 0.279297f
C183 drain_left.n13 a_n3134_n1288# 0.729666f
C184 drain_left.t13 a_n3134_n1288# 0.044458f
C185 drain_left.t18 a_n3134_n1288# 0.044458f
C186 drain_left.n14 a_n3134_n1288# 0.279297f
C187 drain_left.n15 a_n3134_n1288# 0.360635f
C188 drain_left.t19 a_n3134_n1288# 0.044458f
C189 drain_left.t20 a_n3134_n1288# 0.044458f
C190 drain_left.n16 a_n3134_n1288# 0.279297f
C191 drain_left.n17 a_n3134_n1288# 0.360635f
C192 drain_left.t21 a_n3134_n1288# 0.044458f
C193 drain_left.t23 a_n3134_n1288# 0.044458f
C194 drain_left.n18 a_n3134_n1288# 0.279297f
C195 drain_left.n19 a_n3134_n1288# 0.360635f
C196 drain_left.t4 a_n3134_n1288# 0.044458f
C197 drain_left.t7 a_n3134_n1288# 0.044458f
C198 drain_left.n20 a_n3134_n1288# 0.279297f
C199 drain_left.n21 a_n3134_n1288# 0.605922f
C200 source.n0 a_n3134_n1288# 0.047451f
C201 source.n1 a_n3134_n1288# 0.104991f
C202 source.t45 a_n3134_n1288# 0.07879f
C203 source.n2 a_n3134_n1288# 0.08217f
C204 source.n3 a_n3134_n1288# 0.026488f
C205 source.n4 a_n3134_n1288# 0.01747f
C206 source.n5 a_n3134_n1288# 0.231425f
C207 source.n6 a_n3134_n1288# 0.052017f
C208 source.n7 a_n3134_n1288# 0.538888f
C209 source.t22 a_n3134_n1288# 0.051381f
C210 source.t31 a_n3134_n1288# 0.051381f
C211 source.n8 a_n3134_n1288# 0.274683f
C212 source.n9 a_n3134_n1288# 0.420722f
C213 source.t23 a_n3134_n1288# 0.051381f
C214 source.t24 a_n3134_n1288# 0.051381f
C215 source.n10 a_n3134_n1288# 0.274683f
C216 source.n11 a_n3134_n1288# 0.420722f
C217 source.t37 a_n3134_n1288# 0.051381f
C218 source.t33 a_n3134_n1288# 0.051381f
C219 source.n12 a_n3134_n1288# 0.274683f
C220 source.n13 a_n3134_n1288# 0.420722f
C221 source.t39 a_n3134_n1288# 0.051381f
C222 source.t43 a_n3134_n1288# 0.051381f
C223 source.n14 a_n3134_n1288# 0.274683f
C224 source.n15 a_n3134_n1288# 0.420722f
C225 source.t38 a_n3134_n1288# 0.051381f
C226 source.t40 a_n3134_n1288# 0.051381f
C227 source.n16 a_n3134_n1288# 0.274683f
C228 source.n17 a_n3134_n1288# 0.420722f
C229 source.n18 a_n3134_n1288# 0.047451f
C230 source.n19 a_n3134_n1288# 0.104991f
C231 source.t41 a_n3134_n1288# 0.07879f
C232 source.n20 a_n3134_n1288# 0.08217f
C233 source.n21 a_n3134_n1288# 0.026488f
C234 source.n22 a_n3134_n1288# 0.01747f
C235 source.n23 a_n3134_n1288# 0.231425f
C236 source.n24 a_n3134_n1288# 0.052017f
C237 source.n25 a_n3134_n1288# 0.159966f
C238 source.n26 a_n3134_n1288# 0.047451f
C239 source.n27 a_n3134_n1288# 0.104991f
C240 source.t6 a_n3134_n1288# 0.07879f
C241 source.n28 a_n3134_n1288# 0.08217f
C242 source.n29 a_n3134_n1288# 0.026488f
C243 source.n30 a_n3134_n1288# 0.01747f
C244 source.n31 a_n3134_n1288# 0.231425f
C245 source.n32 a_n3134_n1288# 0.052017f
C246 source.n33 a_n3134_n1288# 0.159966f
C247 source.t13 a_n3134_n1288# 0.051381f
C248 source.t17 a_n3134_n1288# 0.051381f
C249 source.n34 a_n3134_n1288# 0.274683f
C250 source.n35 a_n3134_n1288# 0.420722f
C251 source.t47 a_n3134_n1288# 0.051381f
C252 source.t11 a_n3134_n1288# 0.051381f
C253 source.n36 a_n3134_n1288# 0.274683f
C254 source.n37 a_n3134_n1288# 0.420722f
C255 source.t3 a_n3134_n1288# 0.051381f
C256 source.t19 a_n3134_n1288# 0.051381f
C257 source.n38 a_n3134_n1288# 0.274683f
C258 source.n39 a_n3134_n1288# 0.420722f
C259 source.t5 a_n3134_n1288# 0.051381f
C260 source.t15 a_n3134_n1288# 0.051381f
C261 source.n40 a_n3134_n1288# 0.274683f
C262 source.n41 a_n3134_n1288# 0.420722f
C263 source.t20 a_n3134_n1288# 0.051381f
C264 source.t1 a_n3134_n1288# 0.051381f
C265 source.n42 a_n3134_n1288# 0.274683f
C266 source.n43 a_n3134_n1288# 0.420722f
C267 source.n44 a_n3134_n1288# 0.047451f
C268 source.n45 a_n3134_n1288# 0.104991f
C269 source.t7 a_n3134_n1288# 0.07879f
C270 source.n46 a_n3134_n1288# 0.08217f
C271 source.n47 a_n3134_n1288# 0.026488f
C272 source.n48 a_n3134_n1288# 0.01747f
C273 source.n49 a_n3134_n1288# 0.231425f
C274 source.n50 a_n3134_n1288# 0.052017f
C275 source.n51 a_n3134_n1288# 0.848131f
C276 source.n52 a_n3134_n1288# 0.047451f
C277 source.n53 a_n3134_n1288# 0.104991f
C278 source.t26 a_n3134_n1288# 0.07879f
C279 source.n54 a_n3134_n1288# 0.08217f
C280 source.n55 a_n3134_n1288# 0.026488f
C281 source.n56 a_n3134_n1288# 0.01747f
C282 source.n57 a_n3134_n1288# 0.231425f
C283 source.n58 a_n3134_n1288# 0.052017f
C284 source.n59 a_n3134_n1288# 0.848131f
C285 source.t32 a_n3134_n1288# 0.051381f
C286 source.t27 a_n3134_n1288# 0.051381f
C287 source.n60 a_n3134_n1288# 0.274681f
C288 source.n61 a_n3134_n1288# 0.420724f
C289 source.t36 a_n3134_n1288# 0.051381f
C290 source.t28 a_n3134_n1288# 0.051381f
C291 source.n62 a_n3134_n1288# 0.274681f
C292 source.n63 a_n3134_n1288# 0.420724f
C293 source.t29 a_n3134_n1288# 0.051381f
C294 source.t34 a_n3134_n1288# 0.051381f
C295 source.n64 a_n3134_n1288# 0.274681f
C296 source.n65 a_n3134_n1288# 0.420724f
C297 source.t30 a_n3134_n1288# 0.051381f
C298 source.t35 a_n3134_n1288# 0.051381f
C299 source.n66 a_n3134_n1288# 0.274681f
C300 source.n67 a_n3134_n1288# 0.420724f
C301 source.t42 a_n3134_n1288# 0.051381f
C302 source.t44 a_n3134_n1288# 0.051381f
C303 source.n68 a_n3134_n1288# 0.274681f
C304 source.n69 a_n3134_n1288# 0.420724f
C305 source.n70 a_n3134_n1288# 0.047451f
C306 source.n71 a_n3134_n1288# 0.104991f
C307 source.t25 a_n3134_n1288# 0.07879f
C308 source.n72 a_n3134_n1288# 0.08217f
C309 source.n73 a_n3134_n1288# 0.026488f
C310 source.n74 a_n3134_n1288# 0.01747f
C311 source.n75 a_n3134_n1288# 0.231425f
C312 source.n76 a_n3134_n1288# 0.052017f
C313 source.n77 a_n3134_n1288# 0.159966f
C314 source.n78 a_n3134_n1288# 0.047451f
C315 source.n79 a_n3134_n1288# 0.104991f
C316 source.t2 a_n3134_n1288# 0.07879f
C317 source.n80 a_n3134_n1288# 0.08217f
C318 source.n81 a_n3134_n1288# 0.026488f
C319 source.n82 a_n3134_n1288# 0.01747f
C320 source.n83 a_n3134_n1288# 0.231425f
C321 source.n84 a_n3134_n1288# 0.052017f
C322 source.n85 a_n3134_n1288# 0.159966f
C323 source.t4 a_n3134_n1288# 0.051381f
C324 source.t21 a_n3134_n1288# 0.051381f
C325 source.n86 a_n3134_n1288# 0.274681f
C326 source.n87 a_n3134_n1288# 0.420724f
C327 source.t0 a_n3134_n1288# 0.051381f
C328 source.t12 a_n3134_n1288# 0.051381f
C329 source.n88 a_n3134_n1288# 0.274681f
C330 source.n89 a_n3134_n1288# 0.420724f
C331 source.t46 a_n3134_n1288# 0.051381f
C332 source.t14 a_n3134_n1288# 0.051381f
C333 source.n90 a_n3134_n1288# 0.274681f
C334 source.n91 a_n3134_n1288# 0.420724f
C335 source.t8 a_n3134_n1288# 0.051381f
C336 source.t10 a_n3134_n1288# 0.051381f
C337 source.n92 a_n3134_n1288# 0.274681f
C338 source.n93 a_n3134_n1288# 0.420724f
C339 source.t9 a_n3134_n1288# 0.051381f
C340 source.t16 a_n3134_n1288# 0.051381f
C341 source.n94 a_n3134_n1288# 0.274681f
C342 source.n95 a_n3134_n1288# 0.420724f
C343 source.n96 a_n3134_n1288# 0.047451f
C344 source.n97 a_n3134_n1288# 0.104991f
C345 source.t18 a_n3134_n1288# 0.07879f
C346 source.n98 a_n3134_n1288# 0.08217f
C347 source.n99 a_n3134_n1288# 0.026488f
C348 source.n100 a_n3134_n1288# 0.01747f
C349 source.n101 a_n3134_n1288# 0.231425f
C350 source.n102 a_n3134_n1288# 0.052017f
C351 source.n103 a_n3134_n1288# 0.364955f
C352 source.n104 a_n3134_n1288# 0.815542f
C353 plus.n0 a_n3134_n1288# 0.044435f
C354 plus.t16 a_n3134_n1288# 0.165122f
C355 plus.t19 a_n3134_n1288# 0.165122f
C356 plus.n1 a_n3134_n1288# 0.059292f
C357 plus.t0 a_n3134_n1288# 0.165122f
C358 plus.n2 a_n3134_n1288# 0.059154f
C359 plus.t2 a_n3134_n1288# 0.165122f
C360 plus.n3 a_n3134_n1288# 0.059292f
C361 plus.t3 a_n3134_n1288# 0.165122f
C362 plus.n4 a_n3134_n1288# 0.118845f
C363 plus.n5 a_n3134_n1288# 0.044435f
C364 plus.t4 a_n3134_n1288# 0.165122f
C365 plus.t5 a_n3134_n1288# 0.165122f
C366 plus.n6 a_n3134_n1288# 0.118845f
C367 plus.n7 a_n3134_n1288# 0.044435f
C368 plus.t10 a_n3134_n1288# 0.165122f
C369 plus.t12 a_n3134_n1288# 0.165122f
C370 plus.n8 a_n3134_n1288# 0.117612f
C371 plus.t18 a_n3134_n1288# 0.183016f
C372 plus.n9 a_n3134_n1288# 0.100925f
C373 plus.t13 a_n3134_n1288# 0.165122f
C374 plus.t17 a_n3134_n1288# 0.165122f
C375 plus.n10 a_n3134_n1288# 0.126431f
C376 plus.n11 a_n3134_n1288# 0.12701f
C377 plus.n12 a_n3134_n1288# 0.215044f
C378 plus.n13 a_n3134_n1288# 0.059292f
C379 plus.n14 a_n3134_n1288# 0.044435f
C380 plus.n15 a_n3134_n1288# 0.010083f
C381 plus.n16 a_n3134_n1288# 0.118845f
C382 plus.n17 a_n3134_n1288# 0.010083f
C383 plus.n18 a_n3134_n1288# 0.044435f
C384 plus.n19 a_n3134_n1288# 0.044435f
C385 plus.n20 a_n3134_n1288# 0.044435f
C386 plus.n21 a_n3134_n1288# 0.010083f
C387 plus.n22 a_n3134_n1288# 0.118845f
C388 plus.n23 a_n3134_n1288# 0.010083f
C389 plus.n24 a_n3134_n1288# 0.044435f
C390 plus.n25 a_n3134_n1288# 0.044435f
C391 plus.n26 a_n3134_n1288# 0.044435f
C392 plus.n27 a_n3134_n1288# 0.010083f
C393 plus.n28 a_n3134_n1288# 0.117612f
C394 plus.n29 a_n3134_n1288# 0.12701f
C395 plus.n30 a_n3134_n1288# 0.117338f
C396 plus.n31 a_n3134_n1288# 0.010083f
C397 plus.n32 a_n3134_n1288# 0.116516f
C398 plus.n33 a_n3134_n1288# 0.328949f
C399 plus.n34 a_n3134_n1288# 0.044435f
C400 plus.t15 a_n3134_n1288# 0.165122f
C401 plus.n35 a_n3134_n1288# 0.059292f
C402 plus.t21 a_n3134_n1288# 0.165122f
C403 plus.n36 a_n3134_n1288# 0.059154f
C404 plus.t14 a_n3134_n1288# 0.165122f
C405 plus.n37 a_n3134_n1288# 0.059292f
C406 plus.t1 a_n3134_n1288# 0.165122f
C407 plus.t7 a_n3134_n1288# 0.165122f
C408 plus.n38 a_n3134_n1288# 0.118845f
C409 plus.n39 a_n3134_n1288# 0.044435f
C410 plus.t9 a_n3134_n1288# 0.165122f
C411 plus.t20 a_n3134_n1288# 0.165122f
C412 plus.n40 a_n3134_n1288# 0.118845f
C413 plus.n41 a_n3134_n1288# 0.044435f
C414 plus.t23 a_n3134_n1288# 0.165122f
C415 plus.t6 a_n3134_n1288# 0.165122f
C416 plus.n42 a_n3134_n1288# 0.117612f
C417 plus.t22 a_n3134_n1288# 0.183016f
C418 plus.n43 a_n3134_n1288# 0.100925f
C419 plus.t8 a_n3134_n1288# 0.165122f
C420 plus.t11 a_n3134_n1288# 0.165122f
C421 plus.n44 a_n3134_n1288# 0.126431f
C422 plus.n45 a_n3134_n1288# 0.12701f
C423 plus.n46 a_n3134_n1288# 0.215044f
C424 plus.n47 a_n3134_n1288# 0.059292f
C425 plus.n48 a_n3134_n1288# 0.044435f
C426 plus.n49 a_n3134_n1288# 0.010083f
C427 plus.n50 a_n3134_n1288# 0.118845f
C428 plus.n51 a_n3134_n1288# 0.010083f
C429 plus.n52 a_n3134_n1288# 0.044435f
C430 plus.n53 a_n3134_n1288# 0.044435f
C431 plus.n54 a_n3134_n1288# 0.044435f
C432 plus.n55 a_n3134_n1288# 0.010083f
C433 plus.n56 a_n3134_n1288# 0.118845f
C434 plus.n57 a_n3134_n1288# 0.010083f
C435 plus.n58 a_n3134_n1288# 0.044435f
C436 plus.n59 a_n3134_n1288# 0.044435f
C437 plus.n60 a_n3134_n1288# 0.044435f
C438 plus.n61 a_n3134_n1288# 0.010083f
C439 plus.n62 a_n3134_n1288# 0.117612f
C440 plus.n63 a_n3134_n1288# 0.12701f
C441 plus.n64 a_n3134_n1288# 0.117338f
C442 plus.n65 a_n3134_n1288# 0.010083f
C443 plus.n66 a_n3134_n1288# 0.116516f
C444 plus.n67 a_n3134_n1288# 1.32444f
.ends

