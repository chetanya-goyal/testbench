* NGSPICE file created from diffpair255.ext - technology: sky130A

.subckt diffpair255 minus drain_right drain_left source plus
X0 a_n1458_n2088# a_n1458_n2088# a_n1458_n2088# a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.2
X1 drain_right.t11 minus.t0 source.t14 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X2 source.t13 minus.t1 drain_right.t10 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X3 drain_left.t11 plus.t0 source.t6 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X4 source.t10 plus.t1 drain_left.t10 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X5 source.t12 minus.t2 drain_right.t9 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X6 source.t4 plus.t2 drain_left.t9 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X7 source.t18 minus.t3 drain_right.t8 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X8 a_n1458_n2088# a_n1458_n2088# a_n1458_n2088# a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X9 drain_left.t8 plus.t3 source.t5 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X10 source.t9 plus.t4 drain_left.t7 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X11 drain_left.t6 plus.t5 source.t0 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X12 drain_left.t5 plus.t6 source.t8 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X13 drain_left.t4 plus.t7 source.t11 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X14 drain_right.t7 minus.t4 source.t21 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X15 drain_right.t6 minus.t5 source.t20 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X16 source.t1 plus.t8 drain_left.t3 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X17 a_n1458_n2088# a_n1458_n2088# a_n1458_n2088# a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X18 a_n1458_n2088# a_n1458_n2088# a_n1458_n2088# a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X19 source.t2 plus.t9 drain_left.t2 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X20 drain_left.t1 plus.t10 source.t3 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X21 source.t22 minus.t6 drain_right.t5 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X22 source.t19 minus.t7 drain_right.t4 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X23 source.t15 minus.t8 drain_right.t3 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X24 drain_right.t2 minus.t9 source.t17 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X25 drain_right.t1 minus.t10 source.t16 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X26 source.t7 plus.t11 drain_left.t0 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X27 drain_right.t0 minus.t11 source.t23 a_n1458_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
R0 minus.n11 minus.t2 927.12
R1 minus.n2 minus.t4 927.12
R2 minus.n24 minus.t11 927.12
R3 minus.n15 minus.t7 927.12
R4 minus.n10 minus.t5 879.65
R5 minus.n8 minus.t8 879.65
R6 minus.n1 minus.t0 879.65
R7 minus.n3 minus.t3 879.65
R8 minus.n23 minus.t1 879.65
R9 minus.n21 minus.t9 879.65
R10 minus.n14 minus.t6 879.65
R11 minus.n16 minus.t10 879.65
R12 minus.n5 minus.n2 161.489
R13 minus.n18 minus.n15 161.489
R14 minus.n12 minus.n11 161.3
R15 minus.n9 minus.n0 161.3
R16 minus.n7 minus.n6 161.3
R17 minus.n5 minus.n4 161.3
R18 minus.n25 minus.n24 161.3
R19 minus.n22 minus.n13 161.3
R20 minus.n20 minus.n19 161.3
R21 minus.n18 minus.n17 161.3
R22 minus.n10 minus.n9 43.0884
R23 minus.n4 minus.n3 43.0884
R24 minus.n17 minus.n16 43.0884
R25 minus.n23 minus.n22 43.0884
R26 minus.n8 minus.n7 38.7066
R27 minus.n7 minus.n1 38.7066
R28 minus.n20 minus.n14 38.7066
R29 minus.n21 minus.n20 38.7066
R30 minus.n9 minus.n8 34.3247
R31 minus.n4 minus.n1 34.3247
R32 minus.n17 minus.n14 34.3247
R33 minus.n22 minus.n21 34.3247
R34 minus.n26 minus.n12 30.0535
R35 minus.n11 minus.n10 29.9429
R36 minus.n3 minus.n2 29.9429
R37 minus.n16 minus.n15 29.9429
R38 minus.n24 minus.n23 29.9429
R39 minus.n26 minus.n25 6.45505
R40 minus.n12 minus.n0 0.189894
R41 minus.n6 minus.n0 0.189894
R42 minus.n6 minus.n5 0.189894
R43 minus.n19 minus.n18 0.189894
R44 minus.n19 minus.n13 0.189894
R45 minus.n25 minus.n13 0.189894
R46 minus minus.n26 0.188
R47 source.n266 source.n240 289.615
R48 source.n230 source.n204 289.615
R49 source.n198 source.n172 289.615
R50 source.n162 source.n136 289.615
R51 source.n26 source.n0 289.615
R52 source.n62 source.n36 289.615
R53 source.n94 source.n68 289.615
R54 source.n130 source.n104 289.615
R55 source.n251 source.n250 185
R56 source.n248 source.n247 185
R57 source.n257 source.n256 185
R58 source.n259 source.n258 185
R59 source.n244 source.n243 185
R60 source.n265 source.n264 185
R61 source.n267 source.n266 185
R62 source.n215 source.n214 185
R63 source.n212 source.n211 185
R64 source.n221 source.n220 185
R65 source.n223 source.n222 185
R66 source.n208 source.n207 185
R67 source.n229 source.n228 185
R68 source.n231 source.n230 185
R69 source.n183 source.n182 185
R70 source.n180 source.n179 185
R71 source.n189 source.n188 185
R72 source.n191 source.n190 185
R73 source.n176 source.n175 185
R74 source.n197 source.n196 185
R75 source.n199 source.n198 185
R76 source.n147 source.n146 185
R77 source.n144 source.n143 185
R78 source.n153 source.n152 185
R79 source.n155 source.n154 185
R80 source.n140 source.n139 185
R81 source.n161 source.n160 185
R82 source.n163 source.n162 185
R83 source.n27 source.n26 185
R84 source.n25 source.n24 185
R85 source.n4 source.n3 185
R86 source.n19 source.n18 185
R87 source.n17 source.n16 185
R88 source.n8 source.n7 185
R89 source.n11 source.n10 185
R90 source.n63 source.n62 185
R91 source.n61 source.n60 185
R92 source.n40 source.n39 185
R93 source.n55 source.n54 185
R94 source.n53 source.n52 185
R95 source.n44 source.n43 185
R96 source.n47 source.n46 185
R97 source.n95 source.n94 185
R98 source.n93 source.n92 185
R99 source.n72 source.n71 185
R100 source.n87 source.n86 185
R101 source.n85 source.n84 185
R102 source.n76 source.n75 185
R103 source.n79 source.n78 185
R104 source.n131 source.n130 185
R105 source.n129 source.n128 185
R106 source.n108 source.n107 185
R107 source.n123 source.n122 185
R108 source.n121 source.n120 185
R109 source.n112 source.n111 185
R110 source.n115 source.n114 185
R111 source.t23 source.n249 147.661
R112 source.t19 source.n213 147.661
R113 source.t11 source.n181 147.661
R114 source.t10 source.n145 147.661
R115 source.t5 source.n9 147.661
R116 source.t9 source.n45 147.661
R117 source.t21 source.n77 147.661
R118 source.t12 source.n113 147.661
R119 source.n250 source.n247 104.615
R120 source.n257 source.n247 104.615
R121 source.n258 source.n257 104.615
R122 source.n258 source.n243 104.615
R123 source.n265 source.n243 104.615
R124 source.n266 source.n265 104.615
R125 source.n214 source.n211 104.615
R126 source.n221 source.n211 104.615
R127 source.n222 source.n221 104.615
R128 source.n222 source.n207 104.615
R129 source.n229 source.n207 104.615
R130 source.n230 source.n229 104.615
R131 source.n182 source.n179 104.615
R132 source.n189 source.n179 104.615
R133 source.n190 source.n189 104.615
R134 source.n190 source.n175 104.615
R135 source.n197 source.n175 104.615
R136 source.n198 source.n197 104.615
R137 source.n146 source.n143 104.615
R138 source.n153 source.n143 104.615
R139 source.n154 source.n153 104.615
R140 source.n154 source.n139 104.615
R141 source.n161 source.n139 104.615
R142 source.n162 source.n161 104.615
R143 source.n26 source.n25 104.615
R144 source.n25 source.n3 104.615
R145 source.n18 source.n3 104.615
R146 source.n18 source.n17 104.615
R147 source.n17 source.n7 104.615
R148 source.n10 source.n7 104.615
R149 source.n62 source.n61 104.615
R150 source.n61 source.n39 104.615
R151 source.n54 source.n39 104.615
R152 source.n54 source.n53 104.615
R153 source.n53 source.n43 104.615
R154 source.n46 source.n43 104.615
R155 source.n94 source.n93 104.615
R156 source.n93 source.n71 104.615
R157 source.n86 source.n71 104.615
R158 source.n86 source.n85 104.615
R159 source.n85 source.n75 104.615
R160 source.n78 source.n75 104.615
R161 source.n130 source.n129 104.615
R162 source.n129 source.n107 104.615
R163 source.n122 source.n107 104.615
R164 source.n122 source.n121 104.615
R165 source.n121 source.n111 104.615
R166 source.n114 source.n111 104.615
R167 source.n250 source.t23 52.3082
R168 source.n214 source.t19 52.3082
R169 source.n182 source.t11 52.3082
R170 source.n146 source.t10 52.3082
R171 source.n10 source.t5 52.3082
R172 source.n46 source.t9 52.3082
R173 source.n78 source.t21 52.3082
R174 source.n114 source.t12 52.3082
R175 source.n33 source.n32 50.512
R176 source.n35 source.n34 50.512
R177 source.n101 source.n100 50.512
R178 source.n103 source.n102 50.512
R179 source.n239 source.n238 50.5119
R180 source.n237 source.n236 50.5119
R181 source.n171 source.n170 50.5119
R182 source.n169 source.n168 50.5119
R183 source.n271 source.n270 32.1853
R184 source.n235 source.n234 32.1853
R185 source.n203 source.n202 32.1853
R186 source.n167 source.n166 32.1853
R187 source.n31 source.n30 32.1853
R188 source.n67 source.n66 32.1853
R189 source.n99 source.n98 32.1853
R190 source.n135 source.n134 32.1853
R191 source.n167 source.n135 17.1992
R192 source.n251 source.n249 15.6674
R193 source.n215 source.n213 15.6674
R194 source.n183 source.n181 15.6674
R195 source.n147 source.n145 15.6674
R196 source.n11 source.n9 15.6674
R197 source.n47 source.n45 15.6674
R198 source.n79 source.n77 15.6674
R199 source.n115 source.n113 15.6674
R200 source.n252 source.n248 12.8005
R201 source.n216 source.n212 12.8005
R202 source.n184 source.n180 12.8005
R203 source.n148 source.n144 12.8005
R204 source.n12 source.n8 12.8005
R205 source.n48 source.n44 12.8005
R206 source.n80 source.n76 12.8005
R207 source.n116 source.n112 12.8005
R208 source.n256 source.n255 12.0247
R209 source.n220 source.n219 12.0247
R210 source.n188 source.n187 12.0247
R211 source.n152 source.n151 12.0247
R212 source.n16 source.n15 12.0247
R213 source.n52 source.n51 12.0247
R214 source.n84 source.n83 12.0247
R215 source.n120 source.n119 12.0247
R216 source.n272 source.n31 11.7078
R217 source.n259 source.n246 11.249
R218 source.n223 source.n210 11.249
R219 source.n191 source.n178 11.249
R220 source.n155 source.n142 11.249
R221 source.n19 source.n6 11.249
R222 source.n55 source.n42 11.249
R223 source.n87 source.n74 11.249
R224 source.n123 source.n110 11.249
R225 source.n260 source.n244 10.4732
R226 source.n224 source.n208 10.4732
R227 source.n192 source.n176 10.4732
R228 source.n156 source.n140 10.4732
R229 source.n20 source.n4 10.4732
R230 source.n56 source.n40 10.4732
R231 source.n88 source.n72 10.4732
R232 source.n124 source.n108 10.4732
R233 source.n264 source.n263 9.69747
R234 source.n228 source.n227 9.69747
R235 source.n196 source.n195 9.69747
R236 source.n160 source.n159 9.69747
R237 source.n24 source.n23 9.69747
R238 source.n60 source.n59 9.69747
R239 source.n92 source.n91 9.69747
R240 source.n128 source.n127 9.69747
R241 source.n270 source.n269 9.45567
R242 source.n234 source.n233 9.45567
R243 source.n202 source.n201 9.45567
R244 source.n166 source.n165 9.45567
R245 source.n30 source.n29 9.45567
R246 source.n66 source.n65 9.45567
R247 source.n98 source.n97 9.45567
R248 source.n134 source.n133 9.45567
R249 source.n269 source.n268 9.3005
R250 source.n242 source.n241 9.3005
R251 source.n263 source.n262 9.3005
R252 source.n261 source.n260 9.3005
R253 source.n246 source.n245 9.3005
R254 source.n255 source.n254 9.3005
R255 source.n253 source.n252 9.3005
R256 source.n233 source.n232 9.3005
R257 source.n206 source.n205 9.3005
R258 source.n227 source.n226 9.3005
R259 source.n225 source.n224 9.3005
R260 source.n210 source.n209 9.3005
R261 source.n219 source.n218 9.3005
R262 source.n217 source.n216 9.3005
R263 source.n201 source.n200 9.3005
R264 source.n174 source.n173 9.3005
R265 source.n195 source.n194 9.3005
R266 source.n193 source.n192 9.3005
R267 source.n178 source.n177 9.3005
R268 source.n187 source.n186 9.3005
R269 source.n185 source.n184 9.3005
R270 source.n165 source.n164 9.3005
R271 source.n138 source.n137 9.3005
R272 source.n159 source.n158 9.3005
R273 source.n157 source.n156 9.3005
R274 source.n142 source.n141 9.3005
R275 source.n151 source.n150 9.3005
R276 source.n149 source.n148 9.3005
R277 source.n29 source.n28 9.3005
R278 source.n2 source.n1 9.3005
R279 source.n23 source.n22 9.3005
R280 source.n21 source.n20 9.3005
R281 source.n6 source.n5 9.3005
R282 source.n15 source.n14 9.3005
R283 source.n13 source.n12 9.3005
R284 source.n65 source.n64 9.3005
R285 source.n38 source.n37 9.3005
R286 source.n59 source.n58 9.3005
R287 source.n57 source.n56 9.3005
R288 source.n42 source.n41 9.3005
R289 source.n51 source.n50 9.3005
R290 source.n49 source.n48 9.3005
R291 source.n97 source.n96 9.3005
R292 source.n70 source.n69 9.3005
R293 source.n91 source.n90 9.3005
R294 source.n89 source.n88 9.3005
R295 source.n74 source.n73 9.3005
R296 source.n83 source.n82 9.3005
R297 source.n81 source.n80 9.3005
R298 source.n133 source.n132 9.3005
R299 source.n106 source.n105 9.3005
R300 source.n127 source.n126 9.3005
R301 source.n125 source.n124 9.3005
R302 source.n110 source.n109 9.3005
R303 source.n119 source.n118 9.3005
R304 source.n117 source.n116 9.3005
R305 source.n267 source.n242 8.92171
R306 source.n231 source.n206 8.92171
R307 source.n199 source.n174 8.92171
R308 source.n163 source.n138 8.92171
R309 source.n27 source.n2 8.92171
R310 source.n63 source.n38 8.92171
R311 source.n95 source.n70 8.92171
R312 source.n131 source.n106 8.92171
R313 source.n268 source.n240 8.14595
R314 source.n232 source.n204 8.14595
R315 source.n200 source.n172 8.14595
R316 source.n164 source.n136 8.14595
R317 source.n28 source.n0 8.14595
R318 source.n64 source.n36 8.14595
R319 source.n96 source.n68 8.14595
R320 source.n132 source.n104 8.14595
R321 source.n270 source.n240 5.81868
R322 source.n234 source.n204 5.81868
R323 source.n202 source.n172 5.81868
R324 source.n166 source.n136 5.81868
R325 source.n30 source.n0 5.81868
R326 source.n66 source.n36 5.81868
R327 source.n98 source.n68 5.81868
R328 source.n134 source.n104 5.81868
R329 source.n272 source.n271 5.49188
R330 source.n268 source.n267 5.04292
R331 source.n232 source.n231 5.04292
R332 source.n200 source.n199 5.04292
R333 source.n164 source.n163 5.04292
R334 source.n28 source.n27 5.04292
R335 source.n64 source.n63 5.04292
R336 source.n96 source.n95 5.04292
R337 source.n132 source.n131 5.04292
R338 source.n253 source.n249 4.38594
R339 source.n217 source.n213 4.38594
R340 source.n185 source.n181 4.38594
R341 source.n149 source.n145 4.38594
R342 source.n13 source.n9 4.38594
R343 source.n49 source.n45 4.38594
R344 source.n81 source.n77 4.38594
R345 source.n117 source.n113 4.38594
R346 source.n264 source.n242 4.26717
R347 source.n228 source.n206 4.26717
R348 source.n196 source.n174 4.26717
R349 source.n160 source.n138 4.26717
R350 source.n24 source.n2 4.26717
R351 source.n60 source.n38 4.26717
R352 source.n92 source.n70 4.26717
R353 source.n128 source.n106 4.26717
R354 source.n263 source.n244 3.49141
R355 source.n227 source.n208 3.49141
R356 source.n195 source.n176 3.49141
R357 source.n159 source.n140 3.49141
R358 source.n23 source.n4 3.49141
R359 source.n59 source.n40 3.49141
R360 source.n91 source.n72 3.49141
R361 source.n127 source.n108 3.49141
R362 source.n238 source.t17 3.3005
R363 source.n238 source.t13 3.3005
R364 source.n236 source.t16 3.3005
R365 source.n236 source.t22 3.3005
R366 source.n170 source.t0 3.3005
R367 source.n170 source.t1 3.3005
R368 source.n168 source.t8 3.3005
R369 source.n168 source.t4 3.3005
R370 source.n32 source.t3 3.3005
R371 source.n32 source.t2 3.3005
R372 source.n34 source.t6 3.3005
R373 source.n34 source.t7 3.3005
R374 source.n100 source.t14 3.3005
R375 source.n100 source.t18 3.3005
R376 source.n102 source.t20 3.3005
R377 source.n102 source.t15 3.3005
R378 source.n260 source.n259 2.71565
R379 source.n224 source.n223 2.71565
R380 source.n192 source.n191 2.71565
R381 source.n156 source.n155 2.71565
R382 source.n20 source.n19 2.71565
R383 source.n56 source.n55 2.71565
R384 source.n88 source.n87 2.71565
R385 source.n124 source.n123 2.71565
R386 source.n256 source.n246 1.93989
R387 source.n220 source.n210 1.93989
R388 source.n188 source.n178 1.93989
R389 source.n152 source.n142 1.93989
R390 source.n16 source.n6 1.93989
R391 source.n52 source.n42 1.93989
R392 source.n84 source.n74 1.93989
R393 source.n120 source.n110 1.93989
R394 source.n255 source.n248 1.16414
R395 source.n219 source.n212 1.16414
R396 source.n187 source.n180 1.16414
R397 source.n151 source.n144 1.16414
R398 source.n15 source.n8 1.16414
R399 source.n51 source.n44 1.16414
R400 source.n83 source.n76 1.16414
R401 source.n119 source.n112 1.16414
R402 source.n99 source.n67 0.470328
R403 source.n235 source.n203 0.470328
R404 source.n135 source.n103 0.457397
R405 source.n103 source.n101 0.457397
R406 source.n101 source.n99 0.457397
R407 source.n67 source.n35 0.457397
R408 source.n35 source.n33 0.457397
R409 source.n33 source.n31 0.457397
R410 source.n169 source.n167 0.457397
R411 source.n171 source.n169 0.457397
R412 source.n203 source.n171 0.457397
R413 source.n237 source.n235 0.457397
R414 source.n239 source.n237 0.457397
R415 source.n271 source.n239 0.457397
R416 source.n252 source.n251 0.388379
R417 source.n216 source.n215 0.388379
R418 source.n184 source.n183 0.388379
R419 source.n148 source.n147 0.388379
R420 source.n12 source.n11 0.388379
R421 source.n48 source.n47 0.388379
R422 source.n80 source.n79 0.388379
R423 source.n116 source.n115 0.388379
R424 source source.n272 0.188
R425 source.n254 source.n253 0.155672
R426 source.n254 source.n245 0.155672
R427 source.n261 source.n245 0.155672
R428 source.n262 source.n261 0.155672
R429 source.n262 source.n241 0.155672
R430 source.n269 source.n241 0.155672
R431 source.n218 source.n217 0.155672
R432 source.n218 source.n209 0.155672
R433 source.n225 source.n209 0.155672
R434 source.n226 source.n225 0.155672
R435 source.n226 source.n205 0.155672
R436 source.n233 source.n205 0.155672
R437 source.n186 source.n185 0.155672
R438 source.n186 source.n177 0.155672
R439 source.n193 source.n177 0.155672
R440 source.n194 source.n193 0.155672
R441 source.n194 source.n173 0.155672
R442 source.n201 source.n173 0.155672
R443 source.n150 source.n149 0.155672
R444 source.n150 source.n141 0.155672
R445 source.n157 source.n141 0.155672
R446 source.n158 source.n157 0.155672
R447 source.n158 source.n137 0.155672
R448 source.n165 source.n137 0.155672
R449 source.n29 source.n1 0.155672
R450 source.n22 source.n1 0.155672
R451 source.n22 source.n21 0.155672
R452 source.n21 source.n5 0.155672
R453 source.n14 source.n5 0.155672
R454 source.n14 source.n13 0.155672
R455 source.n65 source.n37 0.155672
R456 source.n58 source.n37 0.155672
R457 source.n58 source.n57 0.155672
R458 source.n57 source.n41 0.155672
R459 source.n50 source.n41 0.155672
R460 source.n50 source.n49 0.155672
R461 source.n97 source.n69 0.155672
R462 source.n90 source.n69 0.155672
R463 source.n90 source.n89 0.155672
R464 source.n89 source.n73 0.155672
R465 source.n82 source.n73 0.155672
R466 source.n82 source.n81 0.155672
R467 source.n133 source.n105 0.155672
R468 source.n126 source.n105 0.155672
R469 source.n126 source.n125 0.155672
R470 source.n125 source.n109 0.155672
R471 source.n118 source.n109 0.155672
R472 source.n118 source.n117 0.155672
R473 drain_right.n6 drain_right.n4 67.6476
R474 drain_right.n3 drain_right.n2 67.5922
R475 drain_right.n3 drain_right.n0 67.5922
R476 drain_right.n6 drain_right.n5 67.1908
R477 drain_right.n8 drain_right.n7 67.1908
R478 drain_right.n3 drain_right.n1 67.1907
R479 drain_right drain_right.n3 24.5529
R480 drain_right drain_right.n8 6.11011
R481 drain_right.n1 drain_right.t5 3.3005
R482 drain_right.n1 drain_right.t2 3.3005
R483 drain_right.n2 drain_right.t10 3.3005
R484 drain_right.n2 drain_right.t0 3.3005
R485 drain_right.n0 drain_right.t4 3.3005
R486 drain_right.n0 drain_right.t1 3.3005
R487 drain_right.n4 drain_right.t8 3.3005
R488 drain_right.n4 drain_right.t7 3.3005
R489 drain_right.n5 drain_right.t3 3.3005
R490 drain_right.n5 drain_right.t11 3.3005
R491 drain_right.n7 drain_right.t9 3.3005
R492 drain_right.n7 drain_right.t6 3.3005
R493 drain_right.n8 drain_right.n6 0.457397
R494 plus.n2 plus.t4 927.12
R495 plus.n11 plus.t3 927.12
R496 plus.n15 plus.t7 927.12
R497 plus.n24 plus.t1 927.12
R498 plus.n3 plus.t0 879.65
R499 plus.n1 plus.t11 879.65
R500 plus.n8 plus.t10 879.65
R501 plus.n10 plus.t9 879.65
R502 plus.n16 plus.t8 879.65
R503 plus.n14 plus.t5 879.65
R504 plus.n21 plus.t2 879.65
R505 plus.n23 plus.t6 879.65
R506 plus.n5 plus.n2 161.489
R507 plus.n18 plus.n15 161.489
R508 plus.n5 plus.n4 161.3
R509 plus.n7 plus.n6 161.3
R510 plus.n9 plus.n0 161.3
R511 plus.n12 plus.n11 161.3
R512 plus.n18 plus.n17 161.3
R513 plus.n20 plus.n19 161.3
R514 plus.n22 plus.n13 161.3
R515 plus.n25 plus.n24 161.3
R516 plus.n4 plus.n3 43.0884
R517 plus.n10 plus.n9 43.0884
R518 plus.n23 plus.n22 43.0884
R519 plus.n17 plus.n16 43.0884
R520 plus.n7 plus.n1 38.7066
R521 plus.n8 plus.n7 38.7066
R522 plus.n21 plus.n20 38.7066
R523 plus.n20 plus.n14 38.7066
R524 plus.n4 plus.n1 34.3247
R525 plus.n9 plus.n8 34.3247
R526 plus.n22 plus.n21 34.3247
R527 plus.n17 plus.n14 34.3247
R528 plus.n3 plus.n2 29.9429
R529 plus.n11 plus.n10 29.9429
R530 plus.n24 plus.n23 29.9429
R531 plus.n16 plus.n15 29.9429
R532 plus plus.n25 26.2074
R533 plus plus.n12 9.82626
R534 plus.n6 plus.n5 0.189894
R535 plus.n6 plus.n0 0.189894
R536 plus.n12 plus.n0 0.189894
R537 plus.n25 plus.n13 0.189894
R538 plus.n19 plus.n13 0.189894
R539 plus.n19 plus.n18 0.189894
R540 drain_left.n6 drain_left.n4 67.6477
R541 drain_left.n3 drain_left.n2 67.5922
R542 drain_left.n3 drain_left.n0 67.5922
R543 drain_left.n6 drain_left.n5 67.1908
R544 drain_left.n8 drain_left.n7 67.1907
R545 drain_left.n3 drain_left.n1 67.1907
R546 drain_left drain_left.n3 25.1061
R547 drain_left drain_left.n8 6.11011
R548 drain_left.n1 drain_left.t9 3.3005
R549 drain_left.n1 drain_left.t6 3.3005
R550 drain_left.n2 drain_left.t3 3.3005
R551 drain_left.n2 drain_left.t4 3.3005
R552 drain_left.n0 drain_left.t10 3.3005
R553 drain_left.n0 drain_left.t5 3.3005
R554 drain_left.n7 drain_left.t2 3.3005
R555 drain_left.n7 drain_left.t8 3.3005
R556 drain_left.n5 drain_left.t0 3.3005
R557 drain_left.n5 drain_left.t1 3.3005
R558 drain_left.n4 drain_left.t7 3.3005
R559 drain_left.n4 drain_left.t11 3.3005
R560 drain_left.n8 drain_left.n6 0.457397
C0 plus source 1.8446f
C1 plus drain_left 2.11597f
C2 drain_right minus 1.97709f
C3 drain_right source 15.1989f
C4 minus source 1.83058f
C5 drain_right drain_left 0.711832f
C6 drain_left minus 0.17046f
C7 drain_left source 15.1998f
C8 drain_right plus 0.292203f
C9 plus minus 3.86167f
C10 drain_right a_n1458_n2088# 4.60082f
C11 drain_left a_n1458_n2088# 5.12728f
C12 source a_n1458_n2088# 5.13588f
C13 minus a_n1458_n2088# 5.154593f
C14 plus a_n1458_n2088# 6.37513f
C15 drain_left.t10 a_n1458_n2088# 0.174685f
C16 drain_left.t5 a_n1458_n2088# 0.174685f
C17 drain_left.n0 a_n1458_n2088# 1.45936f
C18 drain_left.t9 a_n1458_n2088# 0.174685f
C19 drain_left.t6 a_n1458_n2088# 0.174685f
C20 drain_left.n1 a_n1458_n2088# 1.45688f
C21 drain_left.t3 a_n1458_n2088# 0.174685f
C22 drain_left.t4 a_n1458_n2088# 0.174685f
C23 drain_left.n2 a_n1458_n2088# 1.45936f
C24 drain_left.n3 a_n1458_n2088# 2.35862f
C25 drain_left.t7 a_n1458_n2088# 0.174685f
C26 drain_left.t11 a_n1458_n2088# 0.174685f
C27 drain_left.n4 a_n1458_n2088# 1.45974f
C28 drain_left.t0 a_n1458_n2088# 0.174685f
C29 drain_left.t1 a_n1458_n2088# 0.174685f
C30 drain_left.n5 a_n1458_n2088# 1.45688f
C31 drain_left.n6 a_n1458_n2088# 0.826993f
C32 drain_left.t2 a_n1458_n2088# 0.174685f
C33 drain_left.t8 a_n1458_n2088# 0.174685f
C34 drain_left.n7 a_n1458_n2088# 1.45688f
C35 drain_left.n8 a_n1458_n2088# 0.709033f
C36 plus.n0 a_n1458_n2088# 0.043989f
C37 plus.t9 a_n1458_n2088# 0.1504f
C38 plus.t10 a_n1458_n2088# 0.1504f
C39 plus.t11 a_n1458_n2088# 0.1504f
C40 plus.n1 a_n1458_n2088# 0.073556f
C41 plus.t4 a_n1458_n2088# 0.154201f
C42 plus.n2 a_n1458_n2088# 0.085902f
C43 plus.t0 a_n1458_n2088# 0.1504f
C44 plus.n3 a_n1458_n2088# 0.073556f
C45 plus.n4 a_n1458_n2088# 0.015406f
C46 plus.n5 a_n1458_n2088# 0.097408f
C47 plus.n6 a_n1458_n2088# 0.043989f
C48 plus.n7 a_n1458_n2088# 0.015406f
C49 plus.n8 a_n1458_n2088# 0.073556f
C50 plus.n9 a_n1458_n2088# 0.015406f
C51 plus.n10 a_n1458_n2088# 0.073556f
C52 plus.t3 a_n1458_n2088# 0.154201f
C53 plus.n11 a_n1458_n2088# 0.08584f
C54 plus.n12 a_n1458_n2088# 0.372075f
C55 plus.n13 a_n1458_n2088# 0.043989f
C56 plus.t1 a_n1458_n2088# 0.154201f
C57 plus.t6 a_n1458_n2088# 0.1504f
C58 plus.t2 a_n1458_n2088# 0.1504f
C59 plus.t5 a_n1458_n2088# 0.1504f
C60 plus.n14 a_n1458_n2088# 0.073556f
C61 plus.t7 a_n1458_n2088# 0.154201f
C62 plus.n15 a_n1458_n2088# 0.085902f
C63 plus.t8 a_n1458_n2088# 0.1504f
C64 plus.n16 a_n1458_n2088# 0.073556f
C65 plus.n17 a_n1458_n2088# 0.015406f
C66 plus.n18 a_n1458_n2088# 0.097408f
C67 plus.n19 a_n1458_n2088# 0.043989f
C68 plus.n20 a_n1458_n2088# 0.015406f
C69 plus.n21 a_n1458_n2088# 0.073556f
C70 plus.n22 a_n1458_n2088# 0.015406f
C71 plus.n23 a_n1458_n2088# 0.073556f
C72 plus.n24 a_n1458_n2088# 0.08584f
C73 plus.n25 a_n1458_n2088# 1.0355f
C74 drain_right.t4 a_n1458_n2088# 0.15477f
C75 drain_right.t1 a_n1458_n2088# 0.15477f
C76 drain_right.n0 a_n1458_n2088# 1.29298f
C77 drain_right.t5 a_n1458_n2088# 0.15477f
C78 drain_right.t2 a_n1458_n2088# 0.15477f
C79 drain_right.n1 a_n1458_n2088# 1.29078f
C80 drain_right.t10 a_n1458_n2088# 0.15477f
C81 drain_right.t0 a_n1458_n2088# 0.15477f
C82 drain_right.n2 a_n1458_n2088# 1.29298f
C83 drain_right.n3 a_n1458_n2088# 2.02303f
C84 drain_right.t8 a_n1458_n2088# 0.15477f
C85 drain_right.t7 a_n1458_n2088# 0.15477f
C86 drain_right.n4 a_n1458_n2088# 1.29331f
C87 drain_right.t3 a_n1458_n2088# 0.15477f
C88 drain_right.t11 a_n1458_n2088# 0.15477f
C89 drain_right.n5 a_n1458_n2088# 1.29079f
C90 drain_right.n6 a_n1458_n2088# 0.732717f
C91 drain_right.t9 a_n1458_n2088# 0.15477f
C92 drain_right.t6 a_n1458_n2088# 0.15477f
C93 drain_right.n7 a_n1458_n2088# 1.29079f
C94 drain_right.n8 a_n1458_n2088# 0.628193f
C95 source.n0 a_n1458_n2088# 0.038819f
C96 source.n1 a_n1458_n2088# 0.027617f
C97 source.n2 a_n1458_n2088# 0.01484f
C98 source.n3 a_n1458_n2088# 0.035077f
C99 source.n4 a_n1458_n2088# 0.015713f
C100 source.n5 a_n1458_n2088# 0.027617f
C101 source.n6 a_n1458_n2088# 0.01484f
C102 source.n7 a_n1458_n2088# 0.035077f
C103 source.n8 a_n1458_n2088# 0.015713f
C104 source.n9 a_n1458_n2088# 0.118183f
C105 source.t5 a_n1458_n2088# 0.057171f
C106 source.n10 a_n1458_n2088# 0.026308f
C107 source.n11 a_n1458_n2088# 0.02072f
C108 source.n12 a_n1458_n2088# 0.01484f
C109 source.n13 a_n1458_n2088# 0.657129f
C110 source.n14 a_n1458_n2088# 0.027617f
C111 source.n15 a_n1458_n2088# 0.01484f
C112 source.n16 a_n1458_n2088# 0.015713f
C113 source.n17 a_n1458_n2088# 0.035077f
C114 source.n18 a_n1458_n2088# 0.035077f
C115 source.n19 a_n1458_n2088# 0.015713f
C116 source.n20 a_n1458_n2088# 0.01484f
C117 source.n21 a_n1458_n2088# 0.027617f
C118 source.n22 a_n1458_n2088# 0.027617f
C119 source.n23 a_n1458_n2088# 0.01484f
C120 source.n24 a_n1458_n2088# 0.015713f
C121 source.n25 a_n1458_n2088# 0.035077f
C122 source.n26 a_n1458_n2088# 0.075936f
C123 source.n27 a_n1458_n2088# 0.015713f
C124 source.n28 a_n1458_n2088# 0.01484f
C125 source.n29 a_n1458_n2088# 0.063836f
C126 source.n30 a_n1458_n2088# 0.042489f
C127 source.n31 a_n1458_n2088# 0.65579f
C128 source.t3 a_n1458_n2088# 0.130945f
C129 source.t2 a_n1458_n2088# 0.130945f
C130 source.n32 a_n1458_n2088# 1.01981f
C131 source.n33 a_n1458_n2088# 0.340205f
C132 source.t6 a_n1458_n2088# 0.130945f
C133 source.t7 a_n1458_n2088# 0.130945f
C134 source.n34 a_n1458_n2088# 1.01981f
C135 source.n35 a_n1458_n2088# 0.340205f
C136 source.n36 a_n1458_n2088# 0.038819f
C137 source.n37 a_n1458_n2088# 0.027617f
C138 source.n38 a_n1458_n2088# 0.01484f
C139 source.n39 a_n1458_n2088# 0.035077f
C140 source.n40 a_n1458_n2088# 0.015713f
C141 source.n41 a_n1458_n2088# 0.027617f
C142 source.n42 a_n1458_n2088# 0.01484f
C143 source.n43 a_n1458_n2088# 0.035077f
C144 source.n44 a_n1458_n2088# 0.015713f
C145 source.n45 a_n1458_n2088# 0.118183f
C146 source.t9 a_n1458_n2088# 0.057171f
C147 source.n46 a_n1458_n2088# 0.026308f
C148 source.n47 a_n1458_n2088# 0.02072f
C149 source.n48 a_n1458_n2088# 0.01484f
C150 source.n49 a_n1458_n2088# 0.657129f
C151 source.n50 a_n1458_n2088# 0.027617f
C152 source.n51 a_n1458_n2088# 0.01484f
C153 source.n52 a_n1458_n2088# 0.015713f
C154 source.n53 a_n1458_n2088# 0.035077f
C155 source.n54 a_n1458_n2088# 0.035077f
C156 source.n55 a_n1458_n2088# 0.015713f
C157 source.n56 a_n1458_n2088# 0.01484f
C158 source.n57 a_n1458_n2088# 0.027617f
C159 source.n58 a_n1458_n2088# 0.027617f
C160 source.n59 a_n1458_n2088# 0.01484f
C161 source.n60 a_n1458_n2088# 0.015713f
C162 source.n61 a_n1458_n2088# 0.035077f
C163 source.n62 a_n1458_n2088# 0.075936f
C164 source.n63 a_n1458_n2088# 0.015713f
C165 source.n64 a_n1458_n2088# 0.01484f
C166 source.n65 a_n1458_n2088# 0.063836f
C167 source.n66 a_n1458_n2088# 0.042489f
C168 source.n67 a_n1458_n2088# 0.106056f
C169 source.n68 a_n1458_n2088# 0.038819f
C170 source.n69 a_n1458_n2088# 0.027617f
C171 source.n70 a_n1458_n2088# 0.01484f
C172 source.n71 a_n1458_n2088# 0.035077f
C173 source.n72 a_n1458_n2088# 0.015713f
C174 source.n73 a_n1458_n2088# 0.027617f
C175 source.n74 a_n1458_n2088# 0.01484f
C176 source.n75 a_n1458_n2088# 0.035077f
C177 source.n76 a_n1458_n2088# 0.015713f
C178 source.n77 a_n1458_n2088# 0.118183f
C179 source.t21 a_n1458_n2088# 0.057171f
C180 source.n78 a_n1458_n2088# 0.026308f
C181 source.n79 a_n1458_n2088# 0.02072f
C182 source.n80 a_n1458_n2088# 0.01484f
C183 source.n81 a_n1458_n2088# 0.657129f
C184 source.n82 a_n1458_n2088# 0.027617f
C185 source.n83 a_n1458_n2088# 0.01484f
C186 source.n84 a_n1458_n2088# 0.015713f
C187 source.n85 a_n1458_n2088# 0.035077f
C188 source.n86 a_n1458_n2088# 0.035077f
C189 source.n87 a_n1458_n2088# 0.015713f
C190 source.n88 a_n1458_n2088# 0.01484f
C191 source.n89 a_n1458_n2088# 0.027617f
C192 source.n90 a_n1458_n2088# 0.027617f
C193 source.n91 a_n1458_n2088# 0.01484f
C194 source.n92 a_n1458_n2088# 0.015713f
C195 source.n93 a_n1458_n2088# 0.035077f
C196 source.n94 a_n1458_n2088# 0.075936f
C197 source.n95 a_n1458_n2088# 0.015713f
C198 source.n96 a_n1458_n2088# 0.01484f
C199 source.n97 a_n1458_n2088# 0.063836f
C200 source.n98 a_n1458_n2088# 0.042489f
C201 source.n99 a_n1458_n2088# 0.106056f
C202 source.t14 a_n1458_n2088# 0.130945f
C203 source.t18 a_n1458_n2088# 0.130945f
C204 source.n100 a_n1458_n2088# 1.01981f
C205 source.n101 a_n1458_n2088# 0.340205f
C206 source.t20 a_n1458_n2088# 0.130945f
C207 source.t15 a_n1458_n2088# 0.130945f
C208 source.n102 a_n1458_n2088# 1.01981f
C209 source.n103 a_n1458_n2088# 0.340205f
C210 source.n104 a_n1458_n2088# 0.038819f
C211 source.n105 a_n1458_n2088# 0.027617f
C212 source.n106 a_n1458_n2088# 0.01484f
C213 source.n107 a_n1458_n2088# 0.035077f
C214 source.n108 a_n1458_n2088# 0.015713f
C215 source.n109 a_n1458_n2088# 0.027617f
C216 source.n110 a_n1458_n2088# 0.01484f
C217 source.n111 a_n1458_n2088# 0.035077f
C218 source.n112 a_n1458_n2088# 0.015713f
C219 source.n113 a_n1458_n2088# 0.118183f
C220 source.t12 a_n1458_n2088# 0.057171f
C221 source.n114 a_n1458_n2088# 0.026308f
C222 source.n115 a_n1458_n2088# 0.02072f
C223 source.n116 a_n1458_n2088# 0.01484f
C224 source.n117 a_n1458_n2088# 0.657129f
C225 source.n118 a_n1458_n2088# 0.027617f
C226 source.n119 a_n1458_n2088# 0.01484f
C227 source.n120 a_n1458_n2088# 0.015713f
C228 source.n121 a_n1458_n2088# 0.035077f
C229 source.n122 a_n1458_n2088# 0.035077f
C230 source.n123 a_n1458_n2088# 0.015713f
C231 source.n124 a_n1458_n2088# 0.01484f
C232 source.n125 a_n1458_n2088# 0.027617f
C233 source.n126 a_n1458_n2088# 0.027617f
C234 source.n127 a_n1458_n2088# 0.01484f
C235 source.n128 a_n1458_n2088# 0.015713f
C236 source.n129 a_n1458_n2088# 0.035077f
C237 source.n130 a_n1458_n2088# 0.075936f
C238 source.n131 a_n1458_n2088# 0.015713f
C239 source.n132 a_n1458_n2088# 0.01484f
C240 source.n133 a_n1458_n2088# 0.063836f
C241 source.n134 a_n1458_n2088# 0.042489f
C242 source.n135 a_n1458_n2088# 1.00915f
C243 source.n136 a_n1458_n2088# 0.038819f
C244 source.n137 a_n1458_n2088# 0.027617f
C245 source.n138 a_n1458_n2088# 0.01484f
C246 source.n139 a_n1458_n2088# 0.035077f
C247 source.n140 a_n1458_n2088# 0.015713f
C248 source.n141 a_n1458_n2088# 0.027617f
C249 source.n142 a_n1458_n2088# 0.01484f
C250 source.n143 a_n1458_n2088# 0.035077f
C251 source.n144 a_n1458_n2088# 0.015713f
C252 source.n145 a_n1458_n2088# 0.118183f
C253 source.t10 a_n1458_n2088# 0.057171f
C254 source.n146 a_n1458_n2088# 0.026308f
C255 source.n147 a_n1458_n2088# 0.02072f
C256 source.n148 a_n1458_n2088# 0.01484f
C257 source.n149 a_n1458_n2088# 0.657129f
C258 source.n150 a_n1458_n2088# 0.027617f
C259 source.n151 a_n1458_n2088# 0.01484f
C260 source.n152 a_n1458_n2088# 0.015713f
C261 source.n153 a_n1458_n2088# 0.035077f
C262 source.n154 a_n1458_n2088# 0.035077f
C263 source.n155 a_n1458_n2088# 0.015713f
C264 source.n156 a_n1458_n2088# 0.01484f
C265 source.n157 a_n1458_n2088# 0.027617f
C266 source.n158 a_n1458_n2088# 0.027617f
C267 source.n159 a_n1458_n2088# 0.01484f
C268 source.n160 a_n1458_n2088# 0.015713f
C269 source.n161 a_n1458_n2088# 0.035077f
C270 source.n162 a_n1458_n2088# 0.075936f
C271 source.n163 a_n1458_n2088# 0.015713f
C272 source.n164 a_n1458_n2088# 0.01484f
C273 source.n165 a_n1458_n2088# 0.063836f
C274 source.n166 a_n1458_n2088# 0.042489f
C275 source.n167 a_n1458_n2088# 1.00915f
C276 source.t8 a_n1458_n2088# 0.130945f
C277 source.t4 a_n1458_n2088# 0.130945f
C278 source.n168 a_n1458_n2088# 1.0198f
C279 source.n169 a_n1458_n2088# 0.340212f
C280 source.t0 a_n1458_n2088# 0.130945f
C281 source.t1 a_n1458_n2088# 0.130945f
C282 source.n170 a_n1458_n2088# 1.0198f
C283 source.n171 a_n1458_n2088# 0.340212f
C284 source.n172 a_n1458_n2088# 0.038819f
C285 source.n173 a_n1458_n2088# 0.027617f
C286 source.n174 a_n1458_n2088# 0.01484f
C287 source.n175 a_n1458_n2088# 0.035077f
C288 source.n176 a_n1458_n2088# 0.015713f
C289 source.n177 a_n1458_n2088# 0.027617f
C290 source.n178 a_n1458_n2088# 0.01484f
C291 source.n179 a_n1458_n2088# 0.035077f
C292 source.n180 a_n1458_n2088# 0.015713f
C293 source.n181 a_n1458_n2088# 0.118183f
C294 source.t11 a_n1458_n2088# 0.057171f
C295 source.n182 a_n1458_n2088# 0.026308f
C296 source.n183 a_n1458_n2088# 0.02072f
C297 source.n184 a_n1458_n2088# 0.01484f
C298 source.n185 a_n1458_n2088# 0.657129f
C299 source.n186 a_n1458_n2088# 0.027617f
C300 source.n187 a_n1458_n2088# 0.01484f
C301 source.n188 a_n1458_n2088# 0.015713f
C302 source.n189 a_n1458_n2088# 0.035077f
C303 source.n190 a_n1458_n2088# 0.035077f
C304 source.n191 a_n1458_n2088# 0.015713f
C305 source.n192 a_n1458_n2088# 0.01484f
C306 source.n193 a_n1458_n2088# 0.027617f
C307 source.n194 a_n1458_n2088# 0.027617f
C308 source.n195 a_n1458_n2088# 0.01484f
C309 source.n196 a_n1458_n2088# 0.015713f
C310 source.n197 a_n1458_n2088# 0.035077f
C311 source.n198 a_n1458_n2088# 0.075936f
C312 source.n199 a_n1458_n2088# 0.015713f
C313 source.n200 a_n1458_n2088# 0.01484f
C314 source.n201 a_n1458_n2088# 0.063836f
C315 source.n202 a_n1458_n2088# 0.042489f
C316 source.n203 a_n1458_n2088# 0.106056f
C317 source.n204 a_n1458_n2088# 0.038819f
C318 source.n205 a_n1458_n2088# 0.027617f
C319 source.n206 a_n1458_n2088# 0.01484f
C320 source.n207 a_n1458_n2088# 0.035077f
C321 source.n208 a_n1458_n2088# 0.015713f
C322 source.n209 a_n1458_n2088# 0.027617f
C323 source.n210 a_n1458_n2088# 0.01484f
C324 source.n211 a_n1458_n2088# 0.035077f
C325 source.n212 a_n1458_n2088# 0.015713f
C326 source.n213 a_n1458_n2088# 0.118183f
C327 source.t19 a_n1458_n2088# 0.057171f
C328 source.n214 a_n1458_n2088# 0.026308f
C329 source.n215 a_n1458_n2088# 0.02072f
C330 source.n216 a_n1458_n2088# 0.01484f
C331 source.n217 a_n1458_n2088# 0.657129f
C332 source.n218 a_n1458_n2088# 0.027617f
C333 source.n219 a_n1458_n2088# 0.01484f
C334 source.n220 a_n1458_n2088# 0.015713f
C335 source.n221 a_n1458_n2088# 0.035077f
C336 source.n222 a_n1458_n2088# 0.035077f
C337 source.n223 a_n1458_n2088# 0.015713f
C338 source.n224 a_n1458_n2088# 0.01484f
C339 source.n225 a_n1458_n2088# 0.027617f
C340 source.n226 a_n1458_n2088# 0.027617f
C341 source.n227 a_n1458_n2088# 0.01484f
C342 source.n228 a_n1458_n2088# 0.015713f
C343 source.n229 a_n1458_n2088# 0.035077f
C344 source.n230 a_n1458_n2088# 0.075936f
C345 source.n231 a_n1458_n2088# 0.015713f
C346 source.n232 a_n1458_n2088# 0.01484f
C347 source.n233 a_n1458_n2088# 0.063836f
C348 source.n234 a_n1458_n2088# 0.042489f
C349 source.n235 a_n1458_n2088# 0.106056f
C350 source.t16 a_n1458_n2088# 0.130945f
C351 source.t22 a_n1458_n2088# 0.130945f
C352 source.n236 a_n1458_n2088# 1.0198f
C353 source.n237 a_n1458_n2088# 0.340212f
C354 source.t17 a_n1458_n2088# 0.130945f
C355 source.t13 a_n1458_n2088# 0.130945f
C356 source.n238 a_n1458_n2088# 1.0198f
C357 source.n239 a_n1458_n2088# 0.340212f
C358 source.n240 a_n1458_n2088# 0.038819f
C359 source.n241 a_n1458_n2088# 0.027617f
C360 source.n242 a_n1458_n2088# 0.01484f
C361 source.n243 a_n1458_n2088# 0.035077f
C362 source.n244 a_n1458_n2088# 0.015713f
C363 source.n245 a_n1458_n2088# 0.027617f
C364 source.n246 a_n1458_n2088# 0.01484f
C365 source.n247 a_n1458_n2088# 0.035077f
C366 source.n248 a_n1458_n2088# 0.015713f
C367 source.n249 a_n1458_n2088# 0.118183f
C368 source.t23 a_n1458_n2088# 0.057171f
C369 source.n250 a_n1458_n2088# 0.026308f
C370 source.n251 a_n1458_n2088# 0.02072f
C371 source.n252 a_n1458_n2088# 0.01484f
C372 source.n253 a_n1458_n2088# 0.657129f
C373 source.n254 a_n1458_n2088# 0.027617f
C374 source.n255 a_n1458_n2088# 0.01484f
C375 source.n256 a_n1458_n2088# 0.015713f
C376 source.n257 a_n1458_n2088# 0.035077f
C377 source.n258 a_n1458_n2088# 0.035077f
C378 source.n259 a_n1458_n2088# 0.015713f
C379 source.n260 a_n1458_n2088# 0.01484f
C380 source.n261 a_n1458_n2088# 0.027617f
C381 source.n262 a_n1458_n2088# 0.027617f
C382 source.n263 a_n1458_n2088# 0.01484f
C383 source.n264 a_n1458_n2088# 0.015713f
C384 source.n265 a_n1458_n2088# 0.035077f
C385 source.n266 a_n1458_n2088# 0.075936f
C386 source.n267 a_n1458_n2088# 0.015713f
C387 source.n268 a_n1458_n2088# 0.01484f
C388 source.n269 a_n1458_n2088# 0.063836f
C389 source.n270 a_n1458_n2088# 0.042489f
C390 source.n271 a_n1458_n2088# 0.255806f
C391 source.n272 a_n1458_n2088# 1.12635f
C392 minus.n0 a_n1458_n2088# 0.028175f
C393 minus.t2 a_n1458_n2088# 0.098766f
C394 minus.t5 a_n1458_n2088# 0.096332f
C395 minus.t8 a_n1458_n2088# 0.096332f
C396 minus.t0 a_n1458_n2088# 0.096332f
C397 minus.n1 a_n1458_n2088# 0.047113f
C398 minus.t4 a_n1458_n2088# 0.098766f
C399 minus.n2 a_n1458_n2088# 0.055021f
C400 minus.t3 a_n1458_n2088# 0.096332f
C401 minus.n3 a_n1458_n2088# 0.047113f
C402 minus.n4 a_n1458_n2088# 0.009868f
C403 minus.n5 a_n1458_n2088# 0.06239f
C404 minus.n6 a_n1458_n2088# 0.028175f
C405 minus.n7 a_n1458_n2088# 0.009868f
C406 minus.n8 a_n1458_n2088# 0.047113f
C407 minus.n9 a_n1458_n2088# 0.009868f
C408 minus.n10 a_n1458_n2088# 0.047113f
C409 minus.n11 a_n1458_n2088# 0.054981f
C410 minus.n12 a_n1458_n2088# 0.734015f
C411 minus.n13 a_n1458_n2088# 0.028175f
C412 minus.t1 a_n1458_n2088# 0.096332f
C413 minus.t9 a_n1458_n2088# 0.096332f
C414 minus.t6 a_n1458_n2088# 0.096332f
C415 minus.n14 a_n1458_n2088# 0.047113f
C416 minus.t7 a_n1458_n2088# 0.098766f
C417 minus.n15 a_n1458_n2088# 0.055021f
C418 minus.t10 a_n1458_n2088# 0.096332f
C419 minus.n16 a_n1458_n2088# 0.047113f
C420 minus.n17 a_n1458_n2088# 0.009868f
C421 minus.n18 a_n1458_n2088# 0.06239f
C422 minus.n19 a_n1458_n2088# 0.028175f
C423 minus.n20 a_n1458_n2088# 0.009868f
C424 minus.n21 a_n1458_n2088# 0.047113f
C425 minus.n22 a_n1458_n2088# 0.009868f
C426 minus.n23 a_n1458_n2088# 0.047113f
C427 minus.t11 a_n1458_n2088# 0.098766f
C428 minus.n24 a_n1458_n2088# 0.054981f
C429 minus.n25 a_n1458_n2088# 0.181212f
C430 minus.n26 a_n1458_n2088# 0.906957f
.ends

