* NGSPICE file created from diffpair305.ext - technology: sky130A

.subckt diffpair305 minus drain_right drain_left source plus
X0 source.t20 plus.t0 drain_left.t5 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X1 source.t19 plus.t1 drain_left.t4 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X2 source.t23 minus.t0 drain_right.t11 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X3 drain_left.t3 plus.t2 source.t18 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X4 source.t17 plus.t3 drain_left.t2 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X5 source.t16 plus.t4 drain_left.t10 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X6 drain_left.t6 plus.t5 source.t15 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X7 a_n2158_n2088# a_n2158_n2088# a_n2158_n2088# a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.7
X8 drain_right.t10 minus.t1 source.t1 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X9 drain_right.t9 minus.t2 source.t0 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X10 drain_left.t1 plus.t6 source.t14 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X11 drain_right.t8 minus.t3 source.t21 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X12 source.t22 minus.t4 drain_right.t7 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X13 source.t13 plus.t7 drain_left.t7 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X14 drain_left.t8 plus.t8 source.t12 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X15 drain_right.t6 minus.t5 source.t2 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X16 drain_left.t9 plus.t9 source.t11 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X17 a_n2158_n2088# a_n2158_n2088# a_n2158_n2088# a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X18 drain_right.t5 minus.t6 source.t6 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X19 source.t7 minus.t7 drain_right.t4 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X20 a_n2158_n2088# a_n2158_n2088# a_n2158_n2088# a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X21 drain_left.t0 plus.t10 source.t10 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X22 source.t9 plus.t11 drain_left.t11 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X23 source.t4 minus.t8 drain_right.t3 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X24 drain_right.t2 minus.t9 source.t5 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X25 source.t8 minus.t10 drain_right.t1 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X26 source.t3 minus.t11 drain_right.t0 a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X27 a_n2158_n2088# a_n2158_n2088# a_n2158_n2088# a_n2158_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
R0 plus.n5 plus.t4 285.995
R1 plus.n23 plus.t6 285.995
R2 plus.n16 plus.t9 262.69
R3 plus.n14 plus.t3 262.69
R4 plus.n2 plus.t8 262.69
R5 plus.n8 plus.t1 262.69
R6 plus.n4 plus.t10 262.69
R7 plus.n34 plus.t11 262.69
R8 plus.n32 plus.t2 262.69
R9 plus.n20 plus.t0 262.69
R10 plus.n26 plus.t5 262.69
R11 plus.n22 plus.t7 262.69
R12 plus.n7 plus.n6 161.3
R13 plus.n8 plus.n3 161.3
R14 plus.n10 plus.n9 161.3
R15 plus.n11 plus.n2 161.3
R16 plus.n13 plus.n12 161.3
R17 plus.n14 plus.n1 161.3
R18 plus.n15 plus.n0 161.3
R19 plus.n17 plus.n16 161.3
R20 plus.n25 plus.n24 161.3
R21 plus.n26 plus.n21 161.3
R22 plus.n28 plus.n27 161.3
R23 plus.n29 plus.n20 161.3
R24 plus.n31 plus.n30 161.3
R25 plus.n32 plus.n19 161.3
R26 plus.n33 plus.n18 161.3
R27 plus.n35 plus.n34 161.3
R28 plus.n6 plus.n5 44.8907
R29 plus.n24 plus.n23 44.8907
R30 plus.n16 plus.n15 32.8641
R31 plus.n34 plus.n33 32.8641
R32 plus plus.n35 29.0483
R33 plus.n14 plus.n13 28.4823
R34 plus.n7 plus.n4 28.4823
R35 plus.n32 plus.n31 28.4823
R36 plus.n25 plus.n22 28.4823
R37 plus.n9 plus.n8 24.1005
R38 plus.n9 plus.n2 24.1005
R39 plus.n27 plus.n20 24.1005
R40 plus.n27 plus.n26 24.1005
R41 plus.n13 plus.n2 19.7187
R42 plus.n8 plus.n7 19.7187
R43 plus.n31 plus.n20 19.7187
R44 plus.n26 plus.n25 19.7187
R45 plus.n5 plus.n4 18.4104
R46 plus.n23 plus.n22 18.4104
R47 plus.n15 plus.n14 15.3369
R48 plus.n33 plus.n32 15.3369
R49 plus plus.n17 10.0157
R50 plus.n6 plus.n3 0.189894
R51 plus.n10 plus.n3 0.189894
R52 plus.n11 plus.n10 0.189894
R53 plus.n12 plus.n11 0.189894
R54 plus.n12 plus.n1 0.189894
R55 plus.n1 plus.n0 0.189894
R56 plus.n17 plus.n0 0.189894
R57 plus.n35 plus.n18 0.189894
R58 plus.n19 plus.n18 0.189894
R59 plus.n30 plus.n19 0.189894
R60 plus.n30 plus.n29 0.189894
R61 plus.n29 plus.n28 0.189894
R62 plus.n28 plus.n21 0.189894
R63 plus.n24 plus.n21 0.189894
R64 drain_left.n6 drain_left.n4 68.0787
R65 drain_left.n3 drain_left.n2 68.0232
R66 drain_left.n3 drain_left.n0 68.0232
R67 drain_left.n6 drain_left.n5 67.1908
R68 drain_left.n8 drain_left.n7 67.1907
R69 drain_left.n3 drain_left.n1 67.1907
R70 drain_left drain_left.n3 27.2613
R71 drain_left drain_left.n8 6.54115
R72 drain_left.n1 drain_left.t5 3.3005
R73 drain_left.n1 drain_left.t6 3.3005
R74 drain_left.n2 drain_left.t7 3.3005
R75 drain_left.n2 drain_left.t1 3.3005
R76 drain_left.n0 drain_left.t11 3.3005
R77 drain_left.n0 drain_left.t3 3.3005
R78 drain_left.n7 drain_left.t2 3.3005
R79 drain_left.n7 drain_left.t9 3.3005
R80 drain_left.n5 drain_left.t4 3.3005
R81 drain_left.n5 drain_left.t8 3.3005
R82 drain_left.n4 drain_left.t10 3.3005
R83 drain_left.n4 drain_left.t0 3.3005
R84 drain_left.n8 drain_left.n6 0.888431
R85 source.n266 source.n240 289.615
R86 source.n230 source.n204 289.615
R87 source.n198 source.n172 289.615
R88 source.n162 source.n136 289.615
R89 source.n26 source.n0 289.615
R90 source.n62 source.n36 289.615
R91 source.n94 source.n68 289.615
R92 source.n130 source.n104 289.615
R93 source.n251 source.n250 185
R94 source.n248 source.n247 185
R95 source.n257 source.n256 185
R96 source.n259 source.n258 185
R97 source.n244 source.n243 185
R98 source.n265 source.n264 185
R99 source.n267 source.n266 185
R100 source.n215 source.n214 185
R101 source.n212 source.n211 185
R102 source.n221 source.n220 185
R103 source.n223 source.n222 185
R104 source.n208 source.n207 185
R105 source.n229 source.n228 185
R106 source.n231 source.n230 185
R107 source.n183 source.n182 185
R108 source.n180 source.n179 185
R109 source.n189 source.n188 185
R110 source.n191 source.n190 185
R111 source.n176 source.n175 185
R112 source.n197 source.n196 185
R113 source.n199 source.n198 185
R114 source.n147 source.n146 185
R115 source.n144 source.n143 185
R116 source.n153 source.n152 185
R117 source.n155 source.n154 185
R118 source.n140 source.n139 185
R119 source.n161 source.n160 185
R120 source.n163 source.n162 185
R121 source.n27 source.n26 185
R122 source.n25 source.n24 185
R123 source.n4 source.n3 185
R124 source.n19 source.n18 185
R125 source.n17 source.n16 185
R126 source.n8 source.n7 185
R127 source.n11 source.n10 185
R128 source.n63 source.n62 185
R129 source.n61 source.n60 185
R130 source.n40 source.n39 185
R131 source.n55 source.n54 185
R132 source.n53 source.n52 185
R133 source.n44 source.n43 185
R134 source.n47 source.n46 185
R135 source.n95 source.n94 185
R136 source.n93 source.n92 185
R137 source.n72 source.n71 185
R138 source.n87 source.n86 185
R139 source.n85 source.n84 185
R140 source.n76 source.n75 185
R141 source.n79 source.n78 185
R142 source.n131 source.n130 185
R143 source.n129 source.n128 185
R144 source.n108 source.n107 185
R145 source.n123 source.n122 185
R146 source.n121 source.n120 185
R147 source.n112 source.n111 185
R148 source.n115 source.n114 185
R149 source.t1 source.n249 147.661
R150 source.t4 source.n213 147.661
R151 source.t14 source.n181 147.661
R152 source.t9 source.n145 147.661
R153 source.t11 source.n9 147.661
R154 source.t16 source.n45 147.661
R155 source.t6 source.n77 147.661
R156 source.t3 source.n113 147.661
R157 source.n250 source.n247 104.615
R158 source.n257 source.n247 104.615
R159 source.n258 source.n257 104.615
R160 source.n258 source.n243 104.615
R161 source.n265 source.n243 104.615
R162 source.n266 source.n265 104.615
R163 source.n214 source.n211 104.615
R164 source.n221 source.n211 104.615
R165 source.n222 source.n221 104.615
R166 source.n222 source.n207 104.615
R167 source.n229 source.n207 104.615
R168 source.n230 source.n229 104.615
R169 source.n182 source.n179 104.615
R170 source.n189 source.n179 104.615
R171 source.n190 source.n189 104.615
R172 source.n190 source.n175 104.615
R173 source.n197 source.n175 104.615
R174 source.n198 source.n197 104.615
R175 source.n146 source.n143 104.615
R176 source.n153 source.n143 104.615
R177 source.n154 source.n153 104.615
R178 source.n154 source.n139 104.615
R179 source.n161 source.n139 104.615
R180 source.n162 source.n161 104.615
R181 source.n26 source.n25 104.615
R182 source.n25 source.n3 104.615
R183 source.n18 source.n3 104.615
R184 source.n18 source.n17 104.615
R185 source.n17 source.n7 104.615
R186 source.n10 source.n7 104.615
R187 source.n62 source.n61 104.615
R188 source.n61 source.n39 104.615
R189 source.n54 source.n39 104.615
R190 source.n54 source.n53 104.615
R191 source.n53 source.n43 104.615
R192 source.n46 source.n43 104.615
R193 source.n94 source.n93 104.615
R194 source.n93 source.n71 104.615
R195 source.n86 source.n71 104.615
R196 source.n86 source.n85 104.615
R197 source.n85 source.n75 104.615
R198 source.n78 source.n75 104.615
R199 source.n130 source.n129 104.615
R200 source.n129 source.n107 104.615
R201 source.n122 source.n107 104.615
R202 source.n122 source.n121 104.615
R203 source.n121 source.n111 104.615
R204 source.n114 source.n111 104.615
R205 source.n250 source.t1 52.3082
R206 source.n214 source.t4 52.3082
R207 source.n182 source.t14 52.3082
R208 source.n146 source.t9 52.3082
R209 source.n10 source.t11 52.3082
R210 source.n46 source.t16 52.3082
R211 source.n78 source.t6 52.3082
R212 source.n114 source.t3 52.3082
R213 source.n33 source.n32 50.512
R214 source.n35 source.n34 50.512
R215 source.n101 source.n100 50.512
R216 source.n103 source.n102 50.512
R217 source.n239 source.n238 50.5119
R218 source.n237 source.n236 50.5119
R219 source.n171 source.n170 50.5119
R220 source.n169 source.n168 50.5119
R221 source.n271 source.n270 32.1853
R222 source.n235 source.n234 32.1853
R223 source.n203 source.n202 32.1853
R224 source.n167 source.n166 32.1853
R225 source.n31 source.n30 32.1853
R226 source.n67 source.n66 32.1853
R227 source.n99 source.n98 32.1853
R228 source.n135 source.n134 32.1853
R229 source.n167 source.n135 17.6302
R230 source.n251 source.n249 15.6674
R231 source.n215 source.n213 15.6674
R232 source.n183 source.n181 15.6674
R233 source.n147 source.n145 15.6674
R234 source.n11 source.n9 15.6674
R235 source.n47 source.n45 15.6674
R236 source.n79 source.n77 15.6674
R237 source.n115 source.n113 15.6674
R238 source.n252 source.n248 12.8005
R239 source.n216 source.n212 12.8005
R240 source.n184 source.n180 12.8005
R241 source.n148 source.n144 12.8005
R242 source.n12 source.n8 12.8005
R243 source.n48 source.n44 12.8005
R244 source.n80 source.n76 12.8005
R245 source.n116 source.n112 12.8005
R246 source.n256 source.n255 12.0247
R247 source.n220 source.n219 12.0247
R248 source.n188 source.n187 12.0247
R249 source.n152 source.n151 12.0247
R250 source.n16 source.n15 12.0247
R251 source.n52 source.n51 12.0247
R252 source.n84 source.n83 12.0247
R253 source.n120 source.n119 12.0247
R254 source.n272 source.n31 11.9233
R255 source.n259 source.n246 11.249
R256 source.n223 source.n210 11.249
R257 source.n191 source.n178 11.249
R258 source.n155 source.n142 11.249
R259 source.n19 source.n6 11.249
R260 source.n55 source.n42 11.249
R261 source.n87 source.n74 11.249
R262 source.n123 source.n110 11.249
R263 source.n260 source.n244 10.4732
R264 source.n224 source.n208 10.4732
R265 source.n192 source.n176 10.4732
R266 source.n156 source.n140 10.4732
R267 source.n20 source.n4 10.4732
R268 source.n56 source.n40 10.4732
R269 source.n88 source.n72 10.4732
R270 source.n124 source.n108 10.4732
R271 source.n264 source.n263 9.69747
R272 source.n228 source.n227 9.69747
R273 source.n196 source.n195 9.69747
R274 source.n160 source.n159 9.69747
R275 source.n24 source.n23 9.69747
R276 source.n60 source.n59 9.69747
R277 source.n92 source.n91 9.69747
R278 source.n128 source.n127 9.69747
R279 source.n270 source.n269 9.45567
R280 source.n234 source.n233 9.45567
R281 source.n202 source.n201 9.45567
R282 source.n166 source.n165 9.45567
R283 source.n30 source.n29 9.45567
R284 source.n66 source.n65 9.45567
R285 source.n98 source.n97 9.45567
R286 source.n134 source.n133 9.45567
R287 source.n269 source.n268 9.3005
R288 source.n242 source.n241 9.3005
R289 source.n263 source.n262 9.3005
R290 source.n261 source.n260 9.3005
R291 source.n246 source.n245 9.3005
R292 source.n255 source.n254 9.3005
R293 source.n253 source.n252 9.3005
R294 source.n233 source.n232 9.3005
R295 source.n206 source.n205 9.3005
R296 source.n227 source.n226 9.3005
R297 source.n225 source.n224 9.3005
R298 source.n210 source.n209 9.3005
R299 source.n219 source.n218 9.3005
R300 source.n217 source.n216 9.3005
R301 source.n201 source.n200 9.3005
R302 source.n174 source.n173 9.3005
R303 source.n195 source.n194 9.3005
R304 source.n193 source.n192 9.3005
R305 source.n178 source.n177 9.3005
R306 source.n187 source.n186 9.3005
R307 source.n185 source.n184 9.3005
R308 source.n165 source.n164 9.3005
R309 source.n138 source.n137 9.3005
R310 source.n159 source.n158 9.3005
R311 source.n157 source.n156 9.3005
R312 source.n142 source.n141 9.3005
R313 source.n151 source.n150 9.3005
R314 source.n149 source.n148 9.3005
R315 source.n29 source.n28 9.3005
R316 source.n2 source.n1 9.3005
R317 source.n23 source.n22 9.3005
R318 source.n21 source.n20 9.3005
R319 source.n6 source.n5 9.3005
R320 source.n15 source.n14 9.3005
R321 source.n13 source.n12 9.3005
R322 source.n65 source.n64 9.3005
R323 source.n38 source.n37 9.3005
R324 source.n59 source.n58 9.3005
R325 source.n57 source.n56 9.3005
R326 source.n42 source.n41 9.3005
R327 source.n51 source.n50 9.3005
R328 source.n49 source.n48 9.3005
R329 source.n97 source.n96 9.3005
R330 source.n70 source.n69 9.3005
R331 source.n91 source.n90 9.3005
R332 source.n89 source.n88 9.3005
R333 source.n74 source.n73 9.3005
R334 source.n83 source.n82 9.3005
R335 source.n81 source.n80 9.3005
R336 source.n133 source.n132 9.3005
R337 source.n106 source.n105 9.3005
R338 source.n127 source.n126 9.3005
R339 source.n125 source.n124 9.3005
R340 source.n110 source.n109 9.3005
R341 source.n119 source.n118 9.3005
R342 source.n117 source.n116 9.3005
R343 source.n267 source.n242 8.92171
R344 source.n231 source.n206 8.92171
R345 source.n199 source.n174 8.92171
R346 source.n163 source.n138 8.92171
R347 source.n27 source.n2 8.92171
R348 source.n63 source.n38 8.92171
R349 source.n95 source.n70 8.92171
R350 source.n131 source.n106 8.92171
R351 source.n268 source.n240 8.14595
R352 source.n232 source.n204 8.14595
R353 source.n200 source.n172 8.14595
R354 source.n164 source.n136 8.14595
R355 source.n28 source.n0 8.14595
R356 source.n64 source.n36 8.14595
R357 source.n96 source.n68 8.14595
R358 source.n132 source.n104 8.14595
R359 source.n270 source.n240 5.81868
R360 source.n234 source.n204 5.81868
R361 source.n202 source.n172 5.81868
R362 source.n166 source.n136 5.81868
R363 source.n30 source.n0 5.81868
R364 source.n66 source.n36 5.81868
R365 source.n98 source.n68 5.81868
R366 source.n134 source.n104 5.81868
R367 source.n272 source.n271 5.7074
R368 source.n268 source.n267 5.04292
R369 source.n232 source.n231 5.04292
R370 source.n200 source.n199 5.04292
R371 source.n164 source.n163 5.04292
R372 source.n28 source.n27 5.04292
R373 source.n64 source.n63 5.04292
R374 source.n96 source.n95 5.04292
R375 source.n132 source.n131 5.04292
R376 source.n253 source.n249 4.38594
R377 source.n217 source.n213 4.38594
R378 source.n185 source.n181 4.38594
R379 source.n149 source.n145 4.38594
R380 source.n13 source.n9 4.38594
R381 source.n49 source.n45 4.38594
R382 source.n81 source.n77 4.38594
R383 source.n117 source.n113 4.38594
R384 source.n264 source.n242 4.26717
R385 source.n228 source.n206 4.26717
R386 source.n196 source.n174 4.26717
R387 source.n160 source.n138 4.26717
R388 source.n24 source.n2 4.26717
R389 source.n60 source.n38 4.26717
R390 source.n92 source.n70 4.26717
R391 source.n128 source.n106 4.26717
R392 source.n263 source.n244 3.49141
R393 source.n227 source.n208 3.49141
R394 source.n195 source.n176 3.49141
R395 source.n159 source.n140 3.49141
R396 source.n23 source.n4 3.49141
R397 source.n59 source.n40 3.49141
R398 source.n91 source.n72 3.49141
R399 source.n127 source.n108 3.49141
R400 source.n238 source.t2 3.3005
R401 source.n238 source.t7 3.3005
R402 source.n236 source.t5 3.3005
R403 source.n236 source.t22 3.3005
R404 source.n170 source.t15 3.3005
R405 source.n170 source.t13 3.3005
R406 source.n168 source.t18 3.3005
R407 source.n168 source.t20 3.3005
R408 source.n32 source.t12 3.3005
R409 source.n32 source.t17 3.3005
R410 source.n34 source.t10 3.3005
R411 source.n34 source.t19 3.3005
R412 source.n100 source.t21 3.3005
R413 source.n100 source.t23 3.3005
R414 source.n102 source.t0 3.3005
R415 source.n102 source.t8 3.3005
R416 source.n260 source.n259 2.71565
R417 source.n224 source.n223 2.71565
R418 source.n192 source.n191 2.71565
R419 source.n156 source.n155 2.71565
R420 source.n20 source.n19 2.71565
R421 source.n56 source.n55 2.71565
R422 source.n88 source.n87 2.71565
R423 source.n124 source.n123 2.71565
R424 source.n256 source.n246 1.93989
R425 source.n220 source.n210 1.93989
R426 source.n188 source.n178 1.93989
R427 source.n152 source.n142 1.93989
R428 source.n16 source.n6 1.93989
R429 source.n52 source.n42 1.93989
R430 source.n84 source.n74 1.93989
R431 source.n120 source.n110 1.93989
R432 source.n255 source.n248 1.16414
R433 source.n219 source.n212 1.16414
R434 source.n187 source.n180 1.16414
R435 source.n151 source.n144 1.16414
R436 source.n15 source.n8 1.16414
R437 source.n51 source.n44 1.16414
R438 source.n83 source.n76 1.16414
R439 source.n119 source.n112 1.16414
R440 source.n135 source.n103 0.888431
R441 source.n103 source.n101 0.888431
R442 source.n101 source.n99 0.888431
R443 source.n67 source.n35 0.888431
R444 source.n35 source.n33 0.888431
R445 source.n33 source.n31 0.888431
R446 source.n169 source.n167 0.888431
R447 source.n171 source.n169 0.888431
R448 source.n203 source.n171 0.888431
R449 source.n237 source.n235 0.888431
R450 source.n239 source.n237 0.888431
R451 source.n271 source.n239 0.888431
R452 source.n99 source.n67 0.470328
R453 source.n235 source.n203 0.470328
R454 source.n252 source.n251 0.388379
R455 source.n216 source.n215 0.388379
R456 source.n184 source.n183 0.388379
R457 source.n148 source.n147 0.388379
R458 source.n12 source.n11 0.388379
R459 source.n48 source.n47 0.388379
R460 source.n80 source.n79 0.388379
R461 source.n116 source.n115 0.388379
R462 source source.n272 0.188
R463 source.n254 source.n253 0.155672
R464 source.n254 source.n245 0.155672
R465 source.n261 source.n245 0.155672
R466 source.n262 source.n261 0.155672
R467 source.n262 source.n241 0.155672
R468 source.n269 source.n241 0.155672
R469 source.n218 source.n217 0.155672
R470 source.n218 source.n209 0.155672
R471 source.n225 source.n209 0.155672
R472 source.n226 source.n225 0.155672
R473 source.n226 source.n205 0.155672
R474 source.n233 source.n205 0.155672
R475 source.n186 source.n185 0.155672
R476 source.n186 source.n177 0.155672
R477 source.n193 source.n177 0.155672
R478 source.n194 source.n193 0.155672
R479 source.n194 source.n173 0.155672
R480 source.n201 source.n173 0.155672
R481 source.n150 source.n149 0.155672
R482 source.n150 source.n141 0.155672
R483 source.n157 source.n141 0.155672
R484 source.n158 source.n157 0.155672
R485 source.n158 source.n137 0.155672
R486 source.n165 source.n137 0.155672
R487 source.n29 source.n1 0.155672
R488 source.n22 source.n1 0.155672
R489 source.n22 source.n21 0.155672
R490 source.n21 source.n5 0.155672
R491 source.n14 source.n5 0.155672
R492 source.n14 source.n13 0.155672
R493 source.n65 source.n37 0.155672
R494 source.n58 source.n37 0.155672
R495 source.n58 source.n57 0.155672
R496 source.n57 source.n41 0.155672
R497 source.n50 source.n41 0.155672
R498 source.n50 source.n49 0.155672
R499 source.n97 source.n69 0.155672
R500 source.n90 source.n69 0.155672
R501 source.n90 source.n89 0.155672
R502 source.n89 source.n73 0.155672
R503 source.n82 source.n73 0.155672
R504 source.n82 source.n81 0.155672
R505 source.n133 source.n105 0.155672
R506 source.n126 source.n105 0.155672
R507 source.n126 source.n125 0.155672
R508 source.n125 source.n109 0.155672
R509 source.n118 source.n109 0.155672
R510 source.n118 source.n117 0.155672
R511 minus.n5 minus.t6 285.995
R512 minus.n23 minus.t8 285.995
R513 minus.n4 minus.t0 262.69
R514 minus.n8 minus.t3 262.69
R515 minus.n10 minus.t10 262.69
R516 minus.n14 minus.t2 262.69
R517 minus.n16 minus.t11 262.69
R518 minus.n22 minus.t9 262.69
R519 minus.n26 minus.t4 262.69
R520 minus.n28 minus.t5 262.69
R521 minus.n32 minus.t7 262.69
R522 minus.n34 minus.t1 262.69
R523 minus.n17 minus.n16 161.3
R524 minus.n15 minus.n0 161.3
R525 minus.n14 minus.n13 161.3
R526 minus.n12 minus.n1 161.3
R527 minus.n11 minus.n10 161.3
R528 minus.n9 minus.n2 161.3
R529 minus.n8 minus.n7 161.3
R530 minus.n6 minus.n3 161.3
R531 minus.n35 minus.n34 161.3
R532 minus.n33 minus.n18 161.3
R533 minus.n32 minus.n31 161.3
R534 minus.n30 minus.n19 161.3
R535 minus.n29 minus.n28 161.3
R536 minus.n27 minus.n20 161.3
R537 minus.n26 minus.n25 161.3
R538 minus.n24 minus.n21 161.3
R539 minus.n6 minus.n5 44.8907
R540 minus.n24 minus.n23 44.8907
R541 minus.n36 minus.n17 32.8944
R542 minus.n16 minus.n15 32.8641
R543 minus.n34 minus.n33 32.8641
R544 minus.n4 minus.n3 28.4823
R545 minus.n14 minus.n1 28.4823
R546 minus.n22 minus.n21 28.4823
R547 minus.n32 minus.n19 28.4823
R548 minus.n10 minus.n9 24.1005
R549 minus.n9 minus.n8 24.1005
R550 minus.n27 minus.n26 24.1005
R551 minus.n28 minus.n27 24.1005
R552 minus.n8 minus.n3 19.7187
R553 minus.n10 minus.n1 19.7187
R554 minus.n26 minus.n21 19.7187
R555 minus.n28 minus.n19 19.7187
R556 minus.n5 minus.n4 18.4104
R557 minus.n23 minus.n22 18.4104
R558 minus.n15 minus.n14 15.3369
R559 minus.n33 minus.n32 15.3369
R560 minus.n36 minus.n35 6.64444
R561 minus.n17 minus.n0 0.189894
R562 minus.n13 minus.n0 0.189894
R563 minus.n13 minus.n12 0.189894
R564 minus.n12 minus.n11 0.189894
R565 minus.n11 minus.n2 0.189894
R566 minus.n7 minus.n2 0.189894
R567 minus.n7 minus.n6 0.189894
R568 minus.n25 minus.n24 0.189894
R569 minus.n25 minus.n20 0.189894
R570 minus.n29 minus.n20 0.189894
R571 minus.n30 minus.n29 0.189894
R572 minus.n31 minus.n30 0.189894
R573 minus.n31 minus.n18 0.189894
R574 minus.n35 minus.n18 0.189894
R575 minus minus.n36 0.188
R576 drain_right.n6 drain_right.n4 68.0786
R577 drain_right.n3 drain_right.n2 68.0232
R578 drain_right.n3 drain_right.n0 68.0232
R579 drain_right.n6 drain_right.n5 67.1908
R580 drain_right.n8 drain_right.n7 67.1908
R581 drain_right.n3 drain_right.n1 67.1907
R582 drain_right drain_right.n3 26.708
R583 drain_right drain_right.n8 6.54115
R584 drain_right.n1 drain_right.t7 3.3005
R585 drain_right.n1 drain_right.t6 3.3005
R586 drain_right.n2 drain_right.t4 3.3005
R587 drain_right.n2 drain_right.t10 3.3005
R588 drain_right.n0 drain_right.t3 3.3005
R589 drain_right.n0 drain_right.t2 3.3005
R590 drain_right.n4 drain_right.t11 3.3005
R591 drain_right.n4 drain_right.t5 3.3005
R592 drain_right.n5 drain_right.t1 3.3005
R593 drain_right.n5 drain_right.t8 3.3005
R594 drain_right.n7 drain_right.t0 3.3005
R595 drain_right.n7 drain_right.t9 3.3005
R596 drain_right.n8 drain_right.n6 0.888431
C0 drain_left source 9.15878f
C1 minus plus 4.72368f
C2 drain_right source 9.160821f
C3 drain_left plus 4.40447f
C4 drain_left minus 0.17184f
C5 drain_right plus 0.366822f
C6 drain_right minus 4.19273f
C7 drain_right drain_left 1.08491f
C8 source plus 4.41473f
C9 source minus 4.40071f
C10 drain_right a_n2158_n2088# 5.05296f
C11 drain_left a_n2158_n2088# 5.36763f
C12 source a_n2158_n2088# 5.535097f
C13 minus a_n2158_n2088# 8.008983f
C14 plus a_n2158_n2088# 9.42151f
C15 drain_right.t3 a_n2158_n2088# 0.127683f
C16 drain_right.t2 a_n2158_n2088# 0.127683f
C17 drain_right.n0 a_n2158_n2088# 1.06952f
C18 drain_right.t7 a_n2158_n2088# 0.127683f
C19 drain_right.t6 a_n2158_n2088# 0.127683f
C20 drain_right.n1 a_n2158_n2088# 1.06488f
C21 drain_right.t4 a_n2158_n2088# 0.127683f
C22 drain_right.t10 a_n2158_n2088# 0.127683f
C23 drain_right.n2 a_n2158_n2088# 1.06952f
C24 drain_right.n3 a_n2158_n2088# 2.07117f
C25 drain_right.t11 a_n2158_n2088# 0.127683f
C26 drain_right.t5 a_n2158_n2088# 0.127683f
C27 drain_right.n4 a_n2158_n2088# 1.06988f
C28 drain_right.t1 a_n2158_n2088# 0.127683f
C29 drain_right.t8 a_n2158_n2088# 0.127683f
C30 drain_right.n5 a_n2158_n2088# 1.06488f
C31 drain_right.n6 a_n2158_n2088# 0.751171f
C32 drain_right.t0 a_n2158_n2088# 0.127683f
C33 drain_right.t9 a_n2158_n2088# 0.127683f
C34 drain_right.n7 a_n2158_n2088# 1.06488f
C35 drain_right.n8 a_n2158_n2088# 0.610853f
C36 minus.n0 a_n2158_n2088# 0.042703f
C37 minus.n1 a_n2158_n2088# 0.00969f
C38 minus.t2 a_n2158_n2088# 0.520227f
C39 minus.n2 a_n2158_n2088# 0.042703f
C40 minus.n3 a_n2158_n2088# 0.00969f
C41 minus.t3 a_n2158_n2088# 0.520227f
C42 minus.t6 a_n2158_n2088# 0.539811f
C43 minus.t0 a_n2158_n2088# 0.520227f
C44 minus.n4 a_n2158_n2088# 0.245168f
C45 minus.n5 a_n2158_n2088# 0.224631f
C46 minus.n6 a_n2158_n2088# 0.179146f
C47 minus.n7 a_n2158_n2088# 0.042703f
C48 minus.n8 a_n2158_n2088# 0.240392f
C49 minus.n9 a_n2158_n2088# 0.00969f
C50 minus.t10 a_n2158_n2088# 0.520227f
C51 minus.n10 a_n2158_n2088# 0.240392f
C52 minus.n11 a_n2158_n2088# 0.042703f
C53 minus.n12 a_n2158_n2088# 0.042703f
C54 minus.n13 a_n2158_n2088# 0.042703f
C55 minus.n14 a_n2158_n2088# 0.240392f
C56 minus.n15 a_n2158_n2088# 0.00969f
C57 minus.t11 a_n2158_n2088# 0.520227f
C58 minus.n16 a_n2158_n2088# 0.238417f
C59 minus.n17 a_n2158_n2088# 1.30075f
C60 minus.n18 a_n2158_n2088# 0.042703f
C61 minus.n19 a_n2158_n2088# 0.00969f
C62 minus.n20 a_n2158_n2088# 0.042703f
C63 minus.n21 a_n2158_n2088# 0.00969f
C64 minus.t8 a_n2158_n2088# 0.539811f
C65 minus.t9 a_n2158_n2088# 0.520227f
C66 minus.n22 a_n2158_n2088# 0.245168f
C67 minus.n23 a_n2158_n2088# 0.224631f
C68 minus.n24 a_n2158_n2088# 0.179146f
C69 minus.n25 a_n2158_n2088# 0.042703f
C70 minus.t4 a_n2158_n2088# 0.520227f
C71 minus.n26 a_n2158_n2088# 0.240392f
C72 minus.n27 a_n2158_n2088# 0.00969f
C73 minus.t5 a_n2158_n2088# 0.520227f
C74 minus.n28 a_n2158_n2088# 0.240392f
C75 minus.n29 a_n2158_n2088# 0.042703f
C76 minus.n30 a_n2158_n2088# 0.042703f
C77 minus.n31 a_n2158_n2088# 0.042703f
C78 minus.t7 a_n2158_n2088# 0.520227f
C79 minus.n32 a_n2158_n2088# 0.240392f
C80 minus.n33 a_n2158_n2088# 0.00969f
C81 minus.t1 a_n2158_n2088# 0.520227f
C82 minus.n34 a_n2158_n2088# 0.238417f
C83 minus.n35 a_n2158_n2088# 0.293618f
C84 minus.n36 a_n2158_n2088# 1.58866f
C85 source.n0 a_n2158_n2088# 0.033547f
C86 source.n1 a_n2158_n2088# 0.023867f
C87 source.n2 a_n2158_n2088# 0.012825f
C88 source.n3 a_n2158_n2088# 0.030314f
C89 source.n4 a_n2158_n2088# 0.01358f
C90 source.n5 a_n2158_n2088# 0.023867f
C91 source.n6 a_n2158_n2088# 0.012825f
C92 source.n7 a_n2158_n2088# 0.030314f
C93 source.n8 a_n2158_n2088# 0.01358f
C94 source.n9 a_n2158_n2088# 0.102134f
C95 source.t11 a_n2158_n2088# 0.049408f
C96 source.n10 a_n2158_n2088# 0.022736f
C97 source.n11 a_n2158_n2088# 0.017906f
C98 source.n12 a_n2158_n2088# 0.012825f
C99 source.n13 a_n2158_n2088# 0.567895f
C100 source.n14 a_n2158_n2088# 0.023867f
C101 source.n15 a_n2158_n2088# 0.012825f
C102 source.n16 a_n2158_n2088# 0.01358f
C103 source.n17 a_n2158_n2088# 0.030314f
C104 source.n18 a_n2158_n2088# 0.030314f
C105 source.n19 a_n2158_n2088# 0.01358f
C106 source.n20 a_n2158_n2088# 0.012825f
C107 source.n21 a_n2158_n2088# 0.023867f
C108 source.n22 a_n2158_n2088# 0.023867f
C109 source.n23 a_n2158_n2088# 0.012825f
C110 source.n24 a_n2158_n2088# 0.01358f
C111 source.n25 a_n2158_n2088# 0.030314f
C112 source.n26 a_n2158_n2088# 0.065625f
C113 source.n27 a_n2158_n2088# 0.01358f
C114 source.n28 a_n2158_n2088# 0.012825f
C115 source.n29 a_n2158_n2088# 0.055168f
C116 source.n30 a_n2158_n2088# 0.03672f
C117 source.n31 a_n2158_n2088# 0.623494f
C118 source.t12 a_n2158_n2088# 0.113163f
C119 source.t17 a_n2158_n2088# 0.113163f
C120 source.n32 a_n2158_n2088# 0.881323f
C121 source.n33 a_n2158_n2088# 0.360304f
C122 source.t10 a_n2158_n2088# 0.113163f
C123 source.t19 a_n2158_n2088# 0.113163f
C124 source.n34 a_n2158_n2088# 0.881323f
C125 source.n35 a_n2158_n2088# 0.360304f
C126 source.n36 a_n2158_n2088# 0.033547f
C127 source.n37 a_n2158_n2088# 0.023867f
C128 source.n38 a_n2158_n2088# 0.012825f
C129 source.n39 a_n2158_n2088# 0.030314f
C130 source.n40 a_n2158_n2088# 0.01358f
C131 source.n41 a_n2158_n2088# 0.023867f
C132 source.n42 a_n2158_n2088# 0.012825f
C133 source.n43 a_n2158_n2088# 0.030314f
C134 source.n44 a_n2158_n2088# 0.01358f
C135 source.n45 a_n2158_n2088# 0.102134f
C136 source.t16 a_n2158_n2088# 0.049408f
C137 source.n46 a_n2158_n2088# 0.022736f
C138 source.n47 a_n2158_n2088# 0.017906f
C139 source.n48 a_n2158_n2088# 0.012825f
C140 source.n49 a_n2158_n2088# 0.567895f
C141 source.n50 a_n2158_n2088# 0.023867f
C142 source.n51 a_n2158_n2088# 0.012825f
C143 source.n52 a_n2158_n2088# 0.01358f
C144 source.n53 a_n2158_n2088# 0.030314f
C145 source.n54 a_n2158_n2088# 0.030314f
C146 source.n55 a_n2158_n2088# 0.01358f
C147 source.n56 a_n2158_n2088# 0.012825f
C148 source.n57 a_n2158_n2088# 0.023867f
C149 source.n58 a_n2158_n2088# 0.023867f
C150 source.n59 a_n2158_n2088# 0.012825f
C151 source.n60 a_n2158_n2088# 0.01358f
C152 source.n61 a_n2158_n2088# 0.030314f
C153 source.n62 a_n2158_n2088# 0.065625f
C154 source.n63 a_n2158_n2088# 0.01358f
C155 source.n64 a_n2158_n2088# 0.012825f
C156 source.n65 a_n2158_n2088# 0.055168f
C157 source.n66 a_n2158_n2088# 0.03672f
C158 source.n67 a_n2158_n2088# 0.124803f
C159 source.n68 a_n2158_n2088# 0.033547f
C160 source.n69 a_n2158_n2088# 0.023867f
C161 source.n70 a_n2158_n2088# 0.012825f
C162 source.n71 a_n2158_n2088# 0.030314f
C163 source.n72 a_n2158_n2088# 0.01358f
C164 source.n73 a_n2158_n2088# 0.023867f
C165 source.n74 a_n2158_n2088# 0.012825f
C166 source.n75 a_n2158_n2088# 0.030314f
C167 source.n76 a_n2158_n2088# 0.01358f
C168 source.n77 a_n2158_n2088# 0.102134f
C169 source.t6 a_n2158_n2088# 0.049408f
C170 source.n78 a_n2158_n2088# 0.022736f
C171 source.n79 a_n2158_n2088# 0.017906f
C172 source.n80 a_n2158_n2088# 0.012825f
C173 source.n81 a_n2158_n2088# 0.567895f
C174 source.n82 a_n2158_n2088# 0.023867f
C175 source.n83 a_n2158_n2088# 0.012825f
C176 source.n84 a_n2158_n2088# 0.01358f
C177 source.n85 a_n2158_n2088# 0.030314f
C178 source.n86 a_n2158_n2088# 0.030314f
C179 source.n87 a_n2158_n2088# 0.01358f
C180 source.n88 a_n2158_n2088# 0.012825f
C181 source.n89 a_n2158_n2088# 0.023867f
C182 source.n90 a_n2158_n2088# 0.023867f
C183 source.n91 a_n2158_n2088# 0.012825f
C184 source.n92 a_n2158_n2088# 0.01358f
C185 source.n93 a_n2158_n2088# 0.030314f
C186 source.n94 a_n2158_n2088# 0.065625f
C187 source.n95 a_n2158_n2088# 0.01358f
C188 source.n96 a_n2158_n2088# 0.012825f
C189 source.n97 a_n2158_n2088# 0.055168f
C190 source.n98 a_n2158_n2088# 0.03672f
C191 source.n99 a_n2158_n2088# 0.124803f
C192 source.t21 a_n2158_n2088# 0.113163f
C193 source.t23 a_n2158_n2088# 0.113163f
C194 source.n100 a_n2158_n2088# 0.881323f
C195 source.n101 a_n2158_n2088# 0.360304f
C196 source.t0 a_n2158_n2088# 0.113163f
C197 source.t8 a_n2158_n2088# 0.113163f
C198 source.n102 a_n2158_n2088# 0.881323f
C199 source.n103 a_n2158_n2088# 0.360304f
C200 source.n104 a_n2158_n2088# 0.033547f
C201 source.n105 a_n2158_n2088# 0.023867f
C202 source.n106 a_n2158_n2088# 0.012825f
C203 source.n107 a_n2158_n2088# 0.030314f
C204 source.n108 a_n2158_n2088# 0.01358f
C205 source.n109 a_n2158_n2088# 0.023867f
C206 source.n110 a_n2158_n2088# 0.012825f
C207 source.n111 a_n2158_n2088# 0.030314f
C208 source.n112 a_n2158_n2088# 0.01358f
C209 source.n113 a_n2158_n2088# 0.102134f
C210 source.t3 a_n2158_n2088# 0.049408f
C211 source.n114 a_n2158_n2088# 0.022736f
C212 source.n115 a_n2158_n2088# 0.017906f
C213 source.n116 a_n2158_n2088# 0.012825f
C214 source.n117 a_n2158_n2088# 0.567895f
C215 source.n118 a_n2158_n2088# 0.023867f
C216 source.n119 a_n2158_n2088# 0.012825f
C217 source.n120 a_n2158_n2088# 0.01358f
C218 source.n121 a_n2158_n2088# 0.030314f
C219 source.n122 a_n2158_n2088# 0.030314f
C220 source.n123 a_n2158_n2088# 0.01358f
C221 source.n124 a_n2158_n2088# 0.012825f
C222 source.n125 a_n2158_n2088# 0.023867f
C223 source.n126 a_n2158_n2088# 0.023867f
C224 source.n127 a_n2158_n2088# 0.012825f
C225 source.n128 a_n2158_n2088# 0.01358f
C226 source.n129 a_n2158_n2088# 0.030314f
C227 source.n130 a_n2158_n2088# 0.065625f
C228 source.n131 a_n2158_n2088# 0.01358f
C229 source.n132 a_n2158_n2088# 0.012825f
C230 source.n133 a_n2158_n2088# 0.055168f
C231 source.n134 a_n2158_n2088# 0.03672f
C232 source.n135 a_n2158_n2088# 0.938411f
C233 source.n136 a_n2158_n2088# 0.033547f
C234 source.n137 a_n2158_n2088# 0.023867f
C235 source.n138 a_n2158_n2088# 0.012825f
C236 source.n139 a_n2158_n2088# 0.030314f
C237 source.n140 a_n2158_n2088# 0.01358f
C238 source.n141 a_n2158_n2088# 0.023867f
C239 source.n142 a_n2158_n2088# 0.012825f
C240 source.n143 a_n2158_n2088# 0.030314f
C241 source.n144 a_n2158_n2088# 0.01358f
C242 source.n145 a_n2158_n2088# 0.102134f
C243 source.t9 a_n2158_n2088# 0.049408f
C244 source.n146 a_n2158_n2088# 0.022736f
C245 source.n147 a_n2158_n2088# 0.017906f
C246 source.n148 a_n2158_n2088# 0.012825f
C247 source.n149 a_n2158_n2088# 0.567895f
C248 source.n150 a_n2158_n2088# 0.023867f
C249 source.n151 a_n2158_n2088# 0.012825f
C250 source.n152 a_n2158_n2088# 0.01358f
C251 source.n153 a_n2158_n2088# 0.030314f
C252 source.n154 a_n2158_n2088# 0.030314f
C253 source.n155 a_n2158_n2088# 0.01358f
C254 source.n156 a_n2158_n2088# 0.012825f
C255 source.n157 a_n2158_n2088# 0.023867f
C256 source.n158 a_n2158_n2088# 0.023867f
C257 source.n159 a_n2158_n2088# 0.012825f
C258 source.n160 a_n2158_n2088# 0.01358f
C259 source.n161 a_n2158_n2088# 0.030314f
C260 source.n162 a_n2158_n2088# 0.065625f
C261 source.n163 a_n2158_n2088# 0.01358f
C262 source.n164 a_n2158_n2088# 0.012825f
C263 source.n165 a_n2158_n2088# 0.055168f
C264 source.n166 a_n2158_n2088# 0.03672f
C265 source.n167 a_n2158_n2088# 0.938411f
C266 source.t18 a_n2158_n2088# 0.113163f
C267 source.t20 a_n2158_n2088# 0.113163f
C268 source.n168 a_n2158_n2088# 0.881317f
C269 source.n169 a_n2158_n2088# 0.36031f
C270 source.t15 a_n2158_n2088# 0.113163f
C271 source.t13 a_n2158_n2088# 0.113163f
C272 source.n170 a_n2158_n2088# 0.881317f
C273 source.n171 a_n2158_n2088# 0.36031f
C274 source.n172 a_n2158_n2088# 0.033547f
C275 source.n173 a_n2158_n2088# 0.023867f
C276 source.n174 a_n2158_n2088# 0.012825f
C277 source.n175 a_n2158_n2088# 0.030314f
C278 source.n176 a_n2158_n2088# 0.01358f
C279 source.n177 a_n2158_n2088# 0.023867f
C280 source.n178 a_n2158_n2088# 0.012825f
C281 source.n179 a_n2158_n2088# 0.030314f
C282 source.n180 a_n2158_n2088# 0.01358f
C283 source.n181 a_n2158_n2088# 0.102134f
C284 source.t14 a_n2158_n2088# 0.049408f
C285 source.n182 a_n2158_n2088# 0.022736f
C286 source.n183 a_n2158_n2088# 0.017906f
C287 source.n184 a_n2158_n2088# 0.012825f
C288 source.n185 a_n2158_n2088# 0.567895f
C289 source.n186 a_n2158_n2088# 0.023867f
C290 source.n187 a_n2158_n2088# 0.012825f
C291 source.n188 a_n2158_n2088# 0.01358f
C292 source.n189 a_n2158_n2088# 0.030314f
C293 source.n190 a_n2158_n2088# 0.030314f
C294 source.n191 a_n2158_n2088# 0.01358f
C295 source.n192 a_n2158_n2088# 0.012825f
C296 source.n193 a_n2158_n2088# 0.023867f
C297 source.n194 a_n2158_n2088# 0.023867f
C298 source.n195 a_n2158_n2088# 0.012825f
C299 source.n196 a_n2158_n2088# 0.01358f
C300 source.n197 a_n2158_n2088# 0.030314f
C301 source.n198 a_n2158_n2088# 0.065625f
C302 source.n199 a_n2158_n2088# 0.01358f
C303 source.n200 a_n2158_n2088# 0.012825f
C304 source.n201 a_n2158_n2088# 0.055168f
C305 source.n202 a_n2158_n2088# 0.03672f
C306 source.n203 a_n2158_n2088# 0.124803f
C307 source.n204 a_n2158_n2088# 0.033547f
C308 source.n205 a_n2158_n2088# 0.023867f
C309 source.n206 a_n2158_n2088# 0.012825f
C310 source.n207 a_n2158_n2088# 0.030314f
C311 source.n208 a_n2158_n2088# 0.01358f
C312 source.n209 a_n2158_n2088# 0.023867f
C313 source.n210 a_n2158_n2088# 0.012825f
C314 source.n211 a_n2158_n2088# 0.030314f
C315 source.n212 a_n2158_n2088# 0.01358f
C316 source.n213 a_n2158_n2088# 0.102134f
C317 source.t4 a_n2158_n2088# 0.049408f
C318 source.n214 a_n2158_n2088# 0.022736f
C319 source.n215 a_n2158_n2088# 0.017906f
C320 source.n216 a_n2158_n2088# 0.012825f
C321 source.n217 a_n2158_n2088# 0.567895f
C322 source.n218 a_n2158_n2088# 0.023867f
C323 source.n219 a_n2158_n2088# 0.012825f
C324 source.n220 a_n2158_n2088# 0.01358f
C325 source.n221 a_n2158_n2088# 0.030314f
C326 source.n222 a_n2158_n2088# 0.030314f
C327 source.n223 a_n2158_n2088# 0.01358f
C328 source.n224 a_n2158_n2088# 0.012825f
C329 source.n225 a_n2158_n2088# 0.023867f
C330 source.n226 a_n2158_n2088# 0.023867f
C331 source.n227 a_n2158_n2088# 0.012825f
C332 source.n228 a_n2158_n2088# 0.01358f
C333 source.n229 a_n2158_n2088# 0.030314f
C334 source.n230 a_n2158_n2088# 0.065625f
C335 source.n231 a_n2158_n2088# 0.01358f
C336 source.n232 a_n2158_n2088# 0.012825f
C337 source.n233 a_n2158_n2088# 0.055168f
C338 source.n234 a_n2158_n2088# 0.03672f
C339 source.n235 a_n2158_n2088# 0.124803f
C340 source.t5 a_n2158_n2088# 0.113163f
C341 source.t22 a_n2158_n2088# 0.113163f
C342 source.n236 a_n2158_n2088# 0.881317f
C343 source.n237 a_n2158_n2088# 0.36031f
C344 source.t2 a_n2158_n2088# 0.113163f
C345 source.t7 a_n2158_n2088# 0.113163f
C346 source.n238 a_n2158_n2088# 0.881317f
C347 source.n239 a_n2158_n2088# 0.36031f
C348 source.n240 a_n2158_n2088# 0.033547f
C349 source.n241 a_n2158_n2088# 0.023867f
C350 source.n242 a_n2158_n2088# 0.012825f
C351 source.n243 a_n2158_n2088# 0.030314f
C352 source.n244 a_n2158_n2088# 0.01358f
C353 source.n245 a_n2158_n2088# 0.023867f
C354 source.n246 a_n2158_n2088# 0.012825f
C355 source.n247 a_n2158_n2088# 0.030314f
C356 source.n248 a_n2158_n2088# 0.01358f
C357 source.n249 a_n2158_n2088# 0.102134f
C358 source.t1 a_n2158_n2088# 0.049408f
C359 source.n250 a_n2158_n2088# 0.022736f
C360 source.n251 a_n2158_n2088# 0.017906f
C361 source.n252 a_n2158_n2088# 0.012825f
C362 source.n253 a_n2158_n2088# 0.567895f
C363 source.n254 a_n2158_n2088# 0.023867f
C364 source.n255 a_n2158_n2088# 0.012825f
C365 source.n256 a_n2158_n2088# 0.01358f
C366 source.n257 a_n2158_n2088# 0.030314f
C367 source.n258 a_n2158_n2088# 0.030314f
C368 source.n259 a_n2158_n2088# 0.01358f
C369 source.n260 a_n2158_n2088# 0.012825f
C370 source.n261 a_n2158_n2088# 0.023867f
C371 source.n262 a_n2158_n2088# 0.023867f
C372 source.n263 a_n2158_n2088# 0.012825f
C373 source.n264 a_n2158_n2088# 0.01358f
C374 source.n265 a_n2158_n2088# 0.030314f
C375 source.n266 a_n2158_n2088# 0.065625f
C376 source.n267 a_n2158_n2088# 0.01358f
C377 source.n268 a_n2158_n2088# 0.012825f
C378 source.n269 a_n2158_n2088# 0.055168f
C379 source.n270 a_n2158_n2088# 0.03672f
C380 source.n271 a_n2158_n2088# 0.280489f
C381 source.n272 a_n2158_n2088# 0.989815f
C382 drain_left.t11 a_n2158_n2088# 0.128578f
C383 drain_left.t3 a_n2158_n2088# 0.128578f
C384 drain_left.n0 a_n2158_n2088# 1.07702f
C385 drain_left.t5 a_n2158_n2088# 0.128578f
C386 drain_left.t6 a_n2158_n2088# 0.128578f
C387 drain_left.n1 a_n2158_n2088# 1.07234f
C388 drain_left.t7 a_n2158_n2088# 0.128578f
C389 drain_left.t1 a_n2158_n2088# 0.128578f
C390 drain_left.n2 a_n2158_n2088# 1.07702f
C391 drain_left.n3 a_n2158_n2088# 2.14046f
C392 drain_left.t10 a_n2158_n2088# 0.128578f
C393 drain_left.t0 a_n2158_n2088# 0.128578f
C394 drain_left.n4 a_n2158_n2088# 1.07738f
C395 drain_left.t4 a_n2158_n2088# 0.128578f
C396 drain_left.t8 a_n2158_n2088# 0.128578f
C397 drain_left.n5 a_n2158_n2088# 1.07234f
C398 drain_left.n6 a_n2158_n2088# 0.75643f
C399 drain_left.t2 a_n2158_n2088# 0.128578f
C400 drain_left.t9 a_n2158_n2088# 0.128578f
C401 drain_left.n7 a_n2158_n2088# 1.07234f
C402 drain_left.n8 a_n2158_n2088# 0.61514f
C403 plus.n0 a_n2158_n2088# 0.043629f
C404 plus.t9 a_n2158_n2088# 0.531501f
C405 plus.t3 a_n2158_n2088# 0.531501f
C406 plus.n1 a_n2158_n2088# 0.043629f
C407 plus.t8 a_n2158_n2088# 0.531501f
C408 plus.n2 a_n2158_n2088# 0.245601f
C409 plus.n3 a_n2158_n2088# 0.043629f
C410 plus.t1 a_n2158_n2088# 0.531501f
C411 plus.t10 a_n2158_n2088# 0.531501f
C412 plus.n4 a_n2158_n2088# 0.250481f
C413 plus.t4 a_n2158_n2088# 0.551509f
C414 plus.n5 a_n2158_n2088# 0.229499f
C415 plus.n6 a_n2158_n2088# 0.183028f
C416 plus.n7 a_n2158_n2088# 0.0099f
C417 plus.n8 a_n2158_n2088# 0.245601f
C418 plus.n9 a_n2158_n2088# 0.0099f
C419 plus.n10 a_n2158_n2088# 0.043629f
C420 plus.n11 a_n2158_n2088# 0.043629f
C421 plus.n12 a_n2158_n2088# 0.043629f
C422 plus.n13 a_n2158_n2088# 0.0099f
C423 plus.n14 a_n2158_n2088# 0.245601f
C424 plus.n15 a_n2158_n2088# 0.0099f
C425 plus.n16 a_n2158_n2088# 0.243584f
C426 plus.n17 a_n2158_n2088# 0.389263f
C427 plus.n18 a_n2158_n2088# 0.043629f
C428 plus.t11 a_n2158_n2088# 0.531501f
C429 plus.n19 a_n2158_n2088# 0.043629f
C430 plus.t2 a_n2158_n2088# 0.531501f
C431 plus.t0 a_n2158_n2088# 0.531501f
C432 plus.n20 a_n2158_n2088# 0.245601f
C433 plus.n21 a_n2158_n2088# 0.043629f
C434 plus.t5 a_n2158_n2088# 0.531501f
C435 plus.t7 a_n2158_n2088# 0.531501f
C436 plus.n22 a_n2158_n2088# 0.250481f
C437 plus.t6 a_n2158_n2088# 0.551509f
C438 plus.n23 a_n2158_n2088# 0.229499f
C439 plus.n24 a_n2158_n2088# 0.183028f
C440 plus.n25 a_n2158_n2088# 0.0099f
C441 plus.n26 a_n2158_n2088# 0.245601f
C442 plus.n27 a_n2158_n2088# 0.0099f
C443 plus.n28 a_n2158_n2088# 0.043629f
C444 plus.n29 a_n2158_n2088# 0.043629f
C445 plus.n30 a_n2158_n2088# 0.043629f
C446 plus.n31 a_n2158_n2088# 0.0099f
C447 plus.n32 a_n2158_n2088# 0.245601f
C448 plus.n33 a_n2158_n2088# 0.0099f
C449 plus.n34 a_n2158_n2088# 0.243584f
C450 plus.n35 a_n2158_n2088# 1.20211f
.ends

