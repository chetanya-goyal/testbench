* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t11 minus.t0 drain_right.t4 a_n1236_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X1 source.t4 plus.t0 drain_left.t5 a_n1236_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X2 a_n1236_n1488# a_n1236_n1488# a_n1236_n1488# a_n1236_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=11.4 ps=55.6 w=3 l=0.15
X3 drain_left.t4 plus.t1 source.t5 a_n1236_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X4 a_n1236_n1488# a_n1236_n1488# a_n1236_n1488# a_n1236_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X5 a_n1236_n1488# a_n1236_n1488# a_n1236_n1488# a_n1236_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X6 drain_right.t5 minus.t1 source.t10 a_n1236_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X7 source.t9 minus.t2 drain_right.t1 a_n1236_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X8 drain_right.t2 minus.t3 source.t8 a_n1236_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X9 drain_left.t3 plus.t2 source.t3 a_n1236_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X10 drain_left.t2 plus.t3 source.t2 a_n1236_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X11 drain_right.t0 minus.t4 source.t7 a_n1236_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X12 drain_left.t1 plus.t4 source.t1 a_n1236_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X13 source.t0 plus.t5 drain_left.t0 a_n1236_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X14 drain_right.t3 minus.t5 source.t6 a_n1236_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X15 a_n1236_n1488# a_n1236_n1488# a_n1236_n1488# a_n1236_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
R0 minus.n2 minus.t4 749.292
R1 minus.n0 minus.t3 749.292
R2 minus.n6 minus.t5 749.292
R3 minus.n4 minus.t1 749.292
R4 minus.n1 minus.t2 690.867
R5 minus.n5 minus.t0 690.867
R6 minus.n3 minus.n0 161.489
R7 minus.n7 minus.n4 161.489
R8 minus.n3 minus.n2 161.3
R9 minus.n7 minus.n6 161.3
R10 minus.n2 minus.n1 36.5157
R11 minus.n1 minus.n0 36.5157
R12 minus.n5 minus.n4 36.5157
R13 minus.n6 minus.n5 36.5157
R14 minus.n8 minus.n3 27.0365
R15 minus.n8 minus.n7 6.55164
R16 minus minus.n8 0.188
R17 drain_right.n1 drain_right.t5 90.1379
R18 drain_right.n3 drain_right.t0 89.7731
R19 drain_right.n3 drain_right.n2 80.3335
R20 drain_right.n1 drain_right.n0 79.8577
R21 drain_right drain_right.n1 21.5366
R22 drain_right.n0 drain_right.t4 10.0005
R23 drain_right.n0 drain_right.t3 10.0005
R24 drain_right.n2 drain_right.t1 10.0005
R25 drain_right.n2 drain_right.t2 10.0005
R26 drain_right drain_right.n3 5.93339
R27 source.n0 source.t1 73.0943
R28 source.n3 source.t8 73.0943
R29 source.n11 source.t6 73.0942
R30 source.n8 source.t5 73.0942
R31 source.n2 source.n1 63.0943
R32 source.n5 source.n4 63.0943
R33 source.n10 source.n9 63.0942
R34 source.n7 source.n6 63.0942
R35 source.n7 source.n5 15.5902
R36 source.n9 source.t10 10.0005
R37 source.n9 source.t11 10.0005
R38 source.n6 source.t3 10.0005
R39 source.n6 source.t4 10.0005
R40 source.n1 source.t2 10.0005
R41 source.n1 source.t0 10.0005
R42 source.n4 source.t7 10.0005
R43 source.n4 source.t9 10.0005
R44 source.n12 source.n0 9.48679
R45 source.n12 source.n11 5.5436
R46 source.n3 source.n2 0.7505
R47 source.n10 source.n8 0.7505
R48 source.n5 source.n3 0.560845
R49 source.n2 source.n0 0.560845
R50 source.n8 source.n7 0.560845
R51 source.n11 source.n10 0.560845
R52 source source.n12 0.188
R53 plus.n0 plus.t3 749.292
R54 plus.n2 plus.t4 749.292
R55 plus.n4 plus.t1 749.292
R56 plus.n6 plus.t2 749.292
R57 plus.n1 plus.t5 690.867
R58 plus.n5 plus.t0 690.867
R59 plus.n3 plus.n0 161.489
R60 plus.n7 plus.n4 161.489
R61 plus.n3 plus.n2 161.3
R62 plus.n7 plus.n6 161.3
R63 plus.n1 plus.n0 36.5157
R64 plus.n2 plus.n1 36.5157
R65 plus.n6 plus.n5 36.5157
R66 plus.n5 plus.n4 36.5157
R67 plus plus.n7 24.3267
R68 plus plus.n3 8.78648
R69 drain_left.n3 drain_left.t2 90.3335
R70 drain_left.n1 drain_left.t3 90.1379
R71 drain_left.n1 drain_left.n0 79.8577
R72 drain_left.n3 drain_left.n2 79.7731
R73 drain_left drain_left.n1 22.0898
R74 drain_left.n0 drain_left.t5 10.0005
R75 drain_left.n0 drain_left.t4 10.0005
R76 drain_left.n2 drain_left.t0 10.0005
R77 drain_left.n2 drain_left.t1 10.0005
R78 drain_left drain_left.n3 6.21356
C0 minus drain_right 0.687345f
C1 minus source 0.624644f
C2 drain_left plus 0.802509f
C3 drain_left drain_right 0.572274f
C4 drain_left source 4.84361f
C5 drain_right plus 0.274993f
C6 minus drain_left 0.175499f
C7 source plus 0.638804f
C8 minus plus 3.01468f
C9 source drain_right 4.83941f
C10 drain_right a_n1236_n1488# 3.33018f
C11 drain_left a_n1236_n1488# 3.48846f
C12 source a_n1236_n1488# 2.746948f
C13 minus a_n1236_n1488# 3.80918f
C14 plus a_n1236_n1488# 4.71289f
C15 drain_left.t3 a_n1236_n1488# 0.48338f
C16 drain_left.t5 a_n1236_n1488# 0.073703f
C17 drain_left.t4 a_n1236_n1488# 0.073703f
C18 drain_left.n0 a_n1236_n1488# 0.401169f
C19 drain_left.n1 a_n1236_n1488# 0.964022f
C20 drain_left.t2 a_n1236_n1488# 0.483991f
C21 drain_left.t0 a_n1236_n1488# 0.073703f
C22 drain_left.t1 a_n1236_n1488# 0.073703f
C23 drain_left.n2 a_n1236_n1488# 0.400937f
C24 drain_left.n3 a_n1236_n1488# 0.668875f
C25 plus.t3 a_n1236_n1488# 0.057791f
C26 plus.n0 a_n1236_n1488# 0.054321f
C27 plus.t5 a_n1236_n1488# 0.054709f
C28 plus.n1 a_n1236_n1488# 0.038237f
C29 plus.t4 a_n1236_n1488# 0.057791f
C30 plus.n2 a_n1236_n1488# 0.054258f
C31 plus.n3 a_n1236_n1488# 0.372531f
C32 plus.t1 a_n1236_n1488# 0.057791f
C33 plus.n4 a_n1236_n1488# 0.054321f
C34 plus.t2 a_n1236_n1488# 0.057791f
C35 plus.t0 a_n1236_n1488# 0.054709f
C36 plus.n5 a_n1236_n1488# 0.038237f
C37 plus.n6 a_n1236_n1488# 0.054258f
C38 plus.n7 a_n1236_n1488# 0.916902f
C39 source.t1 a_n1236_n1488# 0.514876f
C40 source.n0 a_n1236_n1488# 0.679701f
C41 source.t2 a_n1236_n1488# 0.087419f
C42 source.t0 a_n1236_n1488# 0.087419f
C43 source.n1 a_n1236_n1488# 0.425272f
C44 source.n2 a_n1236_n1488# 0.314767f
C45 source.t8 a_n1236_n1488# 0.514876f
C46 source.n3 a_n1236_n1488# 0.382516f
C47 source.t7 a_n1236_n1488# 0.087419f
C48 source.t9 a_n1236_n1488# 0.087419f
C49 source.n4 a_n1236_n1488# 0.425272f
C50 source.n5 a_n1236_n1488# 0.909901f
C51 source.t3 a_n1236_n1488# 0.087419f
C52 source.t4 a_n1236_n1488# 0.087419f
C53 source.n6 a_n1236_n1488# 0.425269f
C54 source.n7 a_n1236_n1488# 0.909903f
C55 source.t5 a_n1236_n1488# 0.514873f
C56 source.n8 a_n1236_n1488# 0.382519f
C57 source.t10 a_n1236_n1488# 0.087419f
C58 source.t11 a_n1236_n1488# 0.087419f
C59 source.n9 a_n1236_n1488# 0.425269f
C60 source.n10 a_n1236_n1488# 0.314769f
C61 source.t6 a_n1236_n1488# 0.514873f
C62 source.n11 a_n1236_n1488# 0.499012f
C63 source.n12 a_n1236_n1488# 0.706016f
C64 drain_right.t5 a_n1236_n1488# 0.491601f
C65 drain_right.t4 a_n1236_n1488# 0.074957f
C66 drain_right.t3 a_n1236_n1488# 0.074957f
C67 drain_right.n0 a_n1236_n1488# 0.407992f
C68 drain_right.n1 a_n1236_n1488# 0.938739f
C69 drain_right.t1 a_n1236_n1488# 0.074957f
C70 drain_right.t2 a_n1236_n1488# 0.074957f
C71 drain_right.n2 a_n1236_n1488# 0.409505f
C72 drain_right.t0 a_n1236_n1488# 0.490577f
C73 drain_right.n3 a_n1236_n1488# 0.689266f
C74 minus.t3 a_n1236_n1488# 0.056201f
C75 minus.n0 a_n1236_n1488# 0.052826f
C76 minus.t4 a_n1236_n1488# 0.056201f
C77 minus.t2 a_n1236_n1488# 0.053203f
C78 minus.n1 a_n1236_n1488# 0.037185f
C79 minus.n2 a_n1236_n1488# 0.052765f
C80 minus.n3 a_n1236_n1488# 0.939142f
C81 minus.t1 a_n1236_n1488# 0.056201f
C82 minus.n4 a_n1236_n1488# 0.052826f
C83 minus.t0 a_n1236_n1488# 0.053203f
C84 minus.n5 a_n1236_n1488# 0.037185f
C85 minus.t5 a_n1236_n1488# 0.056201f
C86 minus.n6 a_n1236_n1488# 0.052765f
C87 minus.n7 a_n1236_n1488# 0.323961f
C88 minus.n8 a_n1236_n1488# 1.09332f
.ends

