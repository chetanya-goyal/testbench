* NGSPICE file created from diffpair235.ext - technology: sky130A

.subckt diffpair235 minus drain_right drain_left source plus
X0 source.t22 minus.t0 drain_right.t2 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X1 drain_left.t11 plus.t0 source.t2 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X2 source.t21 minus.t1 drain_right.t10 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X3 source.t20 minus.t2 drain_right.t9 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X4 a_n2298_n1488# a_n2298_n1488# a_n2298_n1488# a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.8
X5 a_n2298_n1488# a_n2298_n1488# a_n2298_n1488# a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X6 drain_left.t10 plus.t1 source.t4 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X7 drain_left.t9 plus.t2 source.t9 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X8 a_n2298_n1488# a_n2298_n1488# a_n2298_n1488# a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X9 a_n2298_n1488# a_n2298_n1488# a_n2298_n1488# a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X10 drain_right.t8 minus.t3 source.t19 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X11 drain_right.t7 minus.t4 source.t18 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X12 source.t17 minus.t5 drain_right.t3 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X13 drain_right.t4 minus.t6 source.t16 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X14 drain_right.t11 minus.t7 source.t15 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X15 source.t14 minus.t8 drain_right.t0 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X16 drain_right.t5 minus.t9 source.t13 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X17 source.t10 plus.t3 drain_left.t8 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X18 source.t12 minus.t10 drain_right.t1 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X19 source.t0 plus.t4 drain_left.t7 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X20 source.t23 plus.t5 drain_left.t6 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X21 drain_right.t6 minus.t11 source.t11 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X22 drain_left.t5 plus.t6 source.t1 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X23 drain_left.t4 plus.t7 source.t6 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X24 source.t5 plus.t8 drain_left.t3 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X25 source.t3 plus.t9 drain_left.t2 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X26 drain_left.t1 plus.t10 source.t8 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X27 source.t7 plus.t11 drain_left.t0 a_n2298_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
R0 minus.n15 minus.n14 161.3
R1 minus.n13 minus.n0 161.3
R2 minus.n12 minus.n11 161.3
R3 minus.n10 minus.n1 161.3
R4 minus.n6 minus.n5 161.3
R5 minus.n31 minus.n30 161.3
R6 minus.n29 minus.n16 161.3
R7 minus.n28 minus.n27 161.3
R8 minus.n26 minus.n17 161.3
R9 minus.n22 minus.n21 161.3
R10 minus.n4 minus.t7 160.875
R11 minus.n20 minus.t1 160.875
R12 minus.n3 minus.t5 139.48
R13 minus.n7 minus.t3 139.48
R14 minus.n8 minus.t10 139.48
R15 minus.n12 minus.t11 139.48
R16 minus.n14 minus.t8 139.48
R17 minus.n19 minus.t4 139.48
R18 minus.n23 minus.t2 139.48
R19 minus.n24 minus.t6 139.48
R20 minus.n28 minus.t0 139.48
R21 minus.n30 minus.t9 139.48
R22 minus.n9 minus.n8 80.6037
R23 minus.n7 minus.n2 80.6037
R24 minus.n25 minus.n24 80.6037
R25 minus.n23 minus.n18 80.6037
R26 minus.n8 minus.n7 48.2005
R27 minus.n24 minus.n23 48.2005
R28 minus.n5 minus.n4 44.853
R29 minus.n21 minus.n20 44.853
R30 minus.n7 minus.n6 41.6278
R31 minus.n8 minus.n1 41.6278
R32 minus.n23 minus.n22 41.6278
R33 minus.n24 minus.n17 41.6278
R34 minus.n32 minus.n15 31.2088
R35 minus.n14 minus.n13 25.5611
R36 minus.n30 minus.n29 25.5611
R37 minus.n13 minus.n12 22.6399
R38 minus.n29 minus.n28 22.6399
R39 minus.n4 minus.n3 20.5405
R40 minus.n20 minus.n19 20.5405
R41 minus.n32 minus.n31 6.70126
R42 minus.n6 minus.n3 6.57323
R43 minus.n12 minus.n1 6.57323
R44 minus.n22 minus.n19 6.57323
R45 minus.n28 minus.n17 6.57323
R46 minus.n9 minus.n2 0.380177
R47 minus.n25 minus.n18 0.380177
R48 minus.n10 minus.n9 0.285035
R49 minus.n5 minus.n2 0.285035
R50 minus.n21 minus.n18 0.285035
R51 minus.n26 minus.n25 0.285035
R52 minus.n15 minus.n0 0.189894
R53 minus.n11 minus.n0 0.189894
R54 minus.n11 minus.n10 0.189894
R55 minus.n27 minus.n26 0.189894
R56 minus.n27 minus.n16 0.189894
R57 minus.n31 minus.n16 0.189894
R58 minus minus.n32 0.188
R59 drain_right.n6 drain_right.n4 80.7472
R60 drain_right.n3 drain_right.n2 80.6918
R61 drain_right.n3 drain_right.n0 80.6918
R62 drain_right.n6 drain_right.n5 79.7731
R63 drain_right.n8 drain_right.n7 79.7731
R64 drain_right.n3 drain_right.n1 79.773
R65 drain_right drain_right.n3 24.8664
R66 drain_right drain_right.n8 6.62735
R67 drain_right.n1 drain_right.t9 6.6005
R68 drain_right.n1 drain_right.t4 6.6005
R69 drain_right.n2 drain_right.t2 6.6005
R70 drain_right.n2 drain_right.t5 6.6005
R71 drain_right.n0 drain_right.t10 6.6005
R72 drain_right.n0 drain_right.t7 6.6005
R73 drain_right.n4 drain_right.t3 6.6005
R74 drain_right.n4 drain_right.t11 6.6005
R75 drain_right.n5 drain_right.t1 6.6005
R76 drain_right.n5 drain_right.t8 6.6005
R77 drain_right.n7 drain_right.t0 6.6005
R78 drain_right.n7 drain_right.t6 6.6005
R79 drain_right.n8 drain_right.n6 0.974638
R80 source.n0 source.t1 69.6943
R81 source.n5 source.t7 69.6943
R82 source.n6 source.t15 69.6943
R83 source.n11 source.t14 69.6943
R84 source.n23 source.t13 69.6942
R85 source.n18 source.t21 69.6942
R86 source.n17 source.t4 69.6942
R87 source.n12 source.t23 69.6942
R88 source.n2 source.n1 63.0943
R89 source.n4 source.n3 63.0943
R90 source.n8 source.n7 63.0943
R91 source.n10 source.n9 63.0943
R92 source.n22 source.n21 63.0942
R93 source.n20 source.n19 63.0942
R94 source.n16 source.n15 63.0942
R95 source.n14 source.n13 63.0942
R96 source.n12 source.n11 15.4437
R97 source.n24 source.n0 9.69368
R98 source.n21 source.t16 6.6005
R99 source.n21 source.t22 6.6005
R100 source.n19 source.t18 6.6005
R101 source.n19 source.t20 6.6005
R102 source.n15 source.t9 6.6005
R103 source.n15 source.t10 6.6005
R104 source.n13 source.t2 6.6005
R105 source.n13 source.t0 6.6005
R106 source.n1 source.t6 6.6005
R107 source.n1 source.t3 6.6005
R108 source.n3 source.t8 6.6005
R109 source.n3 source.t5 6.6005
R110 source.n7 source.t19 6.6005
R111 source.n7 source.t17 6.6005
R112 source.n9 source.t11 6.6005
R113 source.n9 source.t12 6.6005
R114 source.n24 source.n23 5.7505
R115 source.n11 source.n10 0.974638
R116 source.n10 source.n8 0.974638
R117 source.n8 source.n6 0.974638
R118 source.n5 source.n4 0.974638
R119 source.n4 source.n2 0.974638
R120 source.n2 source.n0 0.974638
R121 source.n14 source.n12 0.974638
R122 source.n16 source.n14 0.974638
R123 source.n17 source.n16 0.974638
R124 source.n20 source.n18 0.974638
R125 source.n22 source.n20 0.974638
R126 source.n23 source.n22 0.974638
R127 source.n6 source.n5 0.470328
R128 source.n18 source.n17 0.470328
R129 source source.n24 0.188
R130 plus.n6 plus.n3 161.3
R131 plus.n11 plus.n10 161.3
R132 plus.n12 plus.n1 161.3
R133 plus.n13 plus.n0 161.3
R134 plus.n15 plus.n14 161.3
R135 plus.n22 plus.n19 161.3
R136 plus.n27 plus.n26 161.3
R137 plus.n28 plus.n17 161.3
R138 plus.n29 plus.n16 161.3
R139 plus.n31 plus.n30 161.3
R140 plus.n4 plus.t11 160.875
R141 plus.n20 plus.t1 160.875
R142 plus.n14 plus.t6 139.48
R143 plus.n12 plus.t9 139.48
R144 plus.n2 plus.t7 139.48
R145 plus.n7 plus.t8 139.48
R146 plus.n5 plus.t10 139.48
R147 plus.n30 plus.t5 139.48
R148 plus.n28 plus.t0 139.48
R149 plus.n18 plus.t4 139.48
R150 plus.n23 plus.t2 139.48
R151 plus.n21 plus.t3 139.48
R152 plus.n8 plus.n7 80.6037
R153 plus.n9 plus.n2 80.6037
R154 plus.n24 plus.n23 80.6037
R155 plus.n25 plus.n18 80.6037
R156 plus.n7 plus.n2 48.2005
R157 plus.n23 plus.n18 48.2005
R158 plus.n4 plus.n3 44.853
R159 plus.n20 plus.n19 44.853
R160 plus.n11 plus.n2 41.6278
R161 plus.n7 plus.n6 41.6278
R162 plus.n27 plus.n18 41.6278
R163 plus.n23 plus.n22 41.6278
R164 plus plus.n31 28.499
R165 plus.n14 plus.n13 25.5611
R166 plus.n30 plus.n29 25.5611
R167 plus.n13 plus.n12 22.6399
R168 plus.n29 plus.n28 22.6399
R169 plus.n5 plus.n4 20.5405
R170 plus.n21 plus.n20 20.5405
R171 plus plus.n15 8.93611
R172 plus.n12 plus.n11 6.57323
R173 plus.n6 plus.n5 6.57323
R174 plus.n28 plus.n27 6.57323
R175 plus.n22 plus.n21 6.57323
R176 plus.n9 plus.n8 0.380177
R177 plus.n25 plus.n24 0.380177
R178 plus.n8 plus.n3 0.285035
R179 plus.n10 plus.n9 0.285035
R180 plus.n26 plus.n25 0.285035
R181 plus.n24 plus.n19 0.285035
R182 plus.n10 plus.n1 0.189894
R183 plus.n1 plus.n0 0.189894
R184 plus.n15 plus.n0 0.189894
R185 plus.n31 plus.n16 0.189894
R186 plus.n17 plus.n16 0.189894
R187 plus.n26 plus.n17 0.189894
R188 drain_left.n6 drain_left.n4 80.7472
R189 drain_left.n3 drain_left.n2 80.6918
R190 drain_left.n3 drain_left.n0 80.6918
R191 drain_left.n8 drain_left.n7 79.7731
R192 drain_left.n6 drain_left.n5 79.7731
R193 drain_left.n3 drain_left.n1 79.773
R194 drain_left drain_left.n3 25.4196
R195 drain_left drain_left.n8 6.62735
R196 drain_left.n1 drain_left.t7 6.6005
R197 drain_left.n1 drain_left.t9 6.6005
R198 drain_left.n2 drain_left.t8 6.6005
R199 drain_left.n2 drain_left.t10 6.6005
R200 drain_left.n0 drain_left.t6 6.6005
R201 drain_left.n0 drain_left.t11 6.6005
R202 drain_left.n7 drain_left.t2 6.6005
R203 drain_left.n7 drain_left.t5 6.6005
R204 drain_left.n5 drain_left.t3 6.6005
R205 drain_left.n5 drain_left.t4 6.6005
R206 drain_left.n4 drain_left.t0 6.6005
R207 drain_left.n4 drain_left.t1 6.6005
R208 drain_left.n8 drain_left.n6 0.974638
C0 source plus 2.92517f
C1 minus drain_right 2.49097f
C2 drain_left drain_right 1.16188f
C3 minus source 2.91117f
C4 minus plus 4.34547f
C5 source drain_left 5.85299f
C6 drain_left plus 2.71722f
C7 source drain_right 5.85554f
C8 drain_right plus 0.387413f
C9 minus drain_left 0.177211f
C10 drain_right a_n2298_n1488# 4.57488f
C11 drain_left a_n2298_n1488# 4.91004f
C12 source a_n2298_n1488# 3.873853f
C13 minus a_n2298_n1488# 8.33217f
C14 plus a_n2298_n1488# 9.57858f
C15 drain_left.t6 a_n2298_n1488# 0.062706f
C16 drain_left.t11 a_n2298_n1488# 0.062706f
C17 drain_left.n0 a_n2298_n1488# 0.456602f
C18 drain_left.t7 a_n2298_n1488# 0.062706f
C19 drain_left.t9 a_n2298_n1488# 0.062706f
C20 drain_left.n1 a_n2298_n1488# 0.452225f
C21 drain_left.t8 a_n2298_n1488# 0.062706f
C22 drain_left.t10 a_n2298_n1488# 0.062706f
C23 drain_left.n2 a_n2298_n1488# 0.456602f
C24 drain_left.n3 a_n2298_n1488# 2.00662f
C25 drain_left.t0 a_n2298_n1488# 0.062706f
C26 drain_left.t1 a_n2298_n1488# 0.062706f
C27 drain_left.n4 a_n2298_n1488# 0.456914f
C28 drain_left.t3 a_n2298_n1488# 0.062706f
C29 drain_left.t4 a_n2298_n1488# 0.062706f
C30 drain_left.n5 a_n2298_n1488# 0.452228f
C31 drain_left.n6 a_n2298_n1488# 0.761523f
C32 drain_left.t2 a_n2298_n1488# 0.062706f
C33 drain_left.t5 a_n2298_n1488# 0.062706f
C34 drain_left.n7 a_n2298_n1488# 0.452228f
C35 drain_left.n8 a_n2298_n1488# 0.614956f
C36 plus.n0 a_n2298_n1488# 0.043258f
C37 plus.t6 a_n2298_n1488# 0.311318f
C38 plus.t9 a_n2298_n1488# 0.311318f
C39 plus.n1 a_n2298_n1488# 0.043258f
C40 plus.t7 a_n2298_n1488# 0.311318f
C41 plus.n2 a_n2298_n1488# 0.189447f
C42 plus.n3 a_n2298_n1488# 0.198588f
C43 plus.t8 a_n2298_n1488# 0.311318f
C44 plus.t10 a_n2298_n1488# 0.311318f
C45 plus.t11 a_n2298_n1488# 0.335225f
C46 plus.n4 a_n2298_n1488# 0.160148f
C47 plus.n5 a_n2298_n1488# 0.180734f
C48 plus.n6 a_n2298_n1488# 0.009816f
C49 plus.n7 a_n2298_n1488# 0.189447f
C50 plus.n8 a_n2298_n1488# 0.072052f
C51 plus.n9 a_n2298_n1488# 0.072052f
C52 plus.n10 a_n2298_n1488# 0.057723f
C53 plus.n11 a_n2298_n1488# 0.009816f
C54 plus.n12 a_n2298_n1488# 0.177364f
C55 plus.n13 a_n2298_n1488# 0.009816f
C56 plus.n14 a_n2298_n1488# 0.176697f
C57 plus.n15 a_n2298_n1488# 0.344552f
C58 plus.n16 a_n2298_n1488# 0.043258f
C59 plus.t5 a_n2298_n1488# 0.311318f
C60 plus.n17 a_n2298_n1488# 0.043258f
C61 plus.t0 a_n2298_n1488# 0.311318f
C62 plus.t4 a_n2298_n1488# 0.311318f
C63 plus.n18 a_n2298_n1488# 0.189447f
C64 plus.n19 a_n2298_n1488# 0.198588f
C65 plus.t2 a_n2298_n1488# 0.311318f
C66 plus.t1 a_n2298_n1488# 0.335225f
C67 plus.n20 a_n2298_n1488# 0.160148f
C68 plus.t3 a_n2298_n1488# 0.311318f
C69 plus.n21 a_n2298_n1488# 0.180734f
C70 plus.n22 a_n2298_n1488# 0.009816f
C71 plus.n23 a_n2298_n1488# 0.189447f
C72 plus.n24 a_n2298_n1488# 0.072052f
C73 plus.n25 a_n2298_n1488# 0.072052f
C74 plus.n26 a_n2298_n1488# 0.057723f
C75 plus.n27 a_n2298_n1488# 0.009816f
C76 plus.n28 a_n2298_n1488# 0.177364f
C77 plus.n29 a_n2298_n1488# 0.009816f
C78 plus.n30 a_n2298_n1488# 0.176697f
C79 plus.n31 a_n2298_n1488# 1.1378f
C80 source.t1 a_n2298_n1488# 0.525818f
C81 source.n0 a_n2298_n1488# 0.782514f
C82 source.t6 a_n2298_n1488# 0.063322f
C83 source.t3 a_n2298_n1488# 0.063322f
C84 source.n1 a_n2298_n1488# 0.401501f
C85 source.n2 a_n2298_n1488# 0.400366f
C86 source.t8 a_n2298_n1488# 0.063322f
C87 source.t5 a_n2298_n1488# 0.063322f
C88 source.n3 a_n2298_n1488# 0.401501f
C89 source.n4 a_n2298_n1488# 0.400366f
C90 source.t7 a_n2298_n1488# 0.525818f
C91 source.n5 a_n2298_n1488# 0.405341f
C92 source.t15 a_n2298_n1488# 0.525818f
C93 source.n6 a_n2298_n1488# 0.405341f
C94 source.t19 a_n2298_n1488# 0.063322f
C95 source.t17 a_n2298_n1488# 0.063322f
C96 source.n7 a_n2298_n1488# 0.401501f
C97 source.n8 a_n2298_n1488# 0.400366f
C98 source.t11 a_n2298_n1488# 0.063322f
C99 source.t12 a_n2298_n1488# 0.063322f
C100 source.n9 a_n2298_n1488# 0.401501f
C101 source.n10 a_n2298_n1488# 0.400366f
C102 source.t14 a_n2298_n1488# 0.525818f
C103 source.n11 a_n2298_n1488# 1.07001f
C104 source.t23 a_n2298_n1488# 0.525815f
C105 source.n12 a_n2298_n1488# 1.07001f
C106 source.t2 a_n2298_n1488# 0.063322f
C107 source.t0 a_n2298_n1488# 0.063322f
C108 source.n13 a_n2298_n1488# 0.401498f
C109 source.n14 a_n2298_n1488# 0.400369f
C110 source.t9 a_n2298_n1488# 0.063322f
C111 source.t10 a_n2298_n1488# 0.063322f
C112 source.n15 a_n2298_n1488# 0.401498f
C113 source.n16 a_n2298_n1488# 0.400369f
C114 source.t4 a_n2298_n1488# 0.525815f
C115 source.n17 a_n2298_n1488# 0.405344f
C116 source.t21 a_n2298_n1488# 0.525815f
C117 source.n18 a_n2298_n1488# 0.405344f
C118 source.t18 a_n2298_n1488# 0.063322f
C119 source.t20 a_n2298_n1488# 0.063322f
C120 source.n19 a_n2298_n1488# 0.401498f
C121 source.n20 a_n2298_n1488# 0.400369f
C122 source.t16 a_n2298_n1488# 0.063322f
C123 source.t22 a_n2298_n1488# 0.063322f
C124 source.n21 a_n2298_n1488# 0.401498f
C125 source.n22 a_n2298_n1488# 0.400369f
C126 source.t13 a_n2298_n1488# 0.525815f
C127 source.n23 a_n2298_n1488# 0.58536f
C128 source.n24 a_n2298_n1488# 0.791146f
C129 drain_right.t10 a_n2298_n1488# 0.061993f
C130 drain_right.t7 a_n2298_n1488# 0.061993f
C131 drain_right.n0 a_n2298_n1488# 0.451415f
C132 drain_right.t9 a_n2298_n1488# 0.061993f
C133 drain_right.t4 a_n2298_n1488# 0.061993f
C134 drain_right.n1 a_n2298_n1488# 0.447088f
C135 drain_right.t2 a_n2298_n1488# 0.061993f
C136 drain_right.t5 a_n2298_n1488# 0.061993f
C137 drain_right.n2 a_n2298_n1488# 0.451415f
C138 drain_right.n3 a_n2298_n1488# 1.93228f
C139 drain_right.t3 a_n2298_n1488# 0.061993f
C140 drain_right.t11 a_n2298_n1488# 0.061993f
C141 drain_right.n4 a_n2298_n1488# 0.451723f
C142 drain_right.t1 a_n2298_n1488# 0.061993f
C143 drain_right.t8 a_n2298_n1488# 0.061993f
C144 drain_right.n5 a_n2298_n1488# 0.44709f
C145 drain_right.n6 a_n2298_n1488# 0.752871f
C146 drain_right.t0 a_n2298_n1488# 0.061993f
C147 drain_right.t6 a_n2298_n1488# 0.061993f
C148 drain_right.n7 a_n2298_n1488# 0.44709f
C149 drain_right.n8 a_n2298_n1488# 0.607969f
C150 minus.n0 a_n2298_n1488# 0.042013f
C151 minus.n1 a_n2298_n1488# 0.009534f
C152 minus.t11 a_n2298_n1488# 0.302357f
C153 minus.n2 a_n2298_n1488# 0.069978f
C154 minus.t5 a_n2298_n1488# 0.302357f
C155 minus.n3 a_n2298_n1488# 0.175532f
C156 minus.t7 a_n2298_n1488# 0.325576f
C157 minus.n4 a_n2298_n1488# 0.155538f
C158 minus.n5 a_n2298_n1488# 0.192872f
C159 minus.n6 a_n2298_n1488# 0.009534f
C160 minus.t3 a_n2298_n1488# 0.302357f
C161 minus.n7 a_n2298_n1488# 0.183994f
C162 minus.t10 a_n2298_n1488# 0.302357f
C163 minus.n8 a_n2298_n1488# 0.183994f
C164 minus.n9 a_n2298_n1488# 0.069978f
C165 minus.n10 a_n2298_n1488# 0.056061f
C166 minus.n11 a_n2298_n1488# 0.042013f
C167 minus.n12 a_n2298_n1488# 0.172259f
C168 minus.n13 a_n2298_n1488# 0.009534f
C169 minus.t8 a_n2298_n1488# 0.302357f
C170 minus.n14 a_n2298_n1488# 0.171611f
C171 minus.n15 a_n2298_n1488# 1.17599f
C172 minus.n16 a_n2298_n1488# 0.042013f
C173 minus.n17 a_n2298_n1488# 0.009534f
C174 minus.n18 a_n2298_n1488# 0.069978f
C175 minus.t4 a_n2298_n1488# 0.302357f
C176 minus.n19 a_n2298_n1488# 0.175532f
C177 minus.t1 a_n2298_n1488# 0.325576f
C178 minus.n20 a_n2298_n1488# 0.155538f
C179 minus.n21 a_n2298_n1488# 0.192872f
C180 minus.n22 a_n2298_n1488# 0.009534f
C181 minus.t2 a_n2298_n1488# 0.302357f
C182 minus.n23 a_n2298_n1488# 0.183994f
C183 minus.t6 a_n2298_n1488# 0.302357f
C184 minus.n24 a_n2298_n1488# 0.183994f
C185 minus.n25 a_n2298_n1488# 0.069978f
C186 minus.n26 a_n2298_n1488# 0.056061f
C187 minus.n27 a_n2298_n1488# 0.042013f
C188 minus.t0 a_n2298_n1488# 0.302357f
C189 minus.n28 a_n2298_n1488# 0.172259f
C190 minus.n29 a_n2298_n1488# 0.009534f
C191 minus.t9 a_n2298_n1488# 0.302357f
C192 minus.n30 a_n2298_n1488# 0.171611f
C193 minus.n31 a_n2298_n1488# 0.294406f
C194 minus.n32 a_n2298_n1488# 1.4384f
.ends

