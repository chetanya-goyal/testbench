* NGSPICE file created from diffpair196.ext - technology: sky130A

.subckt diffpair196 minus drain_right drain_left source plus
X0 source.t27 minus.t0 drain_right.t7 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X1 source.t26 minus.t1 drain_right.t1 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X2 source.t25 minus.t2 drain_right.t8 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X3 drain_left.t13 plus.t0 source.t11 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X4 drain_right.t2 minus.t3 source.t24 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X5 drain_right.t3 minus.t4 source.t23 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X6 drain_left.t12 plus.t1 source.t1 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X7 drain_left.t11 plus.t2 source.t10 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X8 drain_right.t0 minus.t5 source.t22 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X9 a_n1724_n1488# a_n1724_n1488# a_n1724_n1488# a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.3
X10 drain_right.t4 minus.t6 source.t21 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X11 drain_left.t10 plus.t3 source.t2 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X12 source.t5 plus.t4 drain_left.t9 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X13 source.t13 plus.t5 drain_left.t8 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X14 source.t20 minus.t7 drain_right.t9 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X15 source.t19 minus.t8 drain_right.t11 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X16 drain_left.t7 plus.t6 source.t7 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X17 a_n1724_n1488# a_n1724_n1488# a_n1724_n1488# a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X18 drain_right.t12 minus.t9 source.t18 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X19 source.t9 plus.t7 drain_left.t6 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X20 drain_right.t13 minus.t10 source.t17 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X21 drain_left.t5 plus.t8 source.t4 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X22 a_n1724_n1488# a_n1724_n1488# a_n1724_n1488# a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X23 drain_left.t4 plus.t9 source.t6 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X24 drain_right.t5 minus.t11 source.t16 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X25 a_n1724_n1488# a_n1724_n1488# a_n1724_n1488# a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X26 source.t15 minus.t12 drain_right.t10 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X27 drain_right.t6 minus.t13 source.t14 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X28 source.t8 plus.t10 drain_left.t3 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X29 drain_left.t2 plus.t11 source.t3 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X30 source.t12 plus.t12 drain_left.t1 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X31 source.t0 plus.t13 drain_left.t0 a_n1724_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
R0 minus.n15 minus.t5 402.397
R1 minus.n3 minus.t9 402.397
R2 minus.n32 minus.t10 402.397
R3 minus.n20 minus.t6 402.397
R4 minus.n1 minus.t8 345.433
R5 minus.n14 minus.t1 345.433
R6 minus.n12 minus.t11 345.433
R7 minus.n6 minus.t3 345.433
R8 minus.n4 minus.t12 345.433
R9 minus.n18 minus.t7 345.433
R10 minus.n31 minus.t2 345.433
R11 minus.n29 minus.t4 345.433
R12 minus.n23 minus.t13 345.433
R13 minus.n21 minus.t0 345.433
R14 minus.n3 minus.n2 161.489
R15 minus.n20 minus.n19 161.489
R16 minus.n16 minus.n15 161.3
R17 minus.n13 minus.n0 161.3
R18 minus.n11 minus.n10 161.3
R19 minus.n9 minus.n1 161.3
R20 minus.n8 minus.n7 161.3
R21 minus.n5 minus.n2 161.3
R22 minus.n33 minus.n32 161.3
R23 minus.n30 minus.n17 161.3
R24 minus.n28 minus.n27 161.3
R25 minus.n26 minus.n18 161.3
R26 minus.n25 minus.n24 161.3
R27 minus.n22 minus.n19 161.3
R28 minus.n11 minus.n1 73.0308
R29 minus.n7 minus.n1 73.0308
R30 minus.n24 minus.n18 73.0308
R31 minus.n28 minus.n18 73.0308
R32 minus.n13 minus.n12 54.0429
R33 minus.n6 minus.n5 54.0429
R34 minus.n23 minus.n22 54.0429
R35 minus.n30 minus.n29 54.0429
R36 minus.n14 minus.n13 37.9763
R37 minus.n5 minus.n4 37.9763
R38 minus.n22 minus.n21 37.9763
R39 minus.n31 minus.n30 37.9763
R40 minus.n15 minus.n14 35.055
R41 minus.n4 minus.n3 35.055
R42 minus.n21 minus.n20 35.055
R43 minus.n32 minus.n31 35.055
R44 minus.n34 minus.n16 28.8698
R45 minus.n12 minus.n11 18.9884
R46 minus.n7 minus.n6 18.9884
R47 minus.n24 minus.n23 18.9884
R48 minus.n29 minus.n28 18.9884
R49 minus.n34 minus.n33 6.53648
R50 minus.n16 minus.n0 0.189894
R51 minus.n10 minus.n0 0.189894
R52 minus.n10 minus.n9 0.189894
R53 minus.n9 minus.n8 0.189894
R54 minus.n8 minus.n2 0.189894
R55 minus.n25 minus.n19 0.189894
R56 minus.n26 minus.n25 0.189894
R57 minus.n27 minus.n26 0.189894
R58 minus.n27 minus.n17 0.189894
R59 minus.n33 minus.n17 0.189894
R60 minus minus.n34 0.188
R61 drain_right.n1 drain_right.t4 86.9161
R62 drain_right.n11 drain_right.t0 86.3731
R63 drain_right.n8 drain_right.n6 80.3162
R64 drain_right.n4 drain_right.n2 80.3161
R65 drain_right.n8 drain_right.n7 79.7731
R66 drain_right.n10 drain_right.n9 79.7731
R67 drain_right.n4 drain_right.n3 79.773
R68 drain_right.n1 drain_right.n0 79.773
R69 drain_right drain_right.n5 23.1185
R70 drain_right.n2 drain_right.t8 6.6005
R71 drain_right.n2 drain_right.t13 6.6005
R72 drain_right.n3 drain_right.t9 6.6005
R73 drain_right.n3 drain_right.t3 6.6005
R74 drain_right.n0 drain_right.t7 6.6005
R75 drain_right.n0 drain_right.t6 6.6005
R76 drain_right.n6 drain_right.t10 6.6005
R77 drain_right.n6 drain_right.t12 6.6005
R78 drain_right.n7 drain_right.t11 6.6005
R79 drain_right.n7 drain_right.t2 6.6005
R80 drain_right.n9 drain_right.t1 6.6005
R81 drain_right.n9 drain_right.t5 6.6005
R82 drain_right drain_right.n11 5.92477
R83 drain_right.n11 drain_right.n10 0.543603
R84 drain_right.n10 drain_right.n8 0.543603
R85 drain_right.n5 drain_right.n1 0.352482
R86 drain_right.n5 drain_right.n4 0.0809298
R87 source.n0 source.t3 69.6943
R88 source.n7 source.t18 69.6943
R89 source.n27 source.t17 69.6942
R90 source.n20 source.t10 69.6942
R91 source.n2 source.n1 63.0943
R92 source.n4 source.n3 63.0943
R93 source.n6 source.n5 63.0943
R94 source.n9 source.n8 63.0943
R95 source.n11 source.n10 63.0943
R96 source.n13 source.n12 63.0943
R97 source.n26 source.n25 63.0942
R98 source.n24 source.n23 63.0942
R99 source.n22 source.n21 63.0942
R100 source.n19 source.n18 63.0942
R101 source.n17 source.n16 63.0942
R102 source.n15 source.n14 63.0942
R103 source.n15 source.n13 15.5558
R104 source.n28 source.n0 9.47816
R105 source.n25 source.t23 6.6005
R106 source.n25 source.t25 6.6005
R107 source.n23 source.t14 6.6005
R108 source.n23 source.t20 6.6005
R109 source.n21 source.t21 6.6005
R110 source.n21 source.t27 6.6005
R111 source.n18 source.t6 6.6005
R112 source.n18 source.t8 6.6005
R113 source.n16 source.t11 6.6005
R114 source.n16 source.t5 6.6005
R115 source.n14 source.t7 6.6005
R116 source.n14 source.t12 6.6005
R117 source.n1 source.t2 6.6005
R118 source.n1 source.t9 6.6005
R119 source.n3 source.t4 6.6005
R120 source.n3 source.t0 6.6005
R121 source.n5 source.t1 6.6005
R122 source.n5 source.t13 6.6005
R123 source.n8 source.t24 6.6005
R124 source.n8 source.t15 6.6005
R125 source.n10 source.t16 6.6005
R126 source.n10 source.t19 6.6005
R127 source.n12 source.t22 6.6005
R128 source.n12 source.t26 6.6005
R129 source.n28 source.n27 5.53498
R130 source.n7 source.n6 0.741879
R131 source.n22 source.n20 0.741879
R132 source.n13 source.n11 0.543603
R133 source.n11 source.n9 0.543603
R134 source.n9 source.n7 0.543603
R135 source.n6 source.n4 0.543603
R136 source.n4 source.n2 0.543603
R137 source.n2 source.n0 0.543603
R138 source.n17 source.n15 0.543603
R139 source.n19 source.n17 0.543603
R140 source.n20 source.n19 0.543603
R141 source.n24 source.n22 0.543603
R142 source.n26 source.n24 0.543603
R143 source.n27 source.n26 0.543603
R144 source source.n28 0.188
R145 plus.n3 plus.t1 402.397
R146 plus.n15 plus.t11 402.397
R147 plus.n20 plus.t2 402.397
R148 plus.n32 plus.t6 402.397
R149 plus.n1 plus.t13 345.433
R150 plus.n4 plus.t5 345.433
R151 plus.n6 plus.t8 345.433
R152 plus.n12 plus.t3 345.433
R153 plus.n14 plus.t7 345.433
R154 plus.n18 plus.t4 345.433
R155 plus.n21 plus.t10 345.433
R156 plus.n23 plus.t9 345.433
R157 plus.n29 plus.t0 345.433
R158 plus.n31 plus.t12 345.433
R159 plus.n3 plus.n2 161.489
R160 plus.n20 plus.n19 161.489
R161 plus.n5 plus.n2 161.3
R162 plus.n8 plus.n7 161.3
R163 plus.n9 plus.n1 161.3
R164 plus.n11 plus.n10 161.3
R165 plus.n13 plus.n0 161.3
R166 plus.n16 plus.n15 161.3
R167 plus.n22 plus.n19 161.3
R168 plus.n25 plus.n24 161.3
R169 plus.n26 plus.n18 161.3
R170 plus.n28 plus.n27 161.3
R171 plus.n30 plus.n17 161.3
R172 plus.n33 plus.n32 161.3
R173 plus.n7 plus.n1 73.0308
R174 plus.n11 plus.n1 73.0308
R175 plus.n28 plus.n18 73.0308
R176 plus.n24 plus.n18 73.0308
R177 plus.n6 plus.n5 54.0429
R178 plus.n13 plus.n12 54.0429
R179 plus.n30 plus.n29 54.0429
R180 plus.n23 plus.n22 54.0429
R181 plus.n5 plus.n4 37.9763
R182 plus.n14 plus.n13 37.9763
R183 plus.n31 plus.n30 37.9763
R184 plus.n22 plus.n21 37.9763
R185 plus.n4 plus.n3 35.055
R186 plus.n15 plus.n14 35.055
R187 plus.n32 plus.n31 35.055
R188 plus.n21 plus.n20 35.055
R189 plus plus.n33 26.16
R190 plus.n7 plus.n6 18.9884
R191 plus.n12 plus.n11 18.9884
R192 plus.n29 plus.n28 18.9884
R193 plus.n24 plus.n23 18.9884
R194 plus plus.n16 8.77133
R195 plus.n8 plus.n2 0.189894
R196 plus.n9 plus.n8 0.189894
R197 plus.n10 plus.n9 0.189894
R198 plus.n10 plus.n0 0.189894
R199 plus.n16 plus.n0 0.189894
R200 plus.n33 plus.n17 0.189894
R201 plus.n27 plus.n17 0.189894
R202 plus.n27 plus.n26 0.189894
R203 plus.n26 plus.n25 0.189894
R204 plus.n25 plus.n19 0.189894
R205 drain_left.n7 drain_left.t12 86.9162
R206 drain_left.n1 drain_left.t7 86.9161
R207 drain_left.n4 drain_left.n2 80.3161
R208 drain_left.n11 drain_left.n10 79.7731
R209 drain_left.n9 drain_left.n8 79.7731
R210 drain_left.n7 drain_left.n6 79.7731
R211 drain_left.n4 drain_left.n3 79.773
R212 drain_left.n1 drain_left.n0 79.773
R213 drain_left drain_left.n5 23.6717
R214 drain_left.n2 drain_left.t3 6.6005
R215 drain_left.n2 drain_left.t11 6.6005
R216 drain_left.n3 drain_left.t9 6.6005
R217 drain_left.n3 drain_left.t4 6.6005
R218 drain_left.n0 drain_left.t1 6.6005
R219 drain_left.n0 drain_left.t13 6.6005
R220 drain_left.n10 drain_left.t6 6.6005
R221 drain_left.n10 drain_left.t2 6.6005
R222 drain_left.n8 drain_left.t0 6.6005
R223 drain_left.n8 drain_left.t10 6.6005
R224 drain_left.n6 drain_left.t8 6.6005
R225 drain_left.n6 drain_left.t5 6.6005
R226 drain_left drain_left.n11 6.19632
R227 drain_left.n9 drain_left.n7 0.543603
R228 drain_left.n11 drain_left.n9 0.543603
R229 drain_left.n5 drain_left.n1 0.352482
R230 drain_left.n5 drain_left.n4 0.0809298
C0 drain_right minus 1.67375f
C1 drain_right plus 0.327429f
C2 plus minus 3.63915f
C3 drain_right drain_left 0.880081f
C4 drain_right source 8.98499f
C5 minus drain_left 0.176873f
C6 plus drain_left 1.83968f
C7 minus source 1.79971f
C8 plus source 1.81387f
C9 source drain_left 8.98819f
C10 drain_right a_n1724_n1488# 4.24607f
C11 drain_left a_n1724_n1488# 4.49434f
C12 source a_n1724_n1488# 2.915101f
C13 minus a_n1724_n1488# 5.979425f
C14 plus a_n1724_n1488# 6.572834f
C15 drain_left.t7 a_n1724_n1488# 0.546697f
C16 drain_left.t1 a_n1724_n1488# 0.058866f
C17 drain_left.t13 a_n1724_n1488# 0.058866f
C18 drain_left.n0 a_n1724_n1488# 0.424536f
C19 drain_left.n1 a_n1724_n1488# 0.562622f
C20 drain_left.t3 a_n1724_n1488# 0.058866f
C21 drain_left.t11 a_n1724_n1488# 0.058866f
C22 drain_left.n2 a_n1724_n1488# 0.426535f
C23 drain_left.t9 a_n1724_n1488# 0.058866f
C24 drain_left.t4 a_n1724_n1488# 0.058866f
C25 drain_left.n3 a_n1724_n1488# 0.424536f
C26 drain_left.n4 a_n1724_n1488# 0.549489f
C27 drain_left.n5 a_n1724_n1488# 0.717799f
C28 drain_left.t12 a_n1724_n1488# 0.546699f
C29 drain_left.t8 a_n1724_n1488# 0.058866f
C30 drain_left.t5 a_n1724_n1488# 0.058866f
C31 drain_left.n6 a_n1724_n1488# 0.424538f
C32 drain_left.n7 a_n1724_n1488# 0.576274f
C33 drain_left.t0 a_n1724_n1488# 0.058866f
C34 drain_left.t10 a_n1724_n1488# 0.058866f
C35 drain_left.n8 a_n1724_n1488# 0.424538f
C36 drain_left.n9 a_n1724_n1488# 0.285672f
C37 drain_left.t6 a_n1724_n1488# 0.058866f
C38 drain_left.t2 a_n1724_n1488# 0.058866f
C39 drain_left.n10 a_n1724_n1488# 0.424538f
C40 drain_left.n11 a_n1724_n1488# 0.492354f
C41 plus.n0 a_n1724_n1488# 0.026435f
C42 plus.t7 a_n1724_n1488# 0.068897f
C43 plus.t3 a_n1724_n1488# 0.068897f
C44 plus.t13 a_n1724_n1488# 0.068897f
C45 plus.n1 a_n1724_n1488# 0.048774f
C46 plus.n2 a_n1724_n1488# 0.062281f
C47 plus.t8 a_n1724_n1488# 0.068897f
C48 plus.t5 a_n1724_n1488# 0.068897f
C49 plus.t1 a_n1724_n1488# 0.074998f
C50 plus.n3 a_n1724_n1488# 0.04793f
C51 plus.n4 a_n1724_n1488# 0.040005f
C52 plus.n5 a_n1724_n1488# 0.010888f
C53 plus.n6 a_n1724_n1488# 0.040005f
C54 plus.n7 a_n1724_n1488# 0.010888f
C55 plus.n8 a_n1724_n1488# 0.026435f
C56 plus.n9 a_n1724_n1488# 0.026435f
C57 plus.n10 a_n1724_n1488# 0.026435f
C58 plus.n11 a_n1724_n1488# 0.010888f
C59 plus.n12 a_n1724_n1488# 0.040005f
C60 plus.n13 a_n1724_n1488# 0.010888f
C61 plus.n14 a_n1724_n1488# 0.040005f
C62 plus.t11 a_n1724_n1488# 0.074998f
C63 plus.n15 a_n1724_n1488# 0.047888f
C64 plus.n16 a_n1724_n1488# 0.199853f
C65 plus.n17 a_n1724_n1488# 0.026435f
C66 plus.t6 a_n1724_n1488# 0.074998f
C67 plus.t12 a_n1724_n1488# 0.068897f
C68 plus.t0 a_n1724_n1488# 0.068897f
C69 plus.t4 a_n1724_n1488# 0.068897f
C70 plus.n18 a_n1724_n1488# 0.048774f
C71 plus.n19 a_n1724_n1488# 0.062281f
C72 plus.t9 a_n1724_n1488# 0.068897f
C73 plus.t10 a_n1724_n1488# 0.068897f
C74 plus.t2 a_n1724_n1488# 0.074998f
C75 plus.n20 a_n1724_n1488# 0.04793f
C76 plus.n21 a_n1724_n1488# 0.040005f
C77 plus.n22 a_n1724_n1488# 0.010888f
C78 plus.n23 a_n1724_n1488# 0.040005f
C79 plus.n24 a_n1724_n1488# 0.010888f
C80 plus.n25 a_n1724_n1488# 0.026435f
C81 plus.n26 a_n1724_n1488# 0.026435f
C82 plus.n27 a_n1724_n1488# 0.026435f
C83 plus.n28 a_n1724_n1488# 0.010888f
C84 plus.n29 a_n1724_n1488# 0.040005f
C85 plus.n30 a_n1724_n1488# 0.010888f
C86 plus.n31 a_n1724_n1488# 0.040005f
C87 plus.n32 a_n1724_n1488# 0.047888f
C88 plus.n33 a_n1724_n1488# 0.606893f
C89 source.t3 a_n1724_n1488# 0.571403f
C90 source.n0 a_n1724_n1488# 0.779585f
C91 source.t2 a_n1724_n1488# 0.068812f
C92 source.t9 a_n1724_n1488# 0.068812f
C93 source.n1 a_n1724_n1488# 0.436308f
C94 source.n2 a_n1724_n1488# 0.354447f
C95 source.t4 a_n1724_n1488# 0.068812f
C96 source.t0 a_n1724_n1488# 0.068812f
C97 source.n3 a_n1724_n1488# 0.436308f
C98 source.n4 a_n1724_n1488# 0.354447f
C99 source.t1 a_n1724_n1488# 0.068812f
C100 source.t13 a_n1724_n1488# 0.068812f
C101 source.n5 a_n1724_n1488# 0.436308f
C102 source.n6 a_n1724_n1488# 0.372991f
C103 source.t18 a_n1724_n1488# 0.571403f
C104 source.n7 a_n1724_n1488# 0.425565f
C105 source.t24 a_n1724_n1488# 0.068812f
C106 source.t15 a_n1724_n1488# 0.068812f
C107 source.n8 a_n1724_n1488# 0.436308f
C108 source.n9 a_n1724_n1488# 0.354447f
C109 source.t16 a_n1724_n1488# 0.068812f
C110 source.t19 a_n1724_n1488# 0.068812f
C111 source.n10 a_n1724_n1488# 0.436308f
C112 source.n11 a_n1724_n1488# 0.354447f
C113 source.t22 a_n1724_n1488# 0.068812f
C114 source.t26 a_n1724_n1488# 0.068812f
C115 source.n12 a_n1724_n1488# 0.436308f
C116 source.n13 a_n1724_n1488# 1.08036f
C117 source.t7 a_n1724_n1488# 0.068812f
C118 source.t12 a_n1724_n1488# 0.068812f
C119 source.n14 a_n1724_n1488# 0.436304f
C120 source.n15 a_n1724_n1488# 1.08037f
C121 source.t11 a_n1724_n1488# 0.068812f
C122 source.t5 a_n1724_n1488# 0.068812f
C123 source.n16 a_n1724_n1488# 0.436304f
C124 source.n17 a_n1724_n1488# 0.35445f
C125 source.t6 a_n1724_n1488# 0.068812f
C126 source.t8 a_n1724_n1488# 0.068812f
C127 source.n18 a_n1724_n1488# 0.436304f
C128 source.n19 a_n1724_n1488# 0.35445f
C129 source.t10 a_n1724_n1488# 0.5714f
C130 source.n20 a_n1724_n1488# 0.425568f
C131 source.t21 a_n1724_n1488# 0.068812f
C132 source.t27 a_n1724_n1488# 0.068812f
C133 source.n21 a_n1724_n1488# 0.436304f
C134 source.n22 a_n1724_n1488# 0.372994f
C135 source.t14 a_n1724_n1488# 0.068812f
C136 source.t20 a_n1724_n1488# 0.068812f
C137 source.n23 a_n1724_n1488# 0.436304f
C138 source.n24 a_n1724_n1488# 0.35445f
C139 source.t23 a_n1724_n1488# 0.068812f
C140 source.t25 a_n1724_n1488# 0.068812f
C141 source.n25 a_n1724_n1488# 0.436304f
C142 source.n26 a_n1724_n1488# 0.35445f
C143 source.t17 a_n1724_n1488# 0.5714f
C144 source.n27 a_n1724_n1488# 0.564023f
C145 source.n28 a_n1724_n1488# 0.841327f
C146 drain_right.t4 a_n1724_n1488# 0.552662f
C147 drain_right.t7 a_n1724_n1488# 0.059508f
C148 drain_right.t6 a_n1724_n1488# 0.059508f
C149 drain_right.n0 a_n1724_n1488# 0.429168f
C150 drain_right.n1 a_n1724_n1488# 0.56876f
C151 drain_right.t8 a_n1724_n1488# 0.059508f
C152 drain_right.t13 a_n1724_n1488# 0.059508f
C153 drain_right.n2 a_n1724_n1488# 0.431189f
C154 drain_right.t9 a_n1724_n1488# 0.059508f
C155 drain_right.t3 a_n1724_n1488# 0.059508f
C156 drain_right.n3 a_n1724_n1488# 0.429168f
C157 drain_right.n4 a_n1724_n1488# 0.555484f
C158 drain_right.n5 a_n1724_n1488# 0.675822f
C159 drain_right.t10 a_n1724_n1488# 0.059508f
C160 drain_right.t12 a_n1724_n1488# 0.059508f
C161 drain_right.n6 a_n1724_n1488# 0.431191f
C162 drain_right.t11 a_n1724_n1488# 0.059508f
C163 drain_right.t2 a_n1724_n1488# 0.059508f
C164 drain_right.n7 a_n1724_n1488# 0.42917f
C165 drain_right.n8 a_n1724_n1488# 0.585667f
C166 drain_right.t1 a_n1724_n1488# 0.059508f
C167 drain_right.t5 a_n1724_n1488# 0.059508f
C168 drain_right.n9 a_n1724_n1488# 0.42917f
C169 drain_right.n10 a_n1724_n1488# 0.288789f
C170 drain_right.t0 a_n1724_n1488# 0.550817f
C171 drain_right.n11 a_n1724_n1488# 0.50503f
C172 minus.n0 a_n1724_n1488# 0.026048f
C173 minus.t5 a_n1724_n1488# 0.073901f
C174 minus.t1 a_n1724_n1488# 0.067889f
C175 minus.t11 a_n1724_n1488# 0.067889f
C176 minus.t8 a_n1724_n1488# 0.067889f
C177 minus.n1 a_n1724_n1488# 0.04806f
C178 minus.n2 a_n1724_n1488# 0.061369f
C179 minus.t3 a_n1724_n1488# 0.067889f
C180 minus.t12 a_n1724_n1488# 0.067889f
C181 minus.t9 a_n1724_n1488# 0.073901f
C182 minus.n3 a_n1724_n1488# 0.047229f
C183 minus.n4 a_n1724_n1488# 0.039419f
C184 minus.n5 a_n1724_n1488# 0.010729f
C185 minus.n6 a_n1724_n1488# 0.039419f
C186 minus.n7 a_n1724_n1488# 0.010729f
C187 minus.n8 a_n1724_n1488# 0.026048f
C188 minus.n9 a_n1724_n1488# 0.026048f
C189 minus.n10 a_n1724_n1488# 0.026048f
C190 minus.n11 a_n1724_n1488# 0.010729f
C191 minus.n12 a_n1724_n1488# 0.039419f
C192 minus.n13 a_n1724_n1488# 0.010729f
C193 minus.n14 a_n1724_n1488# 0.039419f
C194 minus.n15 a_n1724_n1488# 0.047187f
C195 minus.n16 a_n1724_n1488# 0.635118f
C196 minus.n17 a_n1724_n1488# 0.026048f
C197 minus.t2 a_n1724_n1488# 0.067889f
C198 minus.t4 a_n1724_n1488# 0.067889f
C199 minus.t7 a_n1724_n1488# 0.067889f
C200 minus.n18 a_n1724_n1488# 0.04806f
C201 minus.n19 a_n1724_n1488# 0.061369f
C202 minus.t13 a_n1724_n1488# 0.067889f
C203 minus.t0 a_n1724_n1488# 0.067889f
C204 minus.t6 a_n1724_n1488# 0.073901f
C205 minus.n20 a_n1724_n1488# 0.047229f
C206 minus.n21 a_n1724_n1488# 0.039419f
C207 minus.n22 a_n1724_n1488# 0.010729f
C208 minus.n23 a_n1724_n1488# 0.039419f
C209 minus.n24 a_n1724_n1488# 0.010729f
C210 minus.n25 a_n1724_n1488# 0.026048f
C211 minus.n26 a_n1724_n1488# 0.026048f
C212 minus.n27 a_n1724_n1488# 0.026048f
C213 minus.n28 a_n1724_n1488# 0.010729f
C214 minus.n29 a_n1724_n1488# 0.039419f
C215 minus.n30 a_n1724_n1488# 0.010729f
C216 minus.n31 a_n1724_n1488# 0.039419f
C217 minus.t10 a_n1724_n1488# 0.073901f
C218 minus.n32 a_n1724_n1488# 0.047187f
C219 minus.n33 a_n1724_n1488# 0.172531f
C220 minus.n34 a_n1724_n1488# 0.783492f
.ends

