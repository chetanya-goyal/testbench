* NGSPICE file created from diffpair309.ext - technology: sky130A

.subckt diffpair309 minus drain_right drain_left source plus
X0 a_n3394_n2088# a_n3394_n2088# a_n3394_n2088# a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.7
X1 a_n3394_n2088# a_n3394_n2088# a_n3394_n2088# a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X2 drain_left.t23 plus.t0 source.t39 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X3 source.t41 plus.t1 drain_left.t22 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X4 source.t26 plus.t2 drain_left.t21 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X5 source.t24 plus.t3 drain_left.t20 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X6 source.t12 minus.t0 drain_right.t23 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X7 drain_left.t19 plus.t4 source.t42 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X8 drain_left.t18 plus.t5 source.t27 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X9 source.t30 plus.t6 drain_left.t17 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X10 source.t28 plus.t7 drain_left.t16 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X11 drain_right.t22 minus.t1 source.t15 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X12 source.t10 minus.t2 drain_right.t21 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X13 drain_right.t20 minus.t3 source.t11 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X14 drain_left.t15 plus.t8 source.t43 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X15 source.t44 plus.t9 drain_left.t14 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X16 drain_left.t13 plus.t10 source.t31 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X17 drain_right.t19 minus.t4 source.t22 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X18 source.t33 plus.t11 drain_left.t12 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X19 drain_left.t11 plus.t12 source.t36 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X20 a_n3394_n2088# a_n3394_n2088# a_n3394_n2088# a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X21 drain_right.t18 minus.t5 source.t13 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X22 drain_right.t17 minus.t6 source.t2 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X23 drain_right.t16 minus.t7 source.t14 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X24 source.t16 minus.t8 drain_right.t15 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X25 source.t45 plus.t13 drain_left.t10 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X26 drain_left.t9 plus.t14 source.t32 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X27 drain_left.t8 plus.t15 source.t34 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X28 drain_right.t14 minus.t9 source.t0 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X29 source.t19 minus.t10 drain_right.t13 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X30 source.t29 plus.t16 drain_left.t7 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X31 drain_left.t6 plus.t17 source.t25 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X32 drain_right.t12 minus.t11 source.t1 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X33 source.t37 plus.t18 drain_left.t5 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X34 drain_left.t4 plus.t19 source.t46 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X35 drain_right.t11 minus.t12 source.t9 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X36 a_n3394_n2088# a_n3394_n2088# a_n3394_n2088# a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X37 source.t5 minus.t13 drain_right.t10 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X38 drain_left.t3 plus.t20 source.t38 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X39 source.t8 minus.t14 drain_right.t9 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X40 source.t6 minus.t15 drain_right.t8 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X41 drain_right.t7 minus.t16 source.t21 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X42 source.t40 plus.t21 drain_left.t2 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X43 drain_left.t1 plus.t22 source.t35 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X44 source.t18 minus.t17 drain_right.t6 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X45 source.t7 minus.t18 drain_right.t5 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X46 drain_right.t4 minus.t19 source.t17 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X47 source.t4 minus.t20 drain_right.t3 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X48 drain_right.t2 minus.t21 source.t20 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X49 source.t3 minus.t22 drain_right.t1 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X50 source.t47 minus.t23 drain_right.t0 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X51 source.t23 plus.t23 drain_left.t0 a_n3394_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
R0 plus.n11 plus.t7 289.048
R1 plus.n53 plus.t15 289.048
R2 plus.n40 plus.t0 262.69
R3 plus.n38 plus.t18 262.69
R4 plus.n2 plus.t5 262.69
R5 plus.n32 plus.t23 262.69
R6 plus.n4 plus.t14 262.69
R7 plus.n26 plus.t1 262.69
R8 plus.n6 plus.t19 262.69
R9 plus.n20 plus.t6 262.69
R10 plus.n8 plus.t17 262.69
R11 plus.n14 plus.t3 262.69
R12 plus.n10 plus.t20 262.69
R13 plus.n82 plus.t11 262.69
R14 plus.n80 plus.t10 262.69
R15 plus.n44 plus.t9 262.69
R16 plus.n74 plus.t8 262.69
R17 plus.n46 plus.t13 262.69
R18 plus.n68 plus.t22 262.69
R19 plus.n48 plus.t21 262.69
R20 plus.n62 plus.t4 262.69
R21 plus.n50 plus.t2 262.69
R22 plus.n56 plus.t12 262.69
R23 plus.n52 plus.t16 262.69
R24 plus.n13 plus.n12 161.3
R25 plus.n14 plus.n9 161.3
R26 plus.n16 plus.n15 161.3
R27 plus.n17 plus.n8 161.3
R28 plus.n19 plus.n18 161.3
R29 plus.n20 plus.n7 161.3
R30 plus.n22 plus.n21 161.3
R31 plus.n23 plus.n6 161.3
R32 plus.n25 plus.n24 161.3
R33 plus.n26 plus.n5 161.3
R34 plus.n28 plus.n27 161.3
R35 plus.n29 plus.n4 161.3
R36 plus.n31 plus.n30 161.3
R37 plus.n32 plus.n3 161.3
R38 plus.n34 plus.n33 161.3
R39 plus.n35 plus.n2 161.3
R40 plus.n37 plus.n36 161.3
R41 plus.n38 plus.n1 161.3
R42 plus.n39 plus.n0 161.3
R43 plus.n41 plus.n40 161.3
R44 plus.n55 plus.n54 161.3
R45 plus.n56 plus.n51 161.3
R46 plus.n58 plus.n57 161.3
R47 plus.n59 plus.n50 161.3
R48 plus.n61 plus.n60 161.3
R49 plus.n62 plus.n49 161.3
R50 plus.n64 plus.n63 161.3
R51 plus.n65 plus.n48 161.3
R52 plus.n67 plus.n66 161.3
R53 plus.n68 plus.n47 161.3
R54 plus.n70 plus.n69 161.3
R55 plus.n71 plus.n46 161.3
R56 plus.n73 plus.n72 161.3
R57 plus.n74 plus.n45 161.3
R58 plus.n76 plus.n75 161.3
R59 plus.n77 plus.n44 161.3
R60 plus.n79 plus.n78 161.3
R61 plus.n80 plus.n43 161.3
R62 plus.n81 plus.n42 161.3
R63 plus.n83 plus.n82 161.3
R64 plus.n40 plus.n39 46.0096
R65 plus.n82 plus.n81 46.0096
R66 plus.n12 plus.n11 45.0871
R67 plus.n54 plus.n53 45.0871
R68 plus.n38 plus.n37 41.6278
R69 plus.n13 plus.n10 41.6278
R70 plus.n80 plus.n79 41.6278
R71 plus.n55 plus.n52 41.6278
R72 plus.n33 plus.n2 37.246
R73 plus.n15 plus.n14 37.246
R74 plus.n75 plus.n44 37.246
R75 plus.n57 plus.n56 37.246
R76 plus plus.n83 33.7642
R77 plus.n32 plus.n31 32.8641
R78 plus.n19 plus.n8 32.8641
R79 plus.n74 plus.n73 32.8641
R80 plus.n61 plus.n50 32.8641
R81 plus.n27 plus.n4 28.4823
R82 plus.n21 plus.n20 28.4823
R83 plus.n69 plus.n46 28.4823
R84 plus.n63 plus.n62 28.4823
R85 plus.n25 plus.n6 24.1005
R86 plus.n26 plus.n25 24.1005
R87 plus.n68 plus.n67 24.1005
R88 plus.n67 plus.n48 24.1005
R89 plus.n27 plus.n26 19.7187
R90 plus.n21 plus.n6 19.7187
R91 plus.n69 plus.n68 19.7187
R92 plus.n63 plus.n48 19.7187
R93 plus.n31 plus.n4 15.3369
R94 plus.n20 plus.n19 15.3369
R95 plus.n73 plus.n46 15.3369
R96 plus.n62 plus.n61 15.3369
R97 plus.n11 plus.n10 14.1472
R98 plus.n53 plus.n52 14.1472
R99 plus.n33 plus.n32 10.955
R100 plus.n15 plus.n8 10.955
R101 plus.n75 plus.n74 10.955
R102 plus.n57 plus.n50 10.955
R103 plus plus.n41 10.0497
R104 plus.n37 plus.n2 6.57323
R105 plus.n14 plus.n13 6.57323
R106 plus.n79 plus.n44 6.57323
R107 plus.n56 plus.n55 6.57323
R108 plus.n39 plus.n38 2.19141
R109 plus.n81 plus.n80 2.19141
R110 plus.n12 plus.n9 0.189894
R111 plus.n16 plus.n9 0.189894
R112 plus.n17 plus.n16 0.189894
R113 plus.n18 plus.n17 0.189894
R114 plus.n18 plus.n7 0.189894
R115 plus.n22 plus.n7 0.189894
R116 plus.n23 plus.n22 0.189894
R117 plus.n24 plus.n23 0.189894
R118 plus.n24 plus.n5 0.189894
R119 plus.n28 plus.n5 0.189894
R120 plus.n29 plus.n28 0.189894
R121 plus.n30 plus.n29 0.189894
R122 plus.n30 plus.n3 0.189894
R123 plus.n34 plus.n3 0.189894
R124 plus.n35 plus.n34 0.189894
R125 plus.n36 plus.n35 0.189894
R126 plus.n36 plus.n1 0.189894
R127 plus.n1 plus.n0 0.189894
R128 plus.n41 plus.n0 0.189894
R129 plus.n83 plus.n42 0.189894
R130 plus.n43 plus.n42 0.189894
R131 plus.n78 plus.n43 0.189894
R132 plus.n78 plus.n77 0.189894
R133 plus.n77 plus.n76 0.189894
R134 plus.n76 plus.n45 0.189894
R135 plus.n72 plus.n45 0.189894
R136 plus.n72 plus.n71 0.189894
R137 plus.n71 plus.n70 0.189894
R138 plus.n70 plus.n47 0.189894
R139 plus.n66 plus.n47 0.189894
R140 plus.n66 plus.n65 0.189894
R141 plus.n65 plus.n64 0.189894
R142 plus.n64 plus.n49 0.189894
R143 plus.n60 plus.n49 0.189894
R144 plus.n60 plus.n59 0.189894
R145 plus.n59 plus.n58 0.189894
R146 plus.n58 plus.n51 0.189894
R147 plus.n54 plus.n51 0.189894
R148 source.n290 source.n264 289.615
R149 source.n248 source.n222 289.615
R150 source.n216 source.n190 289.615
R151 source.n174 source.n148 289.615
R152 source.n26 source.n0 289.615
R153 source.n68 source.n42 289.615
R154 source.n100 source.n74 289.615
R155 source.n142 source.n116 289.615
R156 source.n275 source.n274 185
R157 source.n272 source.n271 185
R158 source.n281 source.n280 185
R159 source.n283 source.n282 185
R160 source.n268 source.n267 185
R161 source.n289 source.n288 185
R162 source.n291 source.n290 185
R163 source.n233 source.n232 185
R164 source.n230 source.n229 185
R165 source.n239 source.n238 185
R166 source.n241 source.n240 185
R167 source.n226 source.n225 185
R168 source.n247 source.n246 185
R169 source.n249 source.n248 185
R170 source.n201 source.n200 185
R171 source.n198 source.n197 185
R172 source.n207 source.n206 185
R173 source.n209 source.n208 185
R174 source.n194 source.n193 185
R175 source.n215 source.n214 185
R176 source.n217 source.n216 185
R177 source.n159 source.n158 185
R178 source.n156 source.n155 185
R179 source.n165 source.n164 185
R180 source.n167 source.n166 185
R181 source.n152 source.n151 185
R182 source.n173 source.n172 185
R183 source.n175 source.n174 185
R184 source.n27 source.n26 185
R185 source.n25 source.n24 185
R186 source.n4 source.n3 185
R187 source.n19 source.n18 185
R188 source.n17 source.n16 185
R189 source.n8 source.n7 185
R190 source.n11 source.n10 185
R191 source.n69 source.n68 185
R192 source.n67 source.n66 185
R193 source.n46 source.n45 185
R194 source.n61 source.n60 185
R195 source.n59 source.n58 185
R196 source.n50 source.n49 185
R197 source.n53 source.n52 185
R198 source.n101 source.n100 185
R199 source.n99 source.n98 185
R200 source.n78 source.n77 185
R201 source.n93 source.n92 185
R202 source.n91 source.n90 185
R203 source.n82 source.n81 185
R204 source.n85 source.n84 185
R205 source.n143 source.n142 185
R206 source.n141 source.n140 185
R207 source.n120 source.n119 185
R208 source.n135 source.n134 185
R209 source.n133 source.n132 185
R210 source.n124 source.n123 185
R211 source.n127 source.n126 185
R212 source.t21 source.n273 147.661
R213 source.t18 source.n231 147.661
R214 source.t34 source.n199 147.661
R215 source.t33 source.n157 147.661
R216 source.t39 source.n9 147.661
R217 source.t28 source.n51 147.661
R218 source.t9 source.n83 147.661
R219 source.t8 source.n125 147.661
R220 source.n274 source.n271 104.615
R221 source.n281 source.n271 104.615
R222 source.n282 source.n281 104.615
R223 source.n282 source.n267 104.615
R224 source.n289 source.n267 104.615
R225 source.n290 source.n289 104.615
R226 source.n232 source.n229 104.615
R227 source.n239 source.n229 104.615
R228 source.n240 source.n239 104.615
R229 source.n240 source.n225 104.615
R230 source.n247 source.n225 104.615
R231 source.n248 source.n247 104.615
R232 source.n200 source.n197 104.615
R233 source.n207 source.n197 104.615
R234 source.n208 source.n207 104.615
R235 source.n208 source.n193 104.615
R236 source.n215 source.n193 104.615
R237 source.n216 source.n215 104.615
R238 source.n158 source.n155 104.615
R239 source.n165 source.n155 104.615
R240 source.n166 source.n165 104.615
R241 source.n166 source.n151 104.615
R242 source.n173 source.n151 104.615
R243 source.n174 source.n173 104.615
R244 source.n26 source.n25 104.615
R245 source.n25 source.n3 104.615
R246 source.n18 source.n3 104.615
R247 source.n18 source.n17 104.615
R248 source.n17 source.n7 104.615
R249 source.n10 source.n7 104.615
R250 source.n68 source.n67 104.615
R251 source.n67 source.n45 104.615
R252 source.n60 source.n45 104.615
R253 source.n60 source.n59 104.615
R254 source.n59 source.n49 104.615
R255 source.n52 source.n49 104.615
R256 source.n100 source.n99 104.615
R257 source.n99 source.n77 104.615
R258 source.n92 source.n77 104.615
R259 source.n92 source.n91 104.615
R260 source.n91 source.n81 104.615
R261 source.n84 source.n81 104.615
R262 source.n142 source.n141 104.615
R263 source.n141 source.n119 104.615
R264 source.n134 source.n119 104.615
R265 source.n134 source.n133 104.615
R266 source.n133 source.n123 104.615
R267 source.n126 source.n123 104.615
R268 source.n274 source.t21 52.3082
R269 source.n232 source.t18 52.3082
R270 source.n200 source.t34 52.3082
R271 source.n158 source.t33 52.3082
R272 source.n10 source.t39 52.3082
R273 source.n52 source.t28 52.3082
R274 source.n84 source.t9 52.3082
R275 source.n126 source.t8 52.3082
R276 source.n33 source.n32 50.512
R277 source.n35 source.n34 50.512
R278 source.n37 source.n36 50.512
R279 source.n39 source.n38 50.512
R280 source.n41 source.n40 50.512
R281 source.n107 source.n106 50.512
R282 source.n109 source.n108 50.512
R283 source.n111 source.n110 50.512
R284 source.n113 source.n112 50.512
R285 source.n115 source.n114 50.512
R286 source.n263 source.n262 50.5119
R287 source.n261 source.n260 50.5119
R288 source.n259 source.n258 50.5119
R289 source.n257 source.n256 50.5119
R290 source.n255 source.n254 50.5119
R291 source.n189 source.n188 50.5119
R292 source.n187 source.n186 50.5119
R293 source.n185 source.n184 50.5119
R294 source.n183 source.n182 50.5119
R295 source.n181 source.n180 50.5119
R296 source.n295 source.n294 32.1853
R297 source.n253 source.n252 32.1853
R298 source.n221 source.n220 32.1853
R299 source.n179 source.n178 32.1853
R300 source.n31 source.n30 32.1853
R301 source.n73 source.n72 32.1853
R302 source.n105 source.n104 32.1853
R303 source.n147 source.n146 32.1853
R304 source.n179 source.n147 17.6302
R305 source.n275 source.n273 15.6674
R306 source.n233 source.n231 15.6674
R307 source.n201 source.n199 15.6674
R308 source.n159 source.n157 15.6674
R309 source.n11 source.n9 15.6674
R310 source.n53 source.n51 15.6674
R311 source.n85 source.n83 15.6674
R312 source.n127 source.n125 15.6674
R313 source.n276 source.n272 12.8005
R314 source.n234 source.n230 12.8005
R315 source.n202 source.n198 12.8005
R316 source.n160 source.n156 12.8005
R317 source.n12 source.n8 12.8005
R318 source.n54 source.n50 12.8005
R319 source.n86 source.n82 12.8005
R320 source.n128 source.n124 12.8005
R321 source.n280 source.n279 12.0247
R322 source.n238 source.n237 12.0247
R323 source.n206 source.n205 12.0247
R324 source.n164 source.n163 12.0247
R325 source.n16 source.n15 12.0247
R326 source.n58 source.n57 12.0247
R327 source.n90 source.n89 12.0247
R328 source.n132 source.n131 12.0247
R329 source.n296 source.n31 11.9233
R330 source.n283 source.n270 11.249
R331 source.n241 source.n228 11.249
R332 source.n209 source.n196 11.249
R333 source.n167 source.n154 11.249
R334 source.n19 source.n6 11.249
R335 source.n61 source.n48 11.249
R336 source.n93 source.n80 11.249
R337 source.n135 source.n122 11.249
R338 source.n284 source.n268 10.4732
R339 source.n242 source.n226 10.4732
R340 source.n210 source.n194 10.4732
R341 source.n168 source.n152 10.4732
R342 source.n20 source.n4 10.4732
R343 source.n62 source.n46 10.4732
R344 source.n94 source.n78 10.4732
R345 source.n136 source.n120 10.4732
R346 source.n288 source.n287 9.69747
R347 source.n246 source.n245 9.69747
R348 source.n214 source.n213 9.69747
R349 source.n172 source.n171 9.69747
R350 source.n24 source.n23 9.69747
R351 source.n66 source.n65 9.69747
R352 source.n98 source.n97 9.69747
R353 source.n140 source.n139 9.69747
R354 source.n294 source.n293 9.45567
R355 source.n252 source.n251 9.45567
R356 source.n220 source.n219 9.45567
R357 source.n178 source.n177 9.45567
R358 source.n30 source.n29 9.45567
R359 source.n72 source.n71 9.45567
R360 source.n104 source.n103 9.45567
R361 source.n146 source.n145 9.45567
R362 source.n293 source.n292 9.3005
R363 source.n266 source.n265 9.3005
R364 source.n287 source.n286 9.3005
R365 source.n285 source.n284 9.3005
R366 source.n270 source.n269 9.3005
R367 source.n279 source.n278 9.3005
R368 source.n277 source.n276 9.3005
R369 source.n251 source.n250 9.3005
R370 source.n224 source.n223 9.3005
R371 source.n245 source.n244 9.3005
R372 source.n243 source.n242 9.3005
R373 source.n228 source.n227 9.3005
R374 source.n237 source.n236 9.3005
R375 source.n235 source.n234 9.3005
R376 source.n219 source.n218 9.3005
R377 source.n192 source.n191 9.3005
R378 source.n213 source.n212 9.3005
R379 source.n211 source.n210 9.3005
R380 source.n196 source.n195 9.3005
R381 source.n205 source.n204 9.3005
R382 source.n203 source.n202 9.3005
R383 source.n177 source.n176 9.3005
R384 source.n150 source.n149 9.3005
R385 source.n171 source.n170 9.3005
R386 source.n169 source.n168 9.3005
R387 source.n154 source.n153 9.3005
R388 source.n163 source.n162 9.3005
R389 source.n161 source.n160 9.3005
R390 source.n29 source.n28 9.3005
R391 source.n2 source.n1 9.3005
R392 source.n23 source.n22 9.3005
R393 source.n21 source.n20 9.3005
R394 source.n6 source.n5 9.3005
R395 source.n15 source.n14 9.3005
R396 source.n13 source.n12 9.3005
R397 source.n71 source.n70 9.3005
R398 source.n44 source.n43 9.3005
R399 source.n65 source.n64 9.3005
R400 source.n63 source.n62 9.3005
R401 source.n48 source.n47 9.3005
R402 source.n57 source.n56 9.3005
R403 source.n55 source.n54 9.3005
R404 source.n103 source.n102 9.3005
R405 source.n76 source.n75 9.3005
R406 source.n97 source.n96 9.3005
R407 source.n95 source.n94 9.3005
R408 source.n80 source.n79 9.3005
R409 source.n89 source.n88 9.3005
R410 source.n87 source.n86 9.3005
R411 source.n145 source.n144 9.3005
R412 source.n118 source.n117 9.3005
R413 source.n139 source.n138 9.3005
R414 source.n137 source.n136 9.3005
R415 source.n122 source.n121 9.3005
R416 source.n131 source.n130 9.3005
R417 source.n129 source.n128 9.3005
R418 source.n291 source.n266 8.92171
R419 source.n249 source.n224 8.92171
R420 source.n217 source.n192 8.92171
R421 source.n175 source.n150 8.92171
R422 source.n27 source.n2 8.92171
R423 source.n69 source.n44 8.92171
R424 source.n101 source.n76 8.92171
R425 source.n143 source.n118 8.92171
R426 source.n292 source.n264 8.14595
R427 source.n250 source.n222 8.14595
R428 source.n218 source.n190 8.14595
R429 source.n176 source.n148 8.14595
R430 source.n28 source.n0 8.14595
R431 source.n70 source.n42 8.14595
R432 source.n102 source.n74 8.14595
R433 source.n144 source.n116 8.14595
R434 source.n294 source.n264 5.81868
R435 source.n252 source.n222 5.81868
R436 source.n220 source.n190 5.81868
R437 source.n178 source.n148 5.81868
R438 source.n30 source.n0 5.81868
R439 source.n72 source.n42 5.81868
R440 source.n104 source.n74 5.81868
R441 source.n146 source.n116 5.81868
R442 source.n296 source.n295 5.7074
R443 source.n292 source.n291 5.04292
R444 source.n250 source.n249 5.04292
R445 source.n218 source.n217 5.04292
R446 source.n176 source.n175 5.04292
R447 source.n28 source.n27 5.04292
R448 source.n70 source.n69 5.04292
R449 source.n102 source.n101 5.04292
R450 source.n144 source.n143 5.04292
R451 source.n277 source.n273 4.38594
R452 source.n235 source.n231 4.38594
R453 source.n203 source.n199 4.38594
R454 source.n161 source.n157 4.38594
R455 source.n13 source.n9 4.38594
R456 source.n55 source.n51 4.38594
R457 source.n87 source.n83 4.38594
R458 source.n129 source.n125 4.38594
R459 source.n288 source.n266 4.26717
R460 source.n246 source.n224 4.26717
R461 source.n214 source.n192 4.26717
R462 source.n172 source.n150 4.26717
R463 source.n24 source.n2 4.26717
R464 source.n66 source.n44 4.26717
R465 source.n98 source.n76 4.26717
R466 source.n140 source.n118 4.26717
R467 source.n287 source.n268 3.49141
R468 source.n245 source.n226 3.49141
R469 source.n213 source.n194 3.49141
R470 source.n171 source.n152 3.49141
R471 source.n23 source.n4 3.49141
R472 source.n65 source.n46 3.49141
R473 source.n97 source.n78 3.49141
R474 source.n139 source.n120 3.49141
R475 source.n262 source.t20 3.3005
R476 source.n262 source.t6 3.3005
R477 source.n260 source.t11 3.3005
R478 source.n260 source.t10 3.3005
R479 source.n258 source.t2 3.3005
R480 source.n258 source.t16 3.3005
R481 source.n256 source.t1 3.3005
R482 source.n256 source.t5 3.3005
R483 source.n254 source.t17 3.3005
R484 source.n254 source.t19 3.3005
R485 source.n188 source.t36 3.3005
R486 source.n188 source.t29 3.3005
R487 source.n186 source.t42 3.3005
R488 source.n186 source.t26 3.3005
R489 source.n184 source.t35 3.3005
R490 source.n184 source.t40 3.3005
R491 source.n182 source.t43 3.3005
R492 source.n182 source.t45 3.3005
R493 source.n180 source.t31 3.3005
R494 source.n180 source.t44 3.3005
R495 source.n32 source.t27 3.3005
R496 source.n32 source.t37 3.3005
R497 source.n34 source.t32 3.3005
R498 source.n34 source.t23 3.3005
R499 source.n36 source.t46 3.3005
R500 source.n36 source.t41 3.3005
R501 source.n38 source.t25 3.3005
R502 source.n38 source.t30 3.3005
R503 source.n40 source.t38 3.3005
R504 source.n40 source.t24 3.3005
R505 source.n106 source.t0 3.3005
R506 source.n106 source.t12 3.3005
R507 source.n108 source.t14 3.3005
R508 source.n108 source.t3 3.3005
R509 source.n110 source.t13 3.3005
R510 source.n110 source.t47 3.3005
R511 source.n112 source.t22 3.3005
R512 source.n112 source.t4 3.3005
R513 source.n114 source.t15 3.3005
R514 source.n114 source.t7 3.3005
R515 source.n284 source.n283 2.71565
R516 source.n242 source.n241 2.71565
R517 source.n210 source.n209 2.71565
R518 source.n168 source.n167 2.71565
R519 source.n20 source.n19 2.71565
R520 source.n62 source.n61 2.71565
R521 source.n94 source.n93 2.71565
R522 source.n136 source.n135 2.71565
R523 source.n280 source.n270 1.93989
R524 source.n238 source.n228 1.93989
R525 source.n206 source.n196 1.93989
R526 source.n164 source.n154 1.93989
R527 source.n16 source.n6 1.93989
R528 source.n58 source.n48 1.93989
R529 source.n90 source.n80 1.93989
R530 source.n132 source.n122 1.93989
R531 source.n279 source.n272 1.16414
R532 source.n237 source.n230 1.16414
R533 source.n205 source.n198 1.16414
R534 source.n163 source.n156 1.16414
R535 source.n15 source.n8 1.16414
R536 source.n57 source.n50 1.16414
R537 source.n89 source.n82 1.16414
R538 source.n131 source.n124 1.16414
R539 source.n147 source.n115 0.888431
R540 source.n115 source.n113 0.888431
R541 source.n113 source.n111 0.888431
R542 source.n111 source.n109 0.888431
R543 source.n109 source.n107 0.888431
R544 source.n107 source.n105 0.888431
R545 source.n73 source.n41 0.888431
R546 source.n41 source.n39 0.888431
R547 source.n39 source.n37 0.888431
R548 source.n37 source.n35 0.888431
R549 source.n35 source.n33 0.888431
R550 source.n33 source.n31 0.888431
R551 source.n181 source.n179 0.888431
R552 source.n183 source.n181 0.888431
R553 source.n185 source.n183 0.888431
R554 source.n187 source.n185 0.888431
R555 source.n189 source.n187 0.888431
R556 source.n221 source.n189 0.888431
R557 source.n255 source.n253 0.888431
R558 source.n257 source.n255 0.888431
R559 source.n259 source.n257 0.888431
R560 source.n261 source.n259 0.888431
R561 source.n263 source.n261 0.888431
R562 source.n295 source.n263 0.888431
R563 source.n105 source.n73 0.470328
R564 source.n253 source.n221 0.470328
R565 source.n276 source.n275 0.388379
R566 source.n234 source.n233 0.388379
R567 source.n202 source.n201 0.388379
R568 source.n160 source.n159 0.388379
R569 source.n12 source.n11 0.388379
R570 source.n54 source.n53 0.388379
R571 source.n86 source.n85 0.388379
R572 source.n128 source.n127 0.388379
R573 source source.n296 0.188
R574 source.n278 source.n277 0.155672
R575 source.n278 source.n269 0.155672
R576 source.n285 source.n269 0.155672
R577 source.n286 source.n285 0.155672
R578 source.n286 source.n265 0.155672
R579 source.n293 source.n265 0.155672
R580 source.n236 source.n235 0.155672
R581 source.n236 source.n227 0.155672
R582 source.n243 source.n227 0.155672
R583 source.n244 source.n243 0.155672
R584 source.n244 source.n223 0.155672
R585 source.n251 source.n223 0.155672
R586 source.n204 source.n203 0.155672
R587 source.n204 source.n195 0.155672
R588 source.n211 source.n195 0.155672
R589 source.n212 source.n211 0.155672
R590 source.n212 source.n191 0.155672
R591 source.n219 source.n191 0.155672
R592 source.n162 source.n161 0.155672
R593 source.n162 source.n153 0.155672
R594 source.n169 source.n153 0.155672
R595 source.n170 source.n169 0.155672
R596 source.n170 source.n149 0.155672
R597 source.n177 source.n149 0.155672
R598 source.n29 source.n1 0.155672
R599 source.n22 source.n1 0.155672
R600 source.n22 source.n21 0.155672
R601 source.n21 source.n5 0.155672
R602 source.n14 source.n5 0.155672
R603 source.n14 source.n13 0.155672
R604 source.n71 source.n43 0.155672
R605 source.n64 source.n43 0.155672
R606 source.n64 source.n63 0.155672
R607 source.n63 source.n47 0.155672
R608 source.n56 source.n47 0.155672
R609 source.n56 source.n55 0.155672
R610 source.n103 source.n75 0.155672
R611 source.n96 source.n75 0.155672
R612 source.n96 source.n95 0.155672
R613 source.n95 source.n79 0.155672
R614 source.n88 source.n79 0.155672
R615 source.n88 source.n87 0.155672
R616 source.n145 source.n117 0.155672
R617 source.n138 source.n117 0.155672
R618 source.n138 source.n137 0.155672
R619 source.n137 source.n121 0.155672
R620 source.n130 source.n121 0.155672
R621 source.n130 source.n129 0.155672
R622 drain_left.n13 drain_left.n11 68.0787
R623 drain_left.n7 drain_left.n5 68.0786
R624 drain_left.n2 drain_left.n0 68.0786
R625 drain_left.n19 drain_left.n18 67.1908
R626 drain_left.n17 drain_left.n16 67.1908
R627 drain_left.n15 drain_left.n14 67.1908
R628 drain_left.n13 drain_left.n12 67.1908
R629 drain_left.n21 drain_left.n20 67.1907
R630 drain_left.n7 drain_left.n6 67.1907
R631 drain_left.n9 drain_left.n8 67.1907
R632 drain_left.n4 drain_left.n3 67.1907
R633 drain_left.n2 drain_left.n1 67.1907
R634 drain_left drain_left.n10 31.257
R635 drain_left drain_left.n21 6.54115
R636 drain_left.n5 drain_left.t7 3.3005
R637 drain_left.n5 drain_left.t8 3.3005
R638 drain_left.n6 drain_left.t21 3.3005
R639 drain_left.n6 drain_left.t11 3.3005
R640 drain_left.n8 drain_left.t2 3.3005
R641 drain_left.n8 drain_left.t19 3.3005
R642 drain_left.n3 drain_left.t10 3.3005
R643 drain_left.n3 drain_left.t1 3.3005
R644 drain_left.n1 drain_left.t14 3.3005
R645 drain_left.n1 drain_left.t15 3.3005
R646 drain_left.n0 drain_left.t12 3.3005
R647 drain_left.n0 drain_left.t13 3.3005
R648 drain_left.n20 drain_left.t5 3.3005
R649 drain_left.n20 drain_left.t23 3.3005
R650 drain_left.n18 drain_left.t0 3.3005
R651 drain_left.n18 drain_left.t18 3.3005
R652 drain_left.n16 drain_left.t22 3.3005
R653 drain_left.n16 drain_left.t9 3.3005
R654 drain_left.n14 drain_left.t17 3.3005
R655 drain_left.n14 drain_left.t4 3.3005
R656 drain_left.n12 drain_left.t20 3.3005
R657 drain_left.n12 drain_left.t6 3.3005
R658 drain_left.n11 drain_left.t16 3.3005
R659 drain_left.n11 drain_left.t3 3.3005
R660 drain_left.n9 drain_left.n7 0.888431
R661 drain_left.n4 drain_left.n2 0.888431
R662 drain_left.n15 drain_left.n13 0.888431
R663 drain_left.n17 drain_left.n15 0.888431
R664 drain_left.n19 drain_left.n17 0.888431
R665 drain_left.n21 drain_left.n19 0.888431
R666 drain_left.n10 drain_left.n9 0.389119
R667 drain_left.n10 drain_left.n4 0.389119
R668 minus.n11 minus.t12 289.048
R669 minus.n53 minus.t17 289.048
R670 minus.n10 minus.t0 262.69
R671 minus.n14 minus.t9 262.69
R672 minus.n16 minus.t22 262.69
R673 minus.n20 minus.t7 262.69
R674 minus.n22 minus.t23 262.69
R675 minus.n26 minus.t5 262.69
R676 minus.n28 minus.t20 262.69
R677 minus.n32 minus.t4 262.69
R678 minus.n34 minus.t18 262.69
R679 minus.n38 minus.t1 262.69
R680 minus.n40 minus.t14 262.69
R681 minus.n52 minus.t19 262.69
R682 minus.n56 minus.t10 262.69
R683 minus.n58 minus.t11 262.69
R684 minus.n62 minus.t13 262.69
R685 minus.n64 minus.t6 262.69
R686 minus.n68 minus.t8 262.69
R687 minus.n70 minus.t3 262.69
R688 minus.n74 minus.t2 262.69
R689 minus.n76 minus.t21 262.69
R690 minus.n80 minus.t15 262.69
R691 minus.n82 minus.t16 262.69
R692 minus.n41 minus.n40 161.3
R693 minus.n39 minus.n0 161.3
R694 minus.n38 minus.n37 161.3
R695 minus.n36 minus.n1 161.3
R696 minus.n35 minus.n34 161.3
R697 minus.n33 minus.n2 161.3
R698 minus.n32 minus.n31 161.3
R699 minus.n30 minus.n3 161.3
R700 minus.n29 minus.n28 161.3
R701 minus.n27 minus.n4 161.3
R702 minus.n26 minus.n25 161.3
R703 minus.n24 minus.n5 161.3
R704 minus.n23 minus.n22 161.3
R705 minus.n21 minus.n6 161.3
R706 minus.n20 minus.n19 161.3
R707 minus.n18 minus.n7 161.3
R708 minus.n17 minus.n16 161.3
R709 minus.n15 minus.n8 161.3
R710 minus.n14 minus.n13 161.3
R711 minus.n12 minus.n9 161.3
R712 minus.n83 minus.n82 161.3
R713 minus.n81 minus.n42 161.3
R714 minus.n80 minus.n79 161.3
R715 minus.n78 minus.n43 161.3
R716 minus.n77 minus.n76 161.3
R717 minus.n75 minus.n44 161.3
R718 minus.n74 minus.n73 161.3
R719 minus.n72 minus.n45 161.3
R720 minus.n71 minus.n70 161.3
R721 minus.n69 minus.n46 161.3
R722 minus.n68 minus.n67 161.3
R723 minus.n66 minus.n47 161.3
R724 minus.n65 minus.n64 161.3
R725 minus.n63 minus.n48 161.3
R726 minus.n62 minus.n61 161.3
R727 minus.n60 minus.n49 161.3
R728 minus.n59 minus.n58 161.3
R729 minus.n57 minus.n50 161.3
R730 minus.n56 minus.n55 161.3
R731 minus.n54 minus.n51 161.3
R732 minus.n40 minus.n39 46.0096
R733 minus.n82 minus.n81 46.0096
R734 minus.n12 minus.n11 45.0871
R735 minus.n54 minus.n53 45.0871
R736 minus.n10 minus.n9 41.6278
R737 minus.n38 minus.n1 41.6278
R738 minus.n52 minus.n51 41.6278
R739 minus.n80 minus.n43 41.6278
R740 minus.n84 minus.n41 37.6104
R741 minus.n15 minus.n14 37.246
R742 minus.n34 minus.n33 37.246
R743 minus.n57 minus.n56 37.246
R744 minus.n76 minus.n75 37.246
R745 minus.n16 minus.n7 32.8641
R746 minus.n32 minus.n3 32.8641
R747 minus.n58 minus.n49 32.8641
R748 minus.n74 minus.n45 32.8641
R749 minus.n21 minus.n20 28.4823
R750 minus.n28 minus.n27 28.4823
R751 minus.n63 minus.n62 28.4823
R752 minus.n70 minus.n69 28.4823
R753 minus.n26 minus.n5 24.1005
R754 minus.n22 minus.n5 24.1005
R755 minus.n64 minus.n47 24.1005
R756 minus.n68 minus.n47 24.1005
R757 minus.n22 minus.n21 19.7187
R758 minus.n27 minus.n26 19.7187
R759 minus.n64 minus.n63 19.7187
R760 minus.n69 minus.n68 19.7187
R761 minus.n20 minus.n7 15.3369
R762 minus.n28 minus.n3 15.3369
R763 minus.n62 minus.n49 15.3369
R764 minus.n70 minus.n45 15.3369
R765 minus.n11 minus.n10 14.1472
R766 minus.n53 minus.n52 14.1472
R767 minus.n16 minus.n15 10.955
R768 minus.n33 minus.n32 10.955
R769 minus.n58 minus.n57 10.955
R770 minus.n75 minus.n74 10.955
R771 minus.n84 minus.n83 6.67853
R772 minus.n14 minus.n9 6.57323
R773 minus.n34 minus.n1 6.57323
R774 minus.n56 minus.n51 6.57323
R775 minus.n76 minus.n43 6.57323
R776 minus.n39 minus.n38 2.19141
R777 minus.n81 minus.n80 2.19141
R778 minus.n41 minus.n0 0.189894
R779 minus.n37 minus.n0 0.189894
R780 minus.n37 minus.n36 0.189894
R781 minus.n36 minus.n35 0.189894
R782 minus.n35 minus.n2 0.189894
R783 minus.n31 minus.n2 0.189894
R784 minus.n31 minus.n30 0.189894
R785 minus.n30 minus.n29 0.189894
R786 minus.n29 minus.n4 0.189894
R787 minus.n25 minus.n4 0.189894
R788 minus.n25 minus.n24 0.189894
R789 minus.n24 minus.n23 0.189894
R790 minus.n23 minus.n6 0.189894
R791 minus.n19 minus.n6 0.189894
R792 minus.n19 minus.n18 0.189894
R793 minus.n18 minus.n17 0.189894
R794 minus.n17 minus.n8 0.189894
R795 minus.n13 minus.n8 0.189894
R796 minus.n13 minus.n12 0.189894
R797 minus.n55 minus.n54 0.189894
R798 minus.n55 minus.n50 0.189894
R799 minus.n59 minus.n50 0.189894
R800 minus.n60 minus.n59 0.189894
R801 minus.n61 minus.n60 0.189894
R802 minus.n61 minus.n48 0.189894
R803 minus.n65 minus.n48 0.189894
R804 minus.n66 minus.n65 0.189894
R805 minus.n67 minus.n66 0.189894
R806 minus.n67 minus.n46 0.189894
R807 minus.n71 minus.n46 0.189894
R808 minus.n72 minus.n71 0.189894
R809 minus.n73 minus.n72 0.189894
R810 minus.n73 minus.n44 0.189894
R811 minus.n77 minus.n44 0.189894
R812 minus.n78 minus.n77 0.189894
R813 minus.n79 minus.n78 0.189894
R814 minus.n79 minus.n42 0.189894
R815 minus.n83 minus.n42 0.189894
R816 minus minus.n84 0.188
R817 drain_right.n13 drain_right.n11 68.0786
R818 drain_right.n7 drain_right.n5 68.0786
R819 drain_right.n2 drain_right.n0 68.0786
R820 drain_right.n13 drain_right.n12 67.1908
R821 drain_right.n15 drain_right.n14 67.1908
R822 drain_right.n17 drain_right.n16 67.1908
R823 drain_right.n19 drain_right.n18 67.1908
R824 drain_right.n21 drain_right.n20 67.1908
R825 drain_right.n7 drain_right.n6 67.1907
R826 drain_right.n9 drain_right.n8 67.1907
R827 drain_right.n4 drain_right.n3 67.1907
R828 drain_right.n2 drain_right.n1 67.1907
R829 drain_right drain_right.n10 30.7037
R830 drain_right drain_right.n21 6.54115
R831 drain_right.n5 drain_right.t8 3.3005
R832 drain_right.n5 drain_right.t7 3.3005
R833 drain_right.n6 drain_right.t21 3.3005
R834 drain_right.n6 drain_right.t2 3.3005
R835 drain_right.n8 drain_right.t15 3.3005
R836 drain_right.n8 drain_right.t20 3.3005
R837 drain_right.n3 drain_right.t10 3.3005
R838 drain_right.n3 drain_right.t17 3.3005
R839 drain_right.n1 drain_right.t13 3.3005
R840 drain_right.n1 drain_right.t12 3.3005
R841 drain_right.n0 drain_right.t6 3.3005
R842 drain_right.n0 drain_right.t4 3.3005
R843 drain_right.n11 drain_right.t23 3.3005
R844 drain_right.n11 drain_right.t11 3.3005
R845 drain_right.n12 drain_right.t1 3.3005
R846 drain_right.n12 drain_right.t14 3.3005
R847 drain_right.n14 drain_right.t0 3.3005
R848 drain_right.n14 drain_right.t16 3.3005
R849 drain_right.n16 drain_right.t3 3.3005
R850 drain_right.n16 drain_right.t18 3.3005
R851 drain_right.n18 drain_right.t5 3.3005
R852 drain_right.n18 drain_right.t19 3.3005
R853 drain_right.n20 drain_right.t9 3.3005
R854 drain_right.n20 drain_right.t22 3.3005
R855 drain_right.n9 drain_right.n7 0.888431
R856 drain_right.n4 drain_right.n2 0.888431
R857 drain_right.n21 drain_right.n19 0.888431
R858 drain_right.n19 drain_right.n17 0.888431
R859 drain_right.n17 drain_right.n15 0.888431
R860 drain_right.n15 drain_right.n13 0.888431
R861 drain_right.n10 drain_right.n9 0.389119
R862 drain_right.n10 drain_right.n4 0.389119
C0 minus plus 6.26978f
C1 source plus 8.534241f
C2 drain_left drain_right 1.87044f
C3 minus drain_right 7.86599f
C4 minus drain_left 0.174517f
C5 source drain_right 16.5602f
C6 source drain_left 16.5576f
C7 plus drain_right 0.498726f
C8 plus drain_left 8.20642f
C9 minus source 8.52023f
C10 drain_right a_n3394_n2088# 6.77301f
C11 drain_left a_n3394_n2088# 7.2476f
C12 source a_n3394_n2088# 5.950564f
C13 minus a_n3394_n2088# 13.194351f
C14 plus a_n3394_n2088# 14.814461f
C15 drain_right.t6 a_n3394_n2088# 0.128995f
C16 drain_right.t4 a_n3394_n2088# 0.128995f
C17 drain_right.n0 a_n3394_n2088# 1.08087f
C18 drain_right.t13 a_n3394_n2088# 0.128995f
C19 drain_right.t12 a_n3394_n2088# 0.128995f
C20 drain_right.n1 a_n3394_n2088# 1.07582f
C21 drain_right.n2 a_n3394_n2088# 0.758892f
C22 drain_right.t10 a_n3394_n2088# 0.128995f
C23 drain_right.t17 a_n3394_n2088# 0.128995f
C24 drain_right.n3 a_n3394_n2088# 1.07582f
C25 drain_right.n4 a_n3394_n2088# 0.334345f
C26 drain_right.t8 a_n3394_n2088# 0.128995f
C27 drain_right.t7 a_n3394_n2088# 0.128995f
C28 drain_right.n5 a_n3394_n2088# 1.08087f
C29 drain_right.t21 a_n3394_n2088# 0.128995f
C30 drain_right.t2 a_n3394_n2088# 0.128995f
C31 drain_right.n6 a_n3394_n2088# 1.07582f
C32 drain_right.n7 a_n3394_n2088# 0.758892f
C33 drain_right.t15 a_n3394_n2088# 0.128995f
C34 drain_right.t20 a_n3394_n2088# 0.128995f
C35 drain_right.n8 a_n3394_n2088# 1.07582f
C36 drain_right.n9 a_n3394_n2088# 0.334345f
C37 drain_right.n10 a_n3394_n2088# 1.37967f
C38 drain_right.t23 a_n3394_n2088# 0.128995f
C39 drain_right.t11 a_n3394_n2088# 0.128995f
C40 drain_right.n11 a_n3394_n2088# 1.08087f
C41 drain_right.t1 a_n3394_n2088# 0.128995f
C42 drain_right.t14 a_n3394_n2088# 0.128995f
C43 drain_right.n12 a_n3394_n2088# 1.07582f
C44 drain_right.n13 a_n3394_n2088# 0.758887f
C45 drain_right.t0 a_n3394_n2088# 0.128995f
C46 drain_right.t16 a_n3394_n2088# 0.128995f
C47 drain_right.n14 a_n3394_n2088# 1.07582f
C48 drain_right.n15 a_n3394_n2088# 0.376489f
C49 drain_right.t3 a_n3394_n2088# 0.128995f
C50 drain_right.t18 a_n3394_n2088# 0.128995f
C51 drain_right.n16 a_n3394_n2088# 1.07582f
C52 drain_right.n17 a_n3394_n2088# 0.376489f
C53 drain_right.t5 a_n3394_n2088# 0.128995f
C54 drain_right.t19 a_n3394_n2088# 0.128995f
C55 drain_right.n18 a_n3394_n2088# 1.07582f
C56 drain_right.n19 a_n3394_n2088# 0.376489f
C57 drain_right.t9 a_n3394_n2088# 0.128995f
C58 drain_right.t22 a_n3394_n2088# 0.128995f
C59 drain_right.n20 a_n3394_n2088# 1.07582f
C60 drain_right.n21 a_n3394_n2088# 0.617128f
C61 minus.n0 a_n3394_n2088# 0.039977f
C62 minus.n1 a_n3394_n2088# 0.009072f
C63 minus.t1 a_n3394_n2088# 0.487019f
C64 minus.n2 a_n3394_n2088# 0.039977f
C65 minus.n3 a_n3394_n2088# 0.009072f
C66 minus.t4 a_n3394_n2088# 0.487019f
C67 minus.n4 a_n3394_n2088# 0.039977f
C68 minus.n5 a_n3394_n2088# 0.009072f
C69 minus.t5 a_n3394_n2088# 0.487019f
C70 minus.n6 a_n3394_n2088# 0.039977f
C71 minus.n7 a_n3394_n2088# 0.009072f
C72 minus.t7 a_n3394_n2088# 0.487019f
C73 minus.n8 a_n3394_n2088# 0.039977f
C74 minus.n9 a_n3394_n2088# 0.009072f
C75 minus.t9 a_n3394_n2088# 0.487019f
C76 minus.t12 a_n3394_n2088# 0.507605f
C77 minus.t0 a_n3394_n2088# 0.487019f
C78 minus.n10 a_n3394_n2088# 0.233227f
C79 minus.n11 a_n3394_n2088# 0.206589f
C80 minus.n12 a_n3394_n2088# 0.172105f
C81 minus.n13 a_n3394_n2088# 0.039977f
C82 minus.n14 a_n3394_n2088# 0.225046f
C83 minus.n15 a_n3394_n2088# 0.009072f
C84 minus.t22 a_n3394_n2088# 0.487019f
C85 minus.n16 a_n3394_n2088# 0.225046f
C86 minus.n17 a_n3394_n2088# 0.039977f
C87 minus.n18 a_n3394_n2088# 0.039977f
C88 minus.n19 a_n3394_n2088# 0.039977f
C89 minus.n20 a_n3394_n2088# 0.225046f
C90 minus.n21 a_n3394_n2088# 0.009072f
C91 minus.t23 a_n3394_n2088# 0.487019f
C92 minus.n22 a_n3394_n2088# 0.225046f
C93 minus.n23 a_n3394_n2088# 0.039977f
C94 minus.n24 a_n3394_n2088# 0.039977f
C95 minus.n25 a_n3394_n2088# 0.039977f
C96 minus.n26 a_n3394_n2088# 0.225046f
C97 minus.n27 a_n3394_n2088# 0.009072f
C98 minus.t20 a_n3394_n2088# 0.487019f
C99 minus.n28 a_n3394_n2088# 0.225046f
C100 minus.n29 a_n3394_n2088# 0.039977f
C101 minus.n30 a_n3394_n2088# 0.039977f
C102 minus.n31 a_n3394_n2088# 0.039977f
C103 minus.n32 a_n3394_n2088# 0.225046f
C104 minus.n33 a_n3394_n2088# 0.009072f
C105 minus.t18 a_n3394_n2088# 0.487019f
C106 minus.n34 a_n3394_n2088# 0.225046f
C107 minus.n35 a_n3394_n2088# 0.039977f
C108 minus.n36 a_n3394_n2088# 0.039977f
C109 minus.n37 a_n3394_n2088# 0.039977f
C110 minus.n38 a_n3394_n2088# 0.225046f
C111 minus.n39 a_n3394_n2088# 0.009072f
C112 minus.t14 a_n3394_n2088# 0.487019f
C113 minus.n40 a_n3394_n2088# 0.225416f
C114 minus.n41 a_n3394_n2088# 1.50482f
C115 minus.n42 a_n3394_n2088# 0.039977f
C116 minus.n43 a_n3394_n2088# 0.009072f
C117 minus.n44 a_n3394_n2088# 0.039977f
C118 minus.n45 a_n3394_n2088# 0.009072f
C119 minus.n46 a_n3394_n2088# 0.039977f
C120 minus.n47 a_n3394_n2088# 0.009072f
C121 minus.n48 a_n3394_n2088# 0.039977f
C122 minus.n49 a_n3394_n2088# 0.009072f
C123 minus.n50 a_n3394_n2088# 0.039977f
C124 minus.n51 a_n3394_n2088# 0.009072f
C125 minus.t17 a_n3394_n2088# 0.507605f
C126 minus.t19 a_n3394_n2088# 0.487019f
C127 minus.n52 a_n3394_n2088# 0.233227f
C128 minus.n53 a_n3394_n2088# 0.206589f
C129 minus.n54 a_n3394_n2088# 0.172105f
C130 minus.n55 a_n3394_n2088# 0.039977f
C131 minus.t10 a_n3394_n2088# 0.487019f
C132 minus.n56 a_n3394_n2088# 0.225046f
C133 minus.n57 a_n3394_n2088# 0.009072f
C134 minus.t11 a_n3394_n2088# 0.487019f
C135 minus.n58 a_n3394_n2088# 0.225046f
C136 minus.n59 a_n3394_n2088# 0.039977f
C137 minus.n60 a_n3394_n2088# 0.039977f
C138 minus.n61 a_n3394_n2088# 0.039977f
C139 minus.t13 a_n3394_n2088# 0.487019f
C140 minus.n62 a_n3394_n2088# 0.225046f
C141 minus.n63 a_n3394_n2088# 0.009072f
C142 minus.t6 a_n3394_n2088# 0.487019f
C143 minus.n64 a_n3394_n2088# 0.225046f
C144 minus.n65 a_n3394_n2088# 0.039977f
C145 minus.n66 a_n3394_n2088# 0.039977f
C146 minus.n67 a_n3394_n2088# 0.039977f
C147 minus.t8 a_n3394_n2088# 0.487019f
C148 minus.n68 a_n3394_n2088# 0.225046f
C149 minus.n69 a_n3394_n2088# 0.009072f
C150 minus.t3 a_n3394_n2088# 0.487019f
C151 minus.n70 a_n3394_n2088# 0.225046f
C152 minus.n71 a_n3394_n2088# 0.039977f
C153 minus.n72 a_n3394_n2088# 0.039977f
C154 minus.n73 a_n3394_n2088# 0.039977f
C155 minus.t2 a_n3394_n2088# 0.487019f
C156 minus.n74 a_n3394_n2088# 0.225046f
C157 minus.n75 a_n3394_n2088# 0.009072f
C158 minus.t21 a_n3394_n2088# 0.487019f
C159 minus.n76 a_n3394_n2088# 0.225046f
C160 minus.n77 a_n3394_n2088# 0.039977f
C161 minus.n78 a_n3394_n2088# 0.039977f
C162 minus.n79 a_n3394_n2088# 0.039977f
C163 minus.t15 a_n3394_n2088# 0.487019f
C164 minus.n80 a_n3394_n2088# 0.225046f
C165 minus.n81 a_n3394_n2088# 0.009072f
C166 minus.t16 a_n3394_n2088# 0.487019f
C167 minus.n82 a_n3394_n2088# 0.225416f
C168 minus.n83 a_n3394_n2088# 0.278038f
C169 minus.n84 a_n3394_n2088# 1.81514f
C170 drain_left.t12 a_n3394_n2088# 0.130009f
C171 drain_left.t13 a_n3394_n2088# 0.130009f
C172 drain_left.n0 a_n3394_n2088# 1.08937f
C173 drain_left.t14 a_n3394_n2088# 0.130009f
C174 drain_left.t15 a_n3394_n2088# 0.130009f
C175 drain_left.n1 a_n3394_n2088# 1.08428f
C176 drain_left.n2 a_n3394_n2088# 0.764862f
C177 drain_left.t10 a_n3394_n2088# 0.130009f
C178 drain_left.t1 a_n3394_n2088# 0.130009f
C179 drain_left.n3 a_n3394_n2088# 1.08428f
C180 drain_left.n4 a_n3394_n2088# 0.336975f
C181 drain_left.t7 a_n3394_n2088# 0.130009f
C182 drain_left.t8 a_n3394_n2088# 0.130009f
C183 drain_left.n5 a_n3394_n2088# 1.08937f
C184 drain_left.t21 a_n3394_n2088# 0.130009f
C185 drain_left.t11 a_n3394_n2088# 0.130009f
C186 drain_left.n6 a_n3394_n2088# 1.08428f
C187 drain_left.n7 a_n3394_n2088# 0.764862f
C188 drain_left.t2 a_n3394_n2088# 0.130009f
C189 drain_left.t19 a_n3394_n2088# 0.130009f
C190 drain_left.n8 a_n3394_n2088# 1.08428f
C191 drain_left.n9 a_n3394_n2088# 0.336975f
C192 drain_left.n10 a_n3394_n2088# 1.44495f
C193 drain_left.t16 a_n3394_n2088# 0.130009f
C194 drain_left.t3 a_n3394_n2088# 0.130009f
C195 drain_left.n11 a_n3394_n2088# 1.08938f
C196 drain_left.t20 a_n3394_n2088# 0.130009f
C197 drain_left.t6 a_n3394_n2088# 0.130009f
C198 drain_left.n12 a_n3394_n2088# 1.08428f
C199 drain_left.n13 a_n3394_n2088# 0.764852f
C200 drain_left.t17 a_n3394_n2088# 0.130009f
C201 drain_left.t4 a_n3394_n2088# 0.130009f
C202 drain_left.n14 a_n3394_n2088# 1.08428f
C203 drain_left.n15 a_n3394_n2088# 0.379451f
C204 drain_left.t22 a_n3394_n2088# 0.130009f
C205 drain_left.t9 a_n3394_n2088# 0.130009f
C206 drain_left.n16 a_n3394_n2088# 1.08428f
C207 drain_left.n17 a_n3394_n2088# 0.379451f
C208 drain_left.t0 a_n3394_n2088# 0.130009f
C209 drain_left.t18 a_n3394_n2088# 0.130009f
C210 drain_left.n18 a_n3394_n2088# 1.08428f
C211 drain_left.n19 a_n3394_n2088# 0.379451f
C212 drain_left.t5 a_n3394_n2088# 0.130009f
C213 drain_left.t23 a_n3394_n2088# 0.130009f
C214 drain_left.n20 a_n3394_n2088# 1.08428f
C215 drain_left.n21 a_n3394_n2088# 0.621988f
C216 source.n0 a_n3394_n2088# 0.037578f
C217 source.n1 a_n3394_n2088# 0.026735f
C218 source.n2 a_n3394_n2088# 0.014366f
C219 source.n3 a_n3394_n2088# 0.033956f
C220 source.n4 a_n3394_n2088# 0.015211f
C221 source.n5 a_n3394_n2088# 0.026735f
C222 source.n6 a_n3394_n2088# 0.014366f
C223 source.n7 a_n3394_n2088# 0.033956f
C224 source.n8 a_n3394_n2088# 0.015211f
C225 source.n9 a_n3394_n2088# 0.114406f
C226 source.t39 a_n3394_n2088# 0.055344f
C227 source.n10 a_n3394_n2088# 0.025467f
C228 source.n11 a_n3394_n2088# 0.020058f
C229 source.n12 a_n3394_n2088# 0.014366f
C230 source.n13 a_n3394_n2088# 0.636127f
C231 source.n14 a_n3394_n2088# 0.026735f
C232 source.n15 a_n3394_n2088# 0.014366f
C233 source.n16 a_n3394_n2088# 0.015211f
C234 source.n17 a_n3394_n2088# 0.033956f
C235 source.n18 a_n3394_n2088# 0.033956f
C236 source.n19 a_n3394_n2088# 0.015211f
C237 source.n20 a_n3394_n2088# 0.014366f
C238 source.n21 a_n3394_n2088# 0.026735f
C239 source.n22 a_n3394_n2088# 0.026735f
C240 source.n23 a_n3394_n2088# 0.014366f
C241 source.n24 a_n3394_n2088# 0.015211f
C242 source.n25 a_n3394_n2088# 0.033956f
C243 source.n26 a_n3394_n2088# 0.073509f
C244 source.n27 a_n3394_n2088# 0.015211f
C245 source.n28 a_n3394_n2088# 0.014366f
C246 source.n29 a_n3394_n2088# 0.061796f
C247 source.n30 a_n3394_n2088# 0.041131f
C248 source.n31 a_n3394_n2088# 0.698406f
C249 source.t27 a_n3394_n2088# 0.12676f
C250 source.t37 a_n3394_n2088# 0.12676f
C251 source.n32 a_n3394_n2088# 0.987213f
C252 source.n33 a_n3394_n2088# 0.403594f
C253 source.t32 a_n3394_n2088# 0.12676f
C254 source.t23 a_n3394_n2088# 0.12676f
C255 source.n34 a_n3394_n2088# 0.987213f
C256 source.n35 a_n3394_n2088# 0.403594f
C257 source.t46 a_n3394_n2088# 0.12676f
C258 source.t41 a_n3394_n2088# 0.12676f
C259 source.n36 a_n3394_n2088# 0.987213f
C260 source.n37 a_n3394_n2088# 0.403594f
C261 source.t25 a_n3394_n2088# 0.12676f
C262 source.t30 a_n3394_n2088# 0.12676f
C263 source.n38 a_n3394_n2088# 0.987213f
C264 source.n39 a_n3394_n2088# 0.403594f
C265 source.t38 a_n3394_n2088# 0.12676f
C266 source.t24 a_n3394_n2088# 0.12676f
C267 source.n40 a_n3394_n2088# 0.987213f
C268 source.n41 a_n3394_n2088# 0.403594f
C269 source.n42 a_n3394_n2088# 0.037578f
C270 source.n43 a_n3394_n2088# 0.026735f
C271 source.n44 a_n3394_n2088# 0.014366f
C272 source.n45 a_n3394_n2088# 0.033956f
C273 source.n46 a_n3394_n2088# 0.015211f
C274 source.n47 a_n3394_n2088# 0.026735f
C275 source.n48 a_n3394_n2088# 0.014366f
C276 source.n49 a_n3394_n2088# 0.033956f
C277 source.n50 a_n3394_n2088# 0.015211f
C278 source.n51 a_n3394_n2088# 0.114406f
C279 source.t28 a_n3394_n2088# 0.055344f
C280 source.n52 a_n3394_n2088# 0.025467f
C281 source.n53 a_n3394_n2088# 0.020058f
C282 source.n54 a_n3394_n2088# 0.014366f
C283 source.n55 a_n3394_n2088# 0.636127f
C284 source.n56 a_n3394_n2088# 0.026735f
C285 source.n57 a_n3394_n2088# 0.014366f
C286 source.n58 a_n3394_n2088# 0.015211f
C287 source.n59 a_n3394_n2088# 0.033956f
C288 source.n60 a_n3394_n2088# 0.033956f
C289 source.n61 a_n3394_n2088# 0.015211f
C290 source.n62 a_n3394_n2088# 0.014366f
C291 source.n63 a_n3394_n2088# 0.026735f
C292 source.n64 a_n3394_n2088# 0.026735f
C293 source.n65 a_n3394_n2088# 0.014366f
C294 source.n66 a_n3394_n2088# 0.015211f
C295 source.n67 a_n3394_n2088# 0.033956f
C296 source.n68 a_n3394_n2088# 0.073509f
C297 source.n69 a_n3394_n2088# 0.015211f
C298 source.n70 a_n3394_n2088# 0.014366f
C299 source.n71 a_n3394_n2088# 0.061796f
C300 source.n72 a_n3394_n2088# 0.041131f
C301 source.n73 a_n3394_n2088# 0.139798f
C302 source.n74 a_n3394_n2088# 0.037578f
C303 source.n75 a_n3394_n2088# 0.026735f
C304 source.n76 a_n3394_n2088# 0.014366f
C305 source.n77 a_n3394_n2088# 0.033956f
C306 source.n78 a_n3394_n2088# 0.015211f
C307 source.n79 a_n3394_n2088# 0.026735f
C308 source.n80 a_n3394_n2088# 0.014366f
C309 source.n81 a_n3394_n2088# 0.033956f
C310 source.n82 a_n3394_n2088# 0.015211f
C311 source.n83 a_n3394_n2088# 0.114406f
C312 source.t9 a_n3394_n2088# 0.055344f
C313 source.n84 a_n3394_n2088# 0.025467f
C314 source.n85 a_n3394_n2088# 0.020058f
C315 source.n86 a_n3394_n2088# 0.014366f
C316 source.n87 a_n3394_n2088# 0.636127f
C317 source.n88 a_n3394_n2088# 0.026735f
C318 source.n89 a_n3394_n2088# 0.014366f
C319 source.n90 a_n3394_n2088# 0.015211f
C320 source.n91 a_n3394_n2088# 0.033956f
C321 source.n92 a_n3394_n2088# 0.033956f
C322 source.n93 a_n3394_n2088# 0.015211f
C323 source.n94 a_n3394_n2088# 0.014366f
C324 source.n95 a_n3394_n2088# 0.026735f
C325 source.n96 a_n3394_n2088# 0.026735f
C326 source.n97 a_n3394_n2088# 0.014366f
C327 source.n98 a_n3394_n2088# 0.015211f
C328 source.n99 a_n3394_n2088# 0.033956f
C329 source.n100 a_n3394_n2088# 0.073509f
C330 source.n101 a_n3394_n2088# 0.015211f
C331 source.n102 a_n3394_n2088# 0.014366f
C332 source.n103 a_n3394_n2088# 0.061796f
C333 source.n104 a_n3394_n2088# 0.041131f
C334 source.n105 a_n3394_n2088# 0.139798f
C335 source.t0 a_n3394_n2088# 0.12676f
C336 source.t12 a_n3394_n2088# 0.12676f
C337 source.n106 a_n3394_n2088# 0.987213f
C338 source.n107 a_n3394_n2088# 0.403594f
C339 source.t14 a_n3394_n2088# 0.12676f
C340 source.t3 a_n3394_n2088# 0.12676f
C341 source.n108 a_n3394_n2088# 0.987213f
C342 source.n109 a_n3394_n2088# 0.403594f
C343 source.t13 a_n3394_n2088# 0.12676f
C344 source.t47 a_n3394_n2088# 0.12676f
C345 source.n110 a_n3394_n2088# 0.987213f
C346 source.n111 a_n3394_n2088# 0.403594f
C347 source.t22 a_n3394_n2088# 0.12676f
C348 source.t4 a_n3394_n2088# 0.12676f
C349 source.n112 a_n3394_n2088# 0.987213f
C350 source.n113 a_n3394_n2088# 0.403594f
C351 source.t15 a_n3394_n2088# 0.12676f
C352 source.t7 a_n3394_n2088# 0.12676f
C353 source.n114 a_n3394_n2088# 0.987213f
C354 source.n115 a_n3394_n2088# 0.403594f
C355 source.n116 a_n3394_n2088# 0.037578f
C356 source.n117 a_n3394_n2088# 0.026735f
C357 source.n118 a_n3394_n2088# 0.014366f
C358 source.n119 a_n3394_n2088# 0.033956f
C359 source.n120 a_n3394_n2088# 0.015211f
C360 source.n121 a_n3394_n2088# 0.026735f
C361 source.n122 a_n3394_n2088# 0.014366f
C362 source.n123 a_n3394_n2088# 0.033956f
C363 source.n124 a_n3394_n2088# 0.015211f
C364 source.n125 a_n3394_n2088# 0.114406f
C365 source.t8 a_n3394_n2088# 0.055344f
C366 source.n126 a_n3394_n2088# 0.025467f
C367 source.n127 a_n3394_n2088# 0.020058f
C368 source.n128 a_n3394_n2088# 0.014366f
C369 source.n129 a_n3394_n2088# 0.636127f
C370 source.n130 a_n3394_n2088# 0.026735f
C371 source.n131 a_n3394_n2088# 0.014366f
C372 source.n132 a_n3394_n2088# 0.015211f
C373 source.n133 a_n3394_n2088# 0.033956f
C374 source.n134 a_n3394_n2088# 0.033956f
C375 source.n135 a_n3394_n2088# 0.015211f
C376 source.n136 a_n3394_n2088# 0.014366f
C377 source.n137 a_n3394_n2088# 0.026735f
C378 source.n138 a_n3394_n2088# 0.026735f
C379 source.n139 a_n3394_n2088# 0.014366f
C380 source.n140 a_n3394_n2088# 0.015211f
C381 source.n141 a_n3394_n2088# 0.033956f
C382 source.n142 a_n3394_n2088# 0.073509f
C383 source.n143 a_n3394_n2088# 0.015211f
C384 source.n144 a_n3394_n2088# 0.014366f
C385 source.n145 a_n3394_n2088# 0.061796f
C386 source.n146 a_n3394_n2088# 0.041131f
C387 source.n147 a_n3394_n2088# 1.05116f
C388 source.n148 a_n3394_n2088# 0.037578f
C389 source.n149 a_n3394_n2088# 0.026735f
C390 source.n150 a_n3394_n2088# 0.014366f
C391 source.n151 a_n3394_n2088# 0.033956f
C392 source.n152 a_n3394_n2088# 0.015211f
C393 source.n153 a_n3394_n2088# 0.026735f
C394 source.n154 a_n3394_n2088# 0.014366f
C395 source.n155 a_n3394_n2088# 0.033956f
C396 source.n156 a_n3394_n2088# 0.015211f
C397 source.n157 a_n3394_n2088# 0.114406f
C398 source.t33 a_n3394_n2088# 0.055344f
C399 source.n158 a_n3394_n2088# 0.025467f
C400 source.n159 a_n3394_n2088# 0.020058f
C401 source.n160 a_n3394_n2088# 0.014366f
C402 source.n161 a_n3394_n2088# 0.636127f
C403 source.n162 a_n3394_n2088# 0.026735f
C404 source.n163 a_n3394_n2088# 0.014366f
C405 source.n164 a_n3394_n2088# 0.015211f
C406 source.n165 a_n3394_n2088# 0.033956f
C407 source.n166 a_n3394_n2088# 0.033956f
C408 source.n167 a_n3394_n2088# 0.015211f
C409 source.n168 a_n3394_n2088# 0.014366f
C410 source.n169 a_n3394_n2088# 0.026735f
C411 source.n170 a_n3394_n2088# 0.026735f
C412 source.n171 a_n3394_n2088# 0.014366f
C413 source.n172 a_n3394_n2088# 0.015211f
C414 source.n173 a_n3394_n2088# 0.033956f
C415 source.n174 a_n3394_n2088# 0.073509f
C416 source.n175 a_n3394_n2088# 0.015211f
C417 source.n176 a_n3394_n2088# 0.014366f
C418 source.n177 a_n3394_n2088# 0.061796f
C419 source.n178 a_n3394_n2088# 0.041131f
C420 source.n179 a_n3394_n2088# 1.05116f
C421 source.t31 a_n3394_n2088# 0.12676f
C422 source.t44 a_n3394_n2088# 0.12676f
C423 source.n180 a_n3394_n2088# 0.987207f
C424 source.n181 a_n3394_n2088# 0.403601f
C425 source.t43 a_n3394_n2088# 0.12676f
C426 source.t45 a_n3394_n2088# 0.12676f
C427 source.n182 a_n3394_n2088# 0.987207f
C428 source.n183 a_n3394_n2088# 0.403601f
C429 source.t35 a_n3394_n2088# 0.12676f
C430 source.t40 a_n3394_n2088# 0.12676f
C431 source.n184 a_n3394_n2088# 0.987207f
C432 source.n185 a_n3394_n2088# 0.403601f
C433 source.t42 a_n3394_n2088# 0.12676f
C434 source.t26 a_n3394_n2088# 0.12676f
C435 source.n186 a_n3394_n2088# 0.987207f
C436 source.n187 a_n3394_n2088# 0.403601f
C437 source.t36 a_n3394_n2088# 0.12676f
C438 source.t29 a_n3394_n2088# 0.12676f
C439 source.n188 a_n3394_n2088# 0.987207f
C440 source.n189 a_n3394_n2088# 0.403601f
C441 source.n190 a_n3394_n2088# 0.037578f
C442 source.n191 a_n3394_n2088# 0.026735f
C443 source.n192 a_n3394_n2088# 0.014366f
C444 source.n193 a_n3394_n2088# 0.033956f
C445 source.n194 a_n3394_n2088# 0.015211f
C446 source.n195 a_n3394_n2088# 0.026735f
C447 source.n196 a_n3394_n2088# 0.014366f
C448 source.n197 a_n3394_n2088# 0.033956f
C449 source.n198 a_n3394_n2088# 0.015211f
C450 source.n199 a_n3394_n2088# 0.114406f
C451 source.t34 a_n3394_n2088# 0.055344f
C452 source.n200 a_n3394_n2088# 0.025467f
C453 source.n201 a_n3394_n2088# 0.020058f
C454 source.n202 a_n3394_n2088# 0.014366f
C455 source.n203 a_n3394_n2088# 0.636127f
C456 source.n204 a_n3394_n2088# 0.026735f
C457 source.n205 a_n3394_n2088# 0.014366f
C458 source.n206 a_n3394_n2088# 0.015211f
C459 source.n207 a_n3394_n2088# 0.033956f
C460 source.n208 a_n3394_n2088# 0.033956f
C461 source.n209 a_n3394_n2088# 0.015211f
C462 source.n210 a_n3394_n2088# 0.014366f
C463 source.n211 a_n3394_n2088# 0.026735f
C464 source.n212 a_n3394_n2088# 0.026735f
C465 source.n213 a_n3394_n2088# 0.014366f
C466 source.n214 a_n3394_n2088# 0.015211f
C467 source.n215 a_n3394_n2088# 0.033956f
C468 source.n216 a_n3394_n2088# 0.073509f
C469 source.n217 a_n3394_n2088# 0.015211f
C470 source.n218 a_n3394_n2088# 0.014366f
C471 source.n219 a_n3394_n2088# 0.061796f
C472 source.n220 a_n3394_n2088# 0.041131f
C473 source.n221 a_n3394_n2088# 0.139798f
C474 source.n222 a_n3394_n2088# 0.037578f
C475 source.n223 a_n3394_n2088# 0.026735f
C476 source.n224 a_n3394_n2088# 0.014366f
C477 source.n225 a_n3394_n2088# 0.033956f
C478 source.n226 a_n3394_n2088# 0.015211f
C479 source.n227 a_n3394_n2088# 0.026735f
C480 source.n228 a_n3394_n2088# 0.014366f
C481 source.n229 a_n3394_n2088# 0.033956f
C482 source.n230 a_n3394_n2088# 0.015211f
C483 source.n231 a_n3394_n2088# 0.114406f
C484 source.t18 a_n3394_n2088# 0.055344f
C485 source.n232 a_n3394_n2088# 0.025467f
C486 source.n233 a_n3394_n2088# 0.020058f
C487 source.n234 a_n3394_n2088# 0.014366f
C488 source.n235 a_n3394_n2088# 0.636127f
C489 source.n236 a_n3394_n2088# 0.026735f
C490 source.n237 a_n3394_n2088# 0.014366f
C491 source.n238 a_n3394_n2088# 0.015211f
C492 source.n239 a_n3394_n2088# 0.033956f
C493 source.n240 a_n3394_n2088# 0.033956f
C494 source.n241 a_n3394_n2088# 0.015211f
C495 source.n242 a_n3394_n2088# 0.014366f
C496 source.n243 a_n3394_n2088# 0.026735f
C497 source.n244 a_n3394_n2088# 0.026735f
C498 source.n245 a_n3394_n2088# 0.014366f
C499 source.n246 a_n3394_n2088# 0.015211f
C500 source.n247 a_n3394_n2088# 0.033956f
C501 source.n248 a_n3394_n2088# 0.073509f
C502 source.n249 a_n3394_n2088# 0.015211f
C503 source.n250 a_n3394_n2088# 0.014366f
C504 source.n251 a_n3394_n2088# 0.061796f
C505 source.n252 a_n3394_n2088# 0.041131f
C506 source.n253 a_n3394_n2088# 0.139798f
C507 source.t17 a_n3394_n2088# 0.12676f
C508 source.t19 a_n3394_n2088# 0.12676f
C509 source.n254 a_n3394_n2088# 0.987207f
C510 source.n255 a_n3394_n2088# 0.403601f
C511 source.t1 a_n3394_n2088# 0.12676f
C512 source.t5 a_n3394_n2088# 0.12676f
C513 source.n256 a_n3394_n2088# 0.987207f
C514 source.n257 a_n3394_n2088# 0.403601f
C515 source.t2 a_n3394_n2088# 0.12676f
C516 source.t16 a_n3394_n2088# 0.12676f
C517 source.n258 a_n3394_n2088# 0.987207f
C518 source.n259 a_n3394_n2088# 0.403601f
C519 source.t11 a_n3394_n2088# 0.12676f
C520 source.t10 a_n3394_n2088# 0.12676f
C521 source.n260 a_n3394_n2088# 0.987207f
C522 source.n261 a_n3394_n2088# 0.403601f
C523 source.t20 a_n3394_n2088# 0.12676f
C524 source.t6 a_n3394_n2088# 0.12676f
C525 source.n262 a_n3394_n2088# 0.987207f
C526 source.n263 a_n3394_n2088# 0.403601f
C527 source.n264 a_n3394_n2088# 0.037578f
C528 source.n265 a_n3394_n2088# 0.026735f
C529 source.n266 a_n3394_n2088# 0.014366f
C530 source.n267 a_n3394_n2088# 0.033956f
C531 source.n268 a_n3394_n2088# 0.015211f
C532 source.n269 a_n3394_n2088# 0.026735f
C533 source.n270 a_n3394_n2088# 0.014366f
C534 source.n271 a_n3394_n2088# 0.033956f
C535 source.n272 a_n3394_n2088# 0.015211f
C536 source.n273 a_n3394_n2088# 0.114406f
C537 source.t21 a_n3394_n2088# 0.055344f
C538 source.n274 a_n3394_n2088# 0.025467f
C539 source.n275 a_n3394_n2088# 0.020058f
C540 source.n276 a_n3394_n2088# 0.014366f
C541 source.n277 a_n3394_n2088# 0.636127f
C542 source.n278 a_n3394_n2088# 0.026735f
C543 source.n279 a_n3394_n2088# 0.014366f
C544 source.n280 a_n3394_n2088# 0.015211f
C545 source.n281 a_n3394_n2088# 0.033956f
C546 source.n282 a_n3394_n2088# 0.033956f
C547 source.n283 a_n3394_n2088# 0.015211f
C548 source.n284 a_n3394_n2088# 0.014366f
C549 source.n285 a_n3394_n2088# 0.026735f
C550 source.n286 a_n3394_n2088# 0.026735f
C551 source.n287 a_n3394_n2088# 0.014366f
C552 source.n288 a_n3394_n2088# 0.015211f
C553 source.n289 a_n3394_n2088# 0.033956f
C554 source.n290 a_n3394_n2088# 0.073509f
C555 source.n291 a_n3394_n2088# 0.015211f
C556 source.n292 a_n3394_n2088# 0.014366f
C557 source.n293 a_n3394_n2088# 0.061796f
C558 source.n294 a_n3394_n2088# 0.041131f
C559 source.n295 a_n3394_n2088# 0.314189f
C560 source.n296 a_n3394_n2088# 1.10874f
C561 plus.n0 a_n3394_n2088# 0.040651f
C562 plus.t0 a_n3394_n2088# 0.495219f
C563 plus.t18 a_n3394_n2088# 0.495219f
C564 plus.n1 a_n3394_n2088# 0.040651f
C565 plus.t5 a_n3394_n2088# 0.495219f
C566 plus.n2 a_n3394_n2088# 0.228836f
C567 plus.n3 a_n3394_n2088# 0.040651f
C568 plus.t23 a_n3394_n2088# 0.495219f
C569 plus.t14 a_n3394_n2088# 0.495219f
C570 plus.n4 a_n3394_n2088# 0.228836f
C571 plus.n5 a_n3394_n2088# 0.040651f
C572 plus.t1 a_n3394_n2088# 0.495219f
C573 plus.t19 a_n3394_n2088# 0.495219f
C574 plus.n6 a_n3394_n2088# 0.228836f
C575 plus.n7 a_n3394_n2088# 0.040651f
C576 plus.t6 a_n3394_n2088# 0.495219f
C577 plus.t17 a_n3394_n2088# 0.495219f
C578 plus.n8 a_n3394_n2088# 0.228836f
C579 plus.n9 a_n3394_n2088# 0.040651f
C580 plus.t3 a_n3394_n2088# 0.495219f
C581 plus.t20 a_n3394_n2088# 0.495219f
C582 plus.n10 a_n3394_n2088# 0.237154f
C583 plus.t7 a_n3394_n2088# 0.516151f
C584 plus.n11 a_n3394_n2088# 0.210067f
C585 plus.n12 a_n3394_n2088# 0.175003f
C586 plus.n13 a_n3394_n2088# 0.009224f
C587 plus.n14 a_n3394_n2088# 0.228836f
C588 plus.n15 a_n3394_n2088# 0.009224f
C589 plus.n16 a_n3394_n2088# 0.040651f
C590 plus.n17 a_n3394_n2088# 0.040651f
C591 plus.n18 a_n3394_n2088# 0.040651f
C592 plus.n19 a_n3394_n2088# 0.009224f
C593 plus.n20 a_n3394_n2088# 0.228836f
C594 plus.n21 a_n3394_n2088# 0.009224f
C595 plus.n22 a_n3394_n2088# 0.040651f
C596 plus.n23 a_n3394_n2088# 0.040651f
C597 plus.n24 a_n3394_n2088# 0.040651f
C598 plus.n25 a_n3394_n2088# 0.009224f
C599 plus.n26 a_n3394_n2088# 0.228836f
C600 plus.n27 a_n3394_n2088# 0.009224f
C601 plus.n28 a_n3394_n2088# 0.040651f
C602 plus.n29 a_n3394_n2088# 0.040651f
C603 plus.n30 a_n3394_n2088# 0.040651f
C604 plus.n31 a_n3394_n2088# 0.009224f
C605 plus.n32 a_n3394_n2088# 0.228836f
C606 plus.n33 a_n3394_n2088# 0.009224f
C607 plus.n34 a_n3394_n2088# 0.040651f
C608 plus.n35 a_n3394_n2088# 0.040651f
C609 plus.n36 a_n3394_n2088# 0.040651f
C610 plus.n37 a_n3394_n2088# 0.009224f
C611 plus.n38 a_n3394_n2088# 0.228836f
C612 plus.n39 a_n3394_n2088# 0.009224f
C613 plus.n40 a_n3394_n2088# 0.229212f
C614 plus.n41 a_n3394_n2088# 0.366059f
C615 plus.n42 a_n3394_n2088# 0.040651f
C616 plus.t11 a_n3394_n2088# 0.495219f
C617 plus.n43 a_n3394_n2088# 0.040651f
C618 plus.t10 a_n3394_n2088# 0.495219f
C619 plus.t9 a_n3394_n2088# 0.495219f
C620 plus.n44 a_n3394_n2088# 0.228836f
C621 plus.n45 a_n3394_n2088# 0.040651f
C622 plus.t8 a_n3394_n2088# 0.495219f
C623 plus.t13 a_n3394_n2088# 0.495219f
C624 plus.n46 a_n3394_n2088# 0.228836f
C625 plus.n47 a_n3394_n2088# 0.040651f
C626 plus.t22 a_n3394_n2088# 0.495219f
C627 plus.t21 a_n3394_n2088# 0.495219f
C628 plus.n48 a_n3394_n2088# 0.228836f
C629 plus.n49 a_n3394_n2088# 0.040651f
C630 plus.t4 a_n3394_n2088# 0.495219f
C631 plus.t2 a_n3394_n2088# 0.495219f
C632 plus.n50 a_n3394_n2088# 0.228836f
C633 plus.n51 a_n3394_n2088# 0.040651f
C634 plus.t12 a_n3394_n2088# 0.495219f
C635 plus.t16 a_n3394_n2088# 0.495219f
C636 plus.n52 a_n3394_n2088# 0.237154f
C637 plus.t15 a_n3394_n2088# 0.516151f
C638 plus.n53 a_n3394_n2088# 0.210067f
C639 plus.n54 a_n3394_n2088# 0.175003f
C640 plus.n55 a_n3394_n2088# 0.009224f
C641 plus.n56 a_n3394_n2088# 0.228836f
C642 plus.n57 a_n3394_n2088# 0.009224f
C643 plus.n58 a_n3394_n2088# 0.040651f
C644 plus.n59 a_n3394_n2088# 0.040651f
C645 plus.n60 a_n3394_n2088# 0.040651f
C646 plus.n61 a_n3394_n2088# 0.009224f
C647 plus.n62 a_n3394_n2088# 0.228836f
C648 plus.n63 a_n3394_n2088# 0.009224f
C649 plus.n64 a_n3394_n2088# 0.040651f
C650 plus.n65 a_n3394_n2088# 0.040651f
C651 plus.n66 a_n3394_n2088# 0.040651f
C652 plus.n67 a_n3394_n2088# 0.009224f
C653 plus.n68 a_n3394_n2088# 0.228836f
C654 plus.n69 a_n3394_n2088# 0.009224f
C655 plus.n70 a_n3394_n2088# 0.040651f
C656 plus.n71 a_n3394_n2088# 0.040651f
C657 plus.n72 a_n3394_n2088# 0.040651f
C658 plus.n73 a_n3394_n2088# 0.009224f
C659 plus.n74 a_n3394_n2088# 0.228836f
C660 plus.n75 a_n3394_n2088# 0.009224f
C661 plus.n76 a_n3394_n2088# 0.040651f
C662 plus.n77 a_n3394_n2088# 0.040651f
C663 plus.n78 a_n3394_n2088# 0.040651f
C664 plus.n79 a_n3394_n2088# 0.009224f
C665 plus.n80 a_n3394_n2088# 0.228836f
C666 plus.n81 a_n3394_n2088# 0.009224f
C667 plus.n82 a_n3394_n2088# 0.229212f
C668 plus.n83 a_n3394_n2088# 1.39065f
.ends

