* NGSPICE file created from diffpair384.ext - technology: sky130A

.subckt diffpair384 minus drain_right drain_left source plus
X0 drain_left.t9 plus.t0 source.t13 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X1 source.t1 minus.t0 drain_right.t9 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X2 a_n1952_n2688# a_n1952_n2688# a_n1952_n2688# a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.7
X3 drain_left.t8 plus.t1 source.t15 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X4 drain_left.t7 plus.t2 source.t12 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X5 source.t14 plus.t3 drain_left.t6 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X6 drain_left.t5 plus.t4 source.t9 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X7 drain_right.t8 minus.t1 source.t6 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X8 a_n1952_n2688# a_n1952_n2688# a_n1952_n2688# a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X9 drain_left.t4 plus.t5 source.t16 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X10 drain_right.t7 minus.t2 source.t0 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X11 source.t17 plus.t6 drain_left.t3 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X12 drain_right.t6 minus.t3 source.t19 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X13 source.t11 plus.t7 drain_left.t2 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X14 drain_left.t1 plus.t8 source.t10 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X15 drain_right.t5 minus.t4 source.t5 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X16 source.t18 plus.t9 drain_left.t0 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X17 source.t4 minus.t5 drain_right.t4 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X18 a_n1952_n2688# a_n1952_n2688# a_n1952_n2688# a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X19 a_n1952_n2688# a_n1952_n2688# a_n1952_n2688# a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X20 drain_right.t3 minus.t6 source.t2 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X21 source.t8 minus.t7 drain_right.t2 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X22 source.t3 minus.t8 drain_right.t1 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X23 drain_right.t0 minus.t9 source.t7 a_n1952_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
R0 plus.n3 plus.t2 388.724
R1 plus.n17 plus.t8 388.724
R2 plus.n12 plus.t1 365.976
R3 plus.n10 plus.t6 365.976
R4 plus.n2 plus.t0 365.976
R5 plus.n4 plus.t7 365.976
R6 plus.n26 plus.t4 365.976
R7 plus.n24 plus.t3 365.976
R8 plus.n16 plus.t5 365.976
R9 plus.n18 plus.t9 365.976
R10 plus.n6 plus.n5 161.3
R11 plus.n7 plus.n2 161.3
R12 plus.n9 plus.n8 161.3
R13 plus.n10 plus.n1 161.3
R14 plus.n11 plus.n0 161.3
R15 plus.n13 plus.n12 161.3
R16 plus.n20 plus.n19 161.3
R17 plus.n21 plus.n16 161.3
R18 plus.n23 plus.n22 161.3
R19 plus.n24 plus.n15 161.3
R20 plus.n25 plus.n14 161.3
R21 plus.n27 plus.n26 161.3
R22 plus.n6 plus.n3 44.8741
R23 plus.n20 plus.n17 44.8741
R24 plus.n12 plus.n11 30.6732
R25 plus.n26 plus.n25 30.6732
R26 plus plus.n27 29.3986
R27 plus.n10 plus.n9 26.2914
R28 plus.n5 plus.n4 26.2914
R29 plus.n24 plus.n23 26.2914
R30 plus.n19 plus.n18 26.2914
R31 plus.n9 plus.n2 21.9096
R32 plus.n5 plus.n2 21.9096
R33 plus.n23 plus.n16 21.9096
R34 plus.n19 plus.n16 21.9096
R35 plus.n4 plus.n3 19.0667
R36 plus.n18 plus.n17 19.0667
R37 plus.n11 plus.n10 17.5278
R38 plus.n25 plus.n24 17.5278
R39 plus plus.n13 11.1463
R40 plus.n7 plus.n6 0.189894
R41 plus.n8 plus.n7 0.189894
R42 plus.n8 plus.n1 0.189894
R43 plus.n1 plus.n0 0.189894
R44 plus.n13 plus.n0 0.189894
R45 plus.n27 plus.n14 0.189894
R46 plus.n15 plus.n14 0.189894
R47 plus.n22 plus.n15 0.189894
R48 plus.n22 plus.n21 0.189894
R49 plus.n21 plus.n20 0.189894
R50 source.n5 source.t19 51.0588
R51 source.n19 source.t2 51.0586
R52 source.n14 source.t10 51.0586
R53 source.n0 source.t15 51.0586
R54 source.n2 source.n1 48.8588
R55 source.n4 source.n3 48.8588
R56 source.n7 source.n6 48.8588
R57 source.n9 source.n8 48.8588
R58 source.n18 source.n17 48.8586
R59 source.n16 source.n15 48.8586
R60 source.n13 source.n12 48.8586
R61 source.n11 source.n10 48.8586
R62 source.n11 source.n9 20.7909
R63 source.n20 source.n0 14.196
R64 source.n20 source.n19 5.7074
R65 source.n17 source.t5 2.2005
R66 source.n17 source.t4 2.2005
R67 source.n15 source.t7 2.2005
R68 source.n15 source.t3 2.2005
R69 source.n12 source.t16 2.2005
R70 source.n12 source.t18 2.2005
R71 source.n10 source.t9 2.2005
R72 source.n10 source.t14 2.2005
R73 source.n1 source.t13 2.2005
R74 source.n1 source.t17 2.2005
R75 source.n3 source.t12 2.2005
R76 source.n3 source.t11 2.2005
R77 source.n6 source.t0 2.2005
R78 source.n6 source.t1 2.2005
R79 source.n8 source.t6 2.2005
R80 source.n8 source.t8 2.2005
R81 source.n5 source.n4 0.914293
R82 source.n16 source.n14 0.914293
R83 source.n9 source.n7 0.888431
R84 source.n7 source.n5 0.888431
R85 source.n4 source.n2 0.888431
R86 source.n2 source.n0 0.888431
R87 source.n13 source.n11 0.888431
R88 source.n14 source.n13 0.888431
R89 source.n18 source.n16 0.888431
R90 source.n19 source.n18 0.888431
R91 source source.n20 0.188
R92 drain_left.n5 drain_left.t7 68.6255
R93 drain_left.n1 drain_left.t5 68.6253
R94 drain_left.n3 drain_left.n2 66.1479
R95 drain_left.n5 drain_left.n4 65.5376
R96 drain_left.n7 drain_left.n6 65.5374
R97 drain_left.n1 drain_left.n0 65.5373
R98 drain_left drain_left.n3 28.8681
R99 drain_left drain_left.n7 6.54115
R100 drain_left.n2 drain_left.t0 2.2005
R101 drain_left.n2 drain_left.t1 2.2005
R102 drain_left.n0 drain_left.t6 2.2005
R103 drain_left.n0 drain_left.t4 2.2005
R104 drain_left.n6 drain_left.t3 2.2005
R105 drain_left.n6 drain_left.t8 2.2005
R106 drain_left.n4 drain_left.t2 2.2005
R107 drain_left.n4 drain_left.t9 2.2005
R108 drain_left.n7 drain_left.n5 0.888431
R109 drain_left.n3 drain_left.n1 0.167137
R110 minus.n3 minus.t3 388.724
R111 minus.n17 minus.t9 388.724
R112 minus.n4 minus.t0 365.976
R113 minus.n6 minus.t2 365.976
R114 minus.n10 minus.t7 365.976
R115 minus.n12 minus.t1 365.976
R116 minus.n18 minus.t8 365.976
R117 minus.n20 minus.t4 365.976
R118 minus.n24 minus.t5 365.976
R119 minus.n26 minus.t6 365.976
R120 minus.n13 minus.n12 161.3
R121 minus.n11 minus.n0 161.3
R122 minus.n10 minus.n9 161.3
R123 minus.n8 minus.n1 161.3
R124 minus.n7 minus.n6 161.3
R125 minus.n5 minus.n2 161.3
R126 minus.n27 minus.n26 161.3
R127 minus.n25 minus.n14 161.3
R128 minus.n24 minus.n23 161.3
R129 minus.n22 minus.n15 161.3
R130 minus.n21 minus.n20 161.3
R131 minus.n19 minus.n16 161.3
R132 minus.n3 minus.n2 44.8741
R133 minus.n17 minus.n16 44.8741
R134 minus.n28 minus.n13 34.3812
R135 minus.n12 minus.n11 30.6732
R136 minus.n26 minus.n25 30.6732
R137 minus.n5 minus.n4 26.2914
R138 minus.n10 minus.n1 26.2914
R139 minus.n19 minus.n18 26.2914
R140 minus.n24 minus.n15 26.2914
R141 minus.n6 minus.n5 21.9096
R142 minus.n6 minus.n1 21.9096
R143 minus.n20 minus.n19 21.9096
R144 minus.n20 minus.n15 21.9096
R145 minus.n4 minus.n3 19.0667
R146 minus.n18 minus.n17 19.0667
R147 minus.n11 minus.n10 17.5278
R148 minus.n25 minus.n24 17.5278
R149 minus.n28 minus.n27 6.63876
R150 minus.n13 minus.n0 0.189894
R151 minus.n9 minus.n0 0.189894
R152 minus.n9 minus.n8 0.189894
R153 minus.n8 minus.n7 0.189894
R154 minus.n7 minus.n2 0.189894
R155 minus.n21 minus.n16 0.189894
R156 minus.n22 minus.n21 0.189894
R157 minus.n23 minus.n22 0.189894
R158 minus.n23 minus.n14 0.189894
R159 minus.n27 minus.n14 0.189894
R160 minus minus.n28 0.188
R161 drain_right.n1 drain_right.t0 68.6253
R162 drain_right.n7 drain_right.t8 67.7376
R163 drain_right.n6 drain_right.n4 66.4254
R164 drain_right.n3 drain_right.n2 66.1479
R165 drain_right.n6 drain_right.n5 65.5376
R166 drain_right.n1 drain_right.n0 65.5373
R167 drain_right drain_right.n3 28.3148
R168 drain_right drain_right.n7 6.09718
R169 drain_right.n2 drain_right.t4 2.2005
R170 drain_right.n2 drain_right.t3 2.2005
R171 drain_right.n0 drain_right.t1 2.2005
R172 drain_right.n0 drain_right.t5 2.2005
R173 drain_right.n4 drain_right.t9 2.2005
R174 drain_right.n4 drain_right.t6 2.2005
R175 drain_right.n5 drain_right.t2 2.2005
R176 drain_right.n5 drain_right.t7 2.2005
R177 drain_right.n7 drain_right.n6 0.888431
R178 drain_right.n3 drain_right.n1 0.167137
C0 source plus 5.10863f
C1 source drain_left 11.4165f
C2 drain_left plus 5.33255f
C3 drain_right minus 5.14403f
C4 source drain_right 11.411901f
C5 drain_right plus 0.34671f
C6 drain_right drain_left 0.968193f
C7 source minus 5.09421f
C8 minus plus 5.02155f
C9 drain_left minus 0.171897f
C10 drain_right a_n1952_n2688# 6.11472f
C11 drain_left a_n1952_n2688# 6.41574f
C12 source a_n1952_n2688# 5.420299f
C13 minus a_n1952_n2688# 7.43419f
C14 plus a_n1952_n2688# 8.96728f
C15 drain_right.t0 a_n1952_n2688# 1.92374f
C16 drain_right.t1 a_n1952_n2688# 0.172398f
C17 drain_right.t5 a_n1952_n2688# 0.172398f
C18 drain_right.n0 a_n1952_n2688# 1.50791f
C19 drain_right.n1 a_n1952_n2688# 0.607545f
C20 drain_right.t4 a_n1952_n2688# 0.172398f
C21 drain_right.t3 a_n1952_n2688# 0.172398f
C22 drain_right.n2 a_n1952_n2688# 1.51088f
C23 drain_right.n3 a_n1952_n2688# 1.34024f
C24 drain_right.t9 a_n1952_n2688# 0.172398f
C25 drain_right.t6 a_n1952_n2688# 0.172398f
C26 drain_right.n4 a_n1952_n2688# 1.51249f
C27 drain_right.t2 a_n1952_n2688# 0.172398f
C28 drain_right.t7 a_n1952_n2688# 0.172398f
C29 drain_right.n5 a_n1952_n2688# 1.50791f
C30 drain_right.n6 a_n1952_n2688# 0.670934f
C31 drain_right.t8 a_n1952_n2688# 1.91945f
C32 drain_right.n7 a_n1952_n2688# 0.55471f
C33 minus.n0 a_n1952_n2688# 0.042867f
C34 minus.n1 a_n1952_n2688# 0.009727f
C35 minus.t7 a_n1952_n2688# 0.77449f
C36 minus.n2 a_n1952_n2688# 0.179044f
C37 minus.t3 a_n1952_n2688# 0.793524f
C38 minus.n3 a_n1952_n2688# 0.310276f
C39 minus.t0 a_n1952_n2688# 0.77449f
C40 minus.n4 a_n1952_n2688# 0.329721f
C41 minus.n5 a_n1952_n2688# 0.009727f
C42 minus.t2 a_n1952_n2688# 0.77449f
C43 minus.n6 a_n1952_n2688# 0.325402f
C44 minus.n7 a_n1952_n2688# 0.042867f
C45 minus.n8 a_n1952_n2688# 0.042867f
C46 minus.n9 a_n1952_n2688# 0.042867f
C47 minus.n10 a_n1952_n2688# 0.325402f
C48 minus.n11 a_n1952_n2688# 0.009727f
C49 minus.t1 a_n1952_n2688# 0.77449f
C50 minus.n12 a_n1952_n2688# 0.323023f
C51 minus.n13 a_n1952_n2688# 1.40157f
C52 minus.n14 a_n1952_n2688# 0.042867f
C53 minus.n15 a_n1952_n2688# 0.009727f
C54 minus.n16 a_n1952_n2688# 0.179044f
C55 minus.t9 a_n1952_n2688# 0.793524f
C56 minus.n17 a_n1952_n2688# 0.310276f
C57 minus.t8 a_n1952_n2688# 0.77449f
C58 minus.n18 a_n1952_n2688# 0.329721f
C59 minus.n19 a_n1952_n2688# 0.009727f
C60 minus.t4 a_n1952_n2688# 0.77449f
C61 minus.n20 a_n1952_n2688# 0.325402f
C62 minus.n21 a_n1952_n2688# 0.042867f
C63 minus.n22 a_n1952_n2688# 0.042867f
C64 minus.n23 a_n1952_n2688# 0.042867f
C65 minus.t5 a_n1952_n2688# 0.77449f
C66 minus.n24 a_n1952_n2688# 0.325402f
C67 minus.n25 a_n1952_n2688# 0.009727f
C68 minus.t6 a_n1952_n2688# 0.77449f
C69 minus.n26 a_n1952_n2688# 0.323023f
C70 minus.n27 a_n1952_n2688# 0.294172f
C71 minus.n28 a_n1952_n2688# 1.70611f
C72 drain_left.t5 a_n1952_n2688# 1.93593f
C73 drain_left.t6 a_n1952_n2688# 0.173491f
C74 drain_left.t4 a_n1952_n2688# 0.173491f
C75 drain_left.n0 a_n1952_n2688# 1.51747f
C76 drain_left.n1 a_n1952_n2688# 0.611396f
C77 drain_left.t0 a_n1952_n2688# 0.173491f
C78 drain_left.t1 a_n1952_n2688# 0.173491f
C79 drain_left.n2 a_n1952_n2688# 1.52046f
C80 drain_left.n3 a_n1952_n2688# 1.39887f
C81 drain_left.t7 a_n1952_n2688# 1.93593f
C82 drain_left.t2 a_n1952_n2688# 0.173491f
C83 drain_left.t9 a_n1952_n2688# 0.173491f
C84 drain_left.n4 a_n1952_n2688# 1.51747f
C85 drain_left.n5 a_n1952_n2688# 0.664692f
C86 drain_left.t3 a_n1952_n2688# 0.173491f
C87 drain_left.t8 a_n1952_n2688# 0.173491f
C88 drain_left.n6 a_n1952_n2688# 1.51746f
C89 drain_left.n7 a_n1952_n2688# 0.550754f
C90 source.t15 a_n1952_n2688# 1.98047f
C91 source.n0 a_n1952_n2688# 1.18734f
C92 source.t13 a_n1952_n2688# 0.185725f
C93 source.t17 a_n1952_n2688# 0.185725f
C94 source.n1 a_n1952_n2688# 1.55477f
C95 source.n2 a_n1952_n2688# 0.392818f
C96 source.t12 a_n1952_n2688# 0.185725f
C97 source.t11 a_n1952_n2688# 0.185725f
C98 source.n3 a_n1952_n2688# 1.55477f
C99 source.n4 a_n1952_n2688# 0.394994f
C100 source.t19 a_n1952_n2688# 1.98048f
C101 source.n5 a_n1952_n2688# 0.475808f
C102 source.t0 a_n1952_n2688# 0.185725f
C103 source.t1 a_n1952_n2688# 0.185725f
C104 source.n6 a_n1952_n2688# 1.55477f
C105 source.n7 a_n1952_n2688# 0.392818f
C106 source.t6 a_n1952_n2688# 0.185725f
C107 source.t8 a_n1952_n2688# 0.185725f
C108 source.n8 a_n1952_n2688# 1.55477f
C109 source.n9 a_n1952_n2688# 1.57019f
C110 source.t9 a_n1952_n2688# 0.185725f
C111 source.t14 a_n1952_n2688# 0.185725f
C112 source.n10 a_n1952_n2688# 1.55476f
C113 source.n11 a_n1952_n2688# 1.57019f
C114 source.t16 a_n1952_n2688# 0.185725f
C115 source.t18 a_n1952_n2688# 0.185725f
C116 source.n12 a_n1952_n2688# 1.55476f
C117 source.n13 a_n1952_n2688# 0.392822f
C118 source.t10 a_n1952_n2688# 1.98047f
C119 source.n14 a_n1952_n2688# 0.475813f
C120 source.t7 a_n1952_n2688# 0.185725f
C121 source.t3 a_n1952_n2688# 0.185725f
C122 source.n15 a_n1952_n2688# 1.55476f
C123 source.n16 a_n1952_n2688# 0.394998f
C124 source.t5 a_n1952_n2688# 0.185725f
C125 source.t4 a_n1952_n2688# 0.185725f
C126 source.n17 a_n1952_n2688# 1.55476f
C127 source.n18 a_n1952_n2688# 0.392822f
C128 source.t2 a_n1952_n2688# 1.98047f
C129 source.n19 a_n1952_n2688# 0.608798f
C130 source.n20 a_n1952_n2688# 1.37502f
C131 plus.n0 a_n1952_n2688# 0.04368f
C132 plus.t1 a_n1952_n2688# 0.789182f
C133 plus.t6 a_n1952_n2688# 0.789182f
C134 plus.n1 a_n1952_n2688# 0.04368f
C135 plus.t0 a_n1952_n2688# 0.789182f
C136 plus.n2 a_n1952_n2688# 0.331574f
C137 plus.t2 a_n1952_n2688# 0.808576f
C138 plus.n3 a_n1952_n2688# 0.316162f
C139 plus.t7 a_n1952_n2688# 0.789182f
C140 plus.n4 a_n1952_n2688# 0.335975f
C141 plus.n5 a_n1952_n2688# 0.009912f
C142 plus.n6 a_n1952_n2688# 0.182441f
C143 plus.n7 a_n1952_n2688# 0.04368f
C144 plus.n8 a_n1952_n2688# 0.04368f
C145 plus.n9 a_n1952_n2688# 0.009912f
C146 plus.n10 a_n1952_n2688# 0.331574f
C147 plus.n11 a_n1952_n2688# 0.009912f
C148 plus.n12 a_n1952_n2688# 0.329151f
C149 plus.n13 a_n1952_n2688# 0.443706f
C150 plus.n14 a_n1952_n2688# 0.04368f
C151 plus.t4 a_n1952_n2688# 0.789182f
C152 plus.n15 a_n1952_n2688# 0.04368f
C153 plus.t3 a_n1952_n2688# 0.789182f
C154 plus.t5 a_n1952_n2688# 0.789182f
C155 plus.n16 a_n1952_n2688# 0.331574f
C156 plus.t8 a_n1952_n2688# 0.808576f
C157 plus.n17 a_n1952_n2688# 0.316162f
C158 plus.t9 a_n1952_n2688# 0.789182f
C159 plus.n18 a_n1952_n2688# 0.335975f
C160 plus.n19 a_n1952_n2688# 0.009912f
C161 plus.n20 a_n1952_n2688# 0.182441f
C162 plus.n21 a_n1952_n2688# 0.04368f
C163 plus.n22 a_n1952_n2688# 0.04368f
C164 plus.n23 a_n1952_n2688# 0.009912f
C165 plus.n24 a_n1952_n2688# 0.331574f
C166 plus.n25 a_n1952_n2688# 0.009912f
C167 plus.n26 a_n1952_n2688# 0.329151f
C168 plus.n27 a_n1952_n2688# 1.24784f
.ends

