* NGSPICE file created from diffpair697.ext - technology: sky130A

.subckt diffpair697 minus drain_right drain_left source plus
X0 source.t31 plus.t0 drain_left.t11 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X1 source.t30 plus.t1 drain_left.t10 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.6
X2 drain_left.t5 plus.t2 source.t29 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.6
X3 source.t28 plus.t3 drain_left.t4 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X4 drain_right.t15 minus.t0 source.t9 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X5 drain_left.t15 plus.t4 source.t27 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X6 source.t6 minus.t1 drain_right.t14 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.6
X7 source.t14 minus.t2 drain_right.t13 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X8 drain_right.t12 minus.t3 source.t15 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X9 drain_left.t14 plus.t5 source.t26 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X10 drain_right.t11 minus.t4 source.t3 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X11 drain_right.t10 minus.t5 source.t10 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X12 source.t4 minus.t6 drain_right.t9 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X13 source.t25 plus.t6 drain_left.t13 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X14 a_n2390_n5888# a_n2390_n5888# a_n2390_n5888# a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.6
X15 a_n2390_n5888# a_n2390_n5888# a_n2390_n5888# a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.6
X16 source.t24 plus.t7 drain_left.t12 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X17 source.t8 minus.t7 drain_right.t8 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X18 source.t11 minus.t8 drain_right.t7 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X19 source.t23 plus.t8 drain_left.t1 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X20 drain_right.t6 minus.t9 source.t0 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X21 a_n2390_n5888# a_n2390_n5888# a_n2390_n5888# a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.6
X22 drain_left.t0 plus.t9 source.t22 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X23 source.t12 minus.t10 drain_right.t5 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X24 source.t21 plus.t10 drain_left.t3 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X25 drain_right.t4 minus.t11 source.t1 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.6
X26 source.t7 minus.t12 drain_right.t3 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X27 drain_left.t2 plus.t11 source.t20 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X28 source.t19 plus.t12 drain_left.t9 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.6
X29 a_n2390_n5888# a_n2390_n5888# a_n2390_n5888# a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.6
X30 source.t2 minus.t13 drain_right.t2 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.6
X31 drain_left.t8 plus.t13 source.t18 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X32 drain_left.t7 plus.t14 source.t17 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X33 drain_right.t1 minus.t14 source.t13 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.6
X34 drain_right.t0 minus.t15 source.t5 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X35 drain_left.t6 plus.t15 source.t16 a_n2390_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.6
R0 plus.n6 plus.t12 1090.62
R1 plus.n30 plus.t15 1090.62
R2 plus.n22 plus.t2 1069.64
R3 plus.n21 plus.t3 1069.64
R4 plus.n1 plus.t4 1069.64
R5 plus.n15 plus.t7 1069.64
R6 plus.n3 plus.t9 1069.64
R7 plus.n9 plus.t10 1069.64
R8 plus.n5 plus.t11 1069.64
R9 plus.n46 plus.t1 1069.64
R10 plus.n45 plus.t14 1069.64
R11 plus.n25 plus.t6 1069.64
R12 plus.n39 plus.t5 1069.64
R13 plus.n27 plus.t0 1069.64
R14 plus.n33 plus.t13 1069.64
R15 plus.n29 plus.t8 1069.64
R16 plus.n8 plus.n7 161.3
R17 plus.n9 plus.n4 161.3
R18 plus.n11 plus.n10 161.3
R19 plus.n12 plus.n3 161.3
R20 plus.n14 plus.n13 161.3
R21 plus.n15 plus.n2 161.3
R22 plus.n17 plus.n16 161.3
R23 plus.n18 plus.n1 161.3
R24 plus.n20 plus.n19 161.3
R25 plus.n21 plus.n0 161.3
R26 plus.n23 plus.n22 161.3
R27 plus.n32 plus.n31 161.3
R28 plus.n33 plus.n28 161.3
R29 plus.n35 plus.n34 161.3
R30 plus.n36 plus.n27 161.3
R31 plus.n38 plus.n37 161.3
R32 plus.n39 plus.n26 161.3
R33 plus.n41 plus.n40 161.3
R34 plus.n42 plus.n25 161.3
R35 plus.n44 plus.n43 161.3
R36 plus.n45 plus.n24 161.3
R37 plus.n47 plus.n46 161.3
R38 plus.n7 plus.n6 70.4033
R39 plus.n31 plus.n30 70.4033
R40 plus.n22 plus.n21 48.2005
R41 plus.n46 plus.n45 48.2005
R42 plus.n20 plus.n1 44.549
R43 plus.n9 plus.n8 44.549
R44 plus.n44 plus.n25 44.549
R45 plus.n33 plus.n32 44.549
R46 plus plus.n47 37.1354
R47 plus.n16 plus.n15 34.3247
R48 plus.n10 plus.n3 34.3247
R49 plus.n40 plus.n39 34.3247
R50 plus.n34 plus.n27 34.3247
R51 plus.n14 plus.n3 24.1005
R52 plus.n15 plus.n14 24.1005
R53 plus.n39 plus.n38 24.1005
R54 plus.n38 plus.n27 24.1005
R55 plus.n6 plus.n5 20.9576
R56 plus.n30 plus.n29 20.9576
R57 plus plus.n23 17.224
R58 plus.n16 plus.n1 13.8763
R59 plus.n10 plus.n9 13.8763
R60 plus.n40 plus.n25 13.8763
R61 plus.n34 plus.n33 13.8763
R62 plus.n21 plus.n20 3.65202
R63 plus.n8 plus.n5 3.65202
R64 plus.n45 plus.n44 3.65202
R65 plus.n32 plus.n29 3.65202
R66 plus.n7 plus.n4 0.189894
R67 plus.n11 plus.n4 0.189894
R68 plus.n12 plus.n11 0.189894
R69 plus.n13 plus.n12 0.189894
R70 plus.n13 plus.n2 0.189894
R71 plus.n17 plus.n2 0.189894
R72 plus.n18 plus.n17 0.189894
R73 plus.n19 plus.n18 0.189894
R74 plus.n19 plus.n0 0.189894
R75 plus.n23 plus.n0 0.189894
R76 plus.n47 plus.n24 0.189894
R77 plus.n43 plus.n24 0.189894
R78 plus.n43 plus.n42 0.189894
R79 plus.n42 plus.n41 0.189894
R80 plus.n41 plus.n26 0.189894
R81 plus.n37 plus.n26 0.189894
R82 plus.n37 plus.n36 0.189894
R83 plus.n36 plus.n35 0.189894
R84 plus.n35 plus.n28 0.189894
R85 plus.n31 plus.n28 0.189894
R86 drain_left.n5 drain_left.n3 59.5172
R87 drain_left.n2 drain_left.n0 59.5172
R88 drain_left.n9 drain_left.n7 59.5172
R89 drain_left.n5 drain_left.n4 58.7154
R90 drain_left.n2 drain_left.n1 58.7154
R91 drain_left.n11 drain_left.n10 58.7154
R92 drain_left.n9 drain_left.n8 58.7154
R93 drain_left.n13 drain_left.n12 58.7153
R94 drain_left drain_left.n6 42.4268
R95 drain_left drain_left.n13 6.45494
R96 drain_left.n11 drain_left.n9 0.802224
R97 drain_left.n13 drain_left.n11 0.802224
R98 drain_left.n3 drain_left.t1 0.7925
R99 drain_left.n3 drain_left.t6 0.7925
R100 drain_left.n4 drain_left.t11 0.7925
R101 drain_left.n4 drain_left.t8 0.7925
R102 drain_left.n1 drain_left.t13 0.7925
R103 drain_left.n1 drain_left.t14 0.7925
R104 drain_left.n0 drain_left.t10 0.7925
R105 drain_left.n0 drain_left.t7 0.7925
R106 drain_left.n12 drain_left.t4 0.7925
R107 drain_left.n12 drain_left.t5 0.7925
R108 drain_left.n10 drain_left.t12 0.7925
R109 drain_left.n10 drain_left.t15 0.7925
R110 drain_left.n8 drain_left.t3 0.7925
R111 drain_left.n8 drain_left.t0 0.7925
R112 drain_left.n7 drain_left.t9 0.7925
R113 drain_left.n7 drain_left.t2 0.7925
R114 drain_left.n6 drain_left.n5 0.346016
R115 drain_left.n6 drain_left.n2 0.346016
R116 source.n1138 source.n1004 289.615
R117 source.n992 source.n858 289.615
R118 source.n852 source.n718 289.615
R119 source.n706 source.n572 289.615
R120 source.n134 source.n0 289.615
R121 source.n280 source.n146 289.615
R122 source.n420 source.n286 289.615
R123 source.n566 source.n432 289.615
R124 source.n1048 source.n1047 185
R125 source.n1053 source.n1052 185
R126 source.n1055 source.n1054 185
R127 source.n1044 source.n1043 185
R128 source.n1061 source.n1060 185
R129 source.n1063 source.n1062 185
R130 source.n1040 source.n1039 185
R131 source.n1070 source.n1069 185
R132 source.n1071 source.n1038 185
R133 source.n1073 source.n1072 185
R134 source.n1036 source.n1035 185
R135 source.n1079 source.n1078 185
R136 source.n1081 source.n1080 185
R137 source.n1032 source.n1031 185
R138 source.n1087 source.n1086 185
R139 source.n1089 source.n1088 185
R140 source.n1028 source.n1027 185
R141 source.n1095 source.n1094 185
R142 source.n1097 source.n1096 185
R143 source.n1024 source.n1023 185
R144 source.n1103 source.n1102 185
R145 source.n1105 source.n1104 185
R146 source.n1020 source.n1019 185
R147 source.n1111 source.n1110 185
R148 source.n1114 source.n1113 185
R149 source.n1112 source.n1016 185
R150 source.n1119 source.n1015 185
R151 source.n1121 source.n1120 185
R152 source.n1123 source.n1122 185
R153 source.n1012 source.n1011 185
R154 source.n1129 source.n1128 185
R155 source.n1131 source.n1130 185
R156 source.n1008 source.n1007 185
R157 source.n1137 source.n1136 185
R158 source.n1139 source.n1138 185
R159 source.n902 source.n901 185
R160 source.n907 source.n906 185
R161 source.n909 source.n908 185
R162 source.n898 source.n897 185
R163 source.n915 source.n914 185
R164 source.n917 source.n916 185
R165 source.n894 source.n893 185
R166 source.n924 source.n923 185
R167 source.n925 source.n892 185
R168 source.n927 source.n926 185
R169 source.n890 source.n889 185
R170 source.n933 source.n932 185
R171 source.n935 source.n934 185
R172 source.n886 source.n885 185
R173 source.n941 source.n940 185
R174 source.n943 source.n942 185
R175 source.n882 source.n881 185
R176 source.n949 source.n948 185
R177 source.n951 source.n950 185
R178 source.n878 source.n877 185
R179 source.n957 source.n956 185
R180 source.n959 source.n958 185
R181 source.n874 source.n873 185
R182 source.n965 source.n964 185
R183 source.n968 source.n967 185
R184 source.n966 source.n870 185
R185 source.n973 source.n869 185
R186 source.n975 source.n974 185
R187 source.n977 source.n976 185
R188 source.n866 source.n865 185
R189 source.n983 source.n982 185
R190 source.n985 source.n984 185
R191 source.n862 source.n861 185
R192 source.n991 source.n990 185
R193 source.n993 source.n992 185
R194 source.n762 source.n761 185
R195 source.n767 source.n766 185
R196 source.n769 source.n768 185
R197 source.n758 source.n757 185
R198 source.n775 source.n774 185
R199 source.n777 source.n776 185
R200 source.n754 source.n753 185
R201 source.n784 source.n783 185
R202 source.n785 source.n752 185
R203 source.n787 source.n786 185
R204 source.n750 source.n749 185
R205 source.n793 source.n792 185
R206 source.n795 source.n794 185
R207 source.n746 source.n745 185
R208 source.n801 source.n800 185
R209 source.n803 source.n802 185
R210 source.n742 source.n741 185
R211 source.n809 source.n808 185
R212 source.n811 source.n810 185
R213 source.n738 source.n737 185
R214 source.n817 source.n816 185
R215 source.n819 source.n818 185
R216 source.n734 source.n733 185
R217 source.n825 source.n824 185
R218 source.n828 source.n827 185
R219 source.n826 source.n730 185
R220 source.n833 source.n729 185
R221 source.n835 source.n834 185
R222 source.n837 source.n836 185
R223 source.n726 source.n725 185
R224 source.n843 source.n842 185
R225 source.n845 source.n844 185
R226 source.n722 source.n721 185
R227 source.n851 source.n850 185
R228 source.n853 source.n852 185
R229 source.n616 source.n615 185
R230 source.n621 source.n620 185
R231 source.n623 source.n622 185
R232 source.n612 source.n611 185
R233 source.n629 source.n628 185
R234 source.n631 source.n630 185
R235 source.n608 source.n607 185
R236 source.n638 source.n637 185
R237 source.n639 source.n606 185
R238 source.n641 source.n640 185
R239 source.n604 source.n603 185
R240 source.n647 source.n646 185
R241 source.n649 source.n648 185
R242 source.n600 source.n599 185
R243 source.n655 source.n654 185
R244 source.n657 source.n656 185
R245 source.n596 source.n595 185
R246 source.n663 source.n662 185
R247 source.n665 source.n664 185
R248 source.n592 source.n591 185
R249 source.n671 source.n670 185
R250 source.n673 source.n672 185
R251 source.n588 source.n587 185
R252 source.n679 source.n678 185
R253 source.n682 source.n681 185
R254 source.n680 source.n584 185
R255 source.n687 source.n583 185
R256 source.n689 source.n688 185
R257 source.n691 source.n690 185
R258 source.n580 source.n579 185
R259 source.n697 source.n696 185
R260 source.n699 source.n698 185
R261 source.n576 source.n575 185
R262 source.n705 source.n704 185
R263 source.n707 source.n706 185
R264 source.n135 source.n134 185
R265 source.n133 source.n132 185
R266 source.n4 source.n3 185
R267 source.n127 source.n126 185
R268 source.n125 source.n124 185
R269 source.n8 source.n7 185
R270 source.n119 source.n118 185
R271 source.n117 source.n116 185
R272 source.n115 source.n11 185
R273 source.n15 source.n12 185
R274 source.n110 source.n109 185
R275 source.n108 source.n107 185
R276 source.n17 source.n16 185
R277 source.n102 source.n101 185
R278 source.n100 source.n99 185
R279 source.n21 source.n20 185
R280 source.n94 source.n93 185
R281 source.n92 source.n91 185
R282 source.n25 source.n24 185
R283 source.n86 source.n85 185
R284 source.n84 source.n83 185
R285 source.n29 source.n28 185
R286 source.n78 source.n77 185
R287 source.n76 source.n75 185
R288 source.n33 source.n32 185
R289 source.n70 source.n69 185
R290 source.n68 source.n35 185
R291 source.n67 source.n66 185
R292 source.n38 source.n36 185
R293 source.n61 source.n60 185
R294 source.n59 source.n58 185
R295 source.n42 source.n41 185
R296 source.n53 source.n52 185
R297 source.n51 source.n50 185
R298 source.n46 source.n45 185
R299 source.n281 source.n280 185
R300 source.n279 source.n278 185
R301 source.n150 source.n149 185
R302 source.n273 source.n272 185
R303 source.n271 source.n270 185
R304 source.n154 source.n153 185
R305 source.n265 source.n264 185
R306 source.n263 source.n262 185
R307 source.n261 source.n157 185
R308 source.n161 source.n158 185
R309 source.n256 source.n255 185
R310 source.n254 source.n253 185
R311 source.n163 source.n162 185
R312 source.n248 source.n247 185
R313 source.n246 source.n245 185
R314 source.n167 source.n166 185
R315 source.n240 source.n239 185
R316 source.n238 source.n237 185
R317 source.n171 source.n170 185
R318 source.n232 source.n231 185
R319 source.n230 source.n229 185
R320 source.n175 source.n174 185
R321 source.n224 source.n223 185
R322 source.n222 source.n221 185
R323 source.n179 source.n178 185
R324 source.n216 source.n215 185
R325 source.n214 source.n181 185
R326 source.n213 source.n212 185
R327 source.n184 source.n182 185
R328 source.n207 source.n206 185
R329 source.n205 source.n204 185
R330 source.n188 source.n187 185
R331 source.n199 source.n198 185
R332 source.n197 source.n196 185
R333 source.n192 source.n191 185
R334 source.n421 source.n420 185
R335 source.n419 source.n418 185
R336 source.n290 source.n289 185
R337 source.n413 source.n412 185
R338 source.n411 source.n410 185
R339 source.n294 source.n293 185
R340 source.n405 source.n404 185
R341 source.n403 source.n402 185
R342 source.n401 source.n297 185
R343 source.n301 source.n298 185
R344 source.n396 source.n395 185
R345 source.n394 source.n393 185
R346 source.n303 source.n302 185
R347 source.n388 source.n387 185
R348 source.n386 source.n385 185
R349 source.n307 source.n306 185
R350 source.n380 source.n379 185
R351 source.n378 source.n377 185
R352 source.n311 source.n310 185
R353 source.n372 source.n371 185
R354 source.n370 source.n369 185
R355 source.n315 source.n314 185
R356 source.n364 source.n363 185
R357 source.n362 source.n361 185
R358 source.n319 source.n318 185
R359 source.n356 source.n355 185
R360 source.n354 source.n321 185
R361 source.n353 source.n352 185
R362 source.n324 source.n322 185
R363 source.n347 source.n346 185
R364 source.n345 source.n344 185
R365 source.n328 source.n327 185
R366 source.n339 source.n338 185
R367 source.n337 source.n336 185
R368 source.n332 source.n331 185
R369 source.n567 source.n566 185
R370 source.n565 source.n564 185
R371 source.n436 source.n435 185
R372 source.n559 source.n558 185
R373 source.n557 source.n556 185
R374 source.n440 source.n439 185
R375 source.n551 source.n550 185
R376 source.n549 source.n548 185
R377 source.n547 source.n443 185
R378 source.n447 source.n444 185
R379 source.n542 source.n541 185
R380 source.n540 source.n539 185
R381 source.n449 source.n448 185
R382 source.n534 source.n533 185
R383 source.n532 source.n531 185
R384 source.n453 source.n452 185
R385 source.n526 source.n525 185
R386 source.n524 source.n523 185
R387 source.n457 source.n456 185
R388 source.n518 source.n517 185
R389 source.n516 source.n515 185
R390 source.n461 source.n460 185
R391 source.n510 source.n509 185
R392 source.n508 source.n507 185
R393 source.n465 source.n464 185
R394 source.n502 source.n501 185
R395 source.n500 source.n467 185
R396 source.n499 source.n498 185
R397 source.n470 source.n468 185
R398 source.n493 source.n492 185
R399 source.n491 source.n490 185
R400 source.n474 source.n473 185
R401 source.n485 source.n484 185
R402 source.n483 source.n482 185
R403 source.n478 source.n477 185
R404 source.n1049 source.t13 149.524
R405 source.n903 source.t2 149.524
R406 source.n763 source.t16 149.524
R407 source.n617 source.t30 149.524
R408 source.n47 source.t29 149.524
R409 source.n193 source.t19 149.524
R410 source.n333 source.t1 149.524
R411 source.n479 source.t6 149.524
R412 source.n1053 source.n1047 104.615
R413 source.n1054 source.n1053 104.615
R414 source.n1054 source.n1043 104.615
R415 source.n1061 source.n1043 104.615
R416 source.n1062 source.n1061 104.615
R417 source.n1062 source.n1039 104.615
R418 source.n1070 source.n1039 104.615
R419 source.n1071 source.n1070 104.615
R420 source.n1072 source.n1071 104.615
R421 source.n1072 source.n1035 104.615
R422 source.n1079 source.n1035 104.615
R423 source.n1080 source.n1079 104.615
R424 source.n1080 source.n1031 104.615
R425 source.n1087 source.n1031 104.615
R426 source.n1088 source.n1087 104.615
R427 source.n1088 source.n1027 104.615
R428 source.n1095 source.n1027 104.615
R429 source.n1096 source.n1095 104.615
R430 source.n1096 source.n1023 104.615
R431 source.n1103 source.n1023 104.615
R432 source.n1104 source.n1103 104.615
R433 source.n1104 source.n1019 104.615
R434 source.n1111 source.n1019 104.615
R435 source.n1113 source.n1111 104.615
R436 source.n1113 source.n1112 104.615
R437 source.n1112 source.n1015 104.615
R438 source.n1121 source.n1015 104.615
R439 source.n1122 source.n1121 104.615
R440 source.n1122 source.n1011 104.615
R441 source.n1129 source.n1011 104.615
R442 source.n1130 source.n1129 104.615
R443 source.n1130 source.n1007 104.615
R444 source.n1137 source.n1007 104.615
R445 source.n1138 source.n1137 104.615
R446 source.n907 source.n901 104.615
R447 source.n908 source.n907 104.615
R448 source.n908 source.n897 104.615
R449 source.n915 source.n897 104.615
R450 source.n916 source.n915 104.615
R451 source.n916 source.n893 104.615
R452 source.n924 source.n893 104.615
R453 source.n925 source.n924 104.615
R454 source.n926 source.n925 104.615
R455 source.n926 source.n889 104.615
R456 source.n933 source.n889 104.615
R457 source.n934 source.n933 104.615
R458 source.n934 source.n885 104.615
R459 source.n941 source.n885 104.615
R460 source.n942 source.n941 104.615
R461 source.n942 source.n881 104.615
R462 source.n949 source.n881 104.615
R463 source.n950 source.n949 104.615
R464 source.n950 source.n877 104.615
R465 source.n957 source.n877 104.615
R466 source.n958 source.n957 104.615
R467 source.n958 source.n873 104.615
R468 source.n965 source.n873 104.615
R469 source.n967 source.n965 104.615
R470 source.n967 source.n966 104.615
R471 source.n966 source.n869 104.615
R472 source.n975 source.n869 104.615
R473 source.n976 source.n975 104.615
R474 source.n976 source.n865 104.615
R475 source.n983 source.n865 104.615
R476 source.n984 source.n983 104.615
R477 source.n984 source.n861 104.615
R478 source.n991 source.n861 104.615
R479 source.n992 source.n991 104.615
R480 source.n767 source.n761 104.615
R481 source.n768 source.n767 104.615
R482 source.n768 source.n757 104.615
R483 source.n775 source.n757 104.615
R484 source.n776 source.n775 104.615
R485 source.n776 source.n753 104.615
R486 source.n784 source.n753 104.615
R487 source.n785 source.n784 104.615
R488 source.n786 source.n785 104.615
R489 source.n786 source.n749 104.615
R490 source.n793 source.n749 104.615
R491 source.n794 source.n793 104.615
R492 source.n794 source.n745 104.615
R493 source.n801 source.n745 104.615
R494 source.n802 source.n801 104.615
R495 source.n802 source.n741 104.615
R496 source.n809 source.n741 104.615
R497 source.n810 source.n809 104.615
R498 source.n810 source.n737 104.615
R499 source.n817 source.n737 104.615
R500 source.n818 source.n817 104.615
R501 source.n818 source.n733 104.615
R502 source.n825 source.n733 104.615
R503 source.n827 source.n825 104.615
R504 source.n827 source.n826 104.615
R505 source.n826 source.n729 104.615
R506 source.n835 source.n729 104.615
R507 source.n836 source.n835 104.615
R508 source.n836 source.n725 104.615
R509 source.n843 source.n725 104.615
R510 source.n844 source.n843 104.615
R511 source.n844 source.n721 104.615
R512 source.n851 source.n721 104.615
R513 source.n852 source.n851 104.615
R514 source.n621 source.n615 104.615
R515 source.n622 source.n621 104.615
R516 source.n622 source.n611 104.615
R517 source.n629 source.n611 104.615
R518 source.n630 source.n629 104.615
R519 source.n630 source.n607 104.615
R520 source.n638 source.n607 104.615
R521 source.n639 source.n638 104.615
R522 source.n640 source.n639 104.615
R523 source.n640 source.n603 104.615
R524 source.n647 source.n603 104.615
R525 source.n648 source.n647 104.615
R526 source.n648 source.n599 104.615
R527 source.n655 source.n599 104.615
R528 source.n656 source.n655 104.615
R529 source.n656 source.n595 104.615
R530 source.n663 source.n595 104.615
R531 source.n664 source.n663 104.615
R532 source.n664 source.n591 104.615
R533 source.n671 source.n591 104.615
R534 source.n672 source.n671 104.615
R535 source.n672 source.n587 104.615
R536 source.n679 source.n587 104.615
R537 source.n681 source.n679 104.615
R538 source.n681 source.n680 104.615
R539 source.n680 source.n583 104.615
R540 source.n689 source.n583 104.615
R541 source.n690 source.n689 104.615
R542 source.n690 source.n579 104.615
R543 source.n697 source.n579 104.615
R544 source.n698 source.n697 104.615
R545 source.n698 source.n575 104.615
R546 source.n705 source.n575 104.615
R547 source.n706 source.n705 104.615
R548 source.n134 source.n133 104.615
R549 source.n133 source.n3 104.615
R550 source.n126 source.n3 104.615
R551 source.n126 source.n125 104.615
R552 source.n125 source.n7 104.615
R553 source.n118 source.n7 104.615
R554 source.n118 source.n117 104.615
R555 source.n117 source.n11 104.615
R556 source.n15 source.n11 104.615
R557 source.n109 source.n15 104.615
R558 source.n109 source.n108 104.615
R559 source.n108 source.n16 104.615
R560 source.n101 source.n16 104.615
R561 source.n101 source.n100 104.615
R562 source.n100 source.n20 104.615
R563 source.n93 source.n20 104.615
R564 source.n93 source.n92 104.615
R565 source.n92 source.n24 104.615
R566 source.n85 source.n24 104.615
R567 source.n85 source.n84 104.615
R568 source.n84 source.n28 104.615
R569 source.n77 source.n28 104.615
R570 source.n77 source.n76 104.615
R571 source.n76 source.n32 104.615
R572 source.n69 source.n32 104.615
R573 source.n69 source.n68 104.615
R574 source.n68 source.n67 104.615
R575 source.n67 source.n36 104.615
R576 source.n60 source.n36 104.615
R577 source.n60 source.n59 104.615
R578 source.n59 source.n41 104.615
R579 source.n52 source.n41 104.615
R580 source.n52 source.n51 104.615
R581 source.n51 source.n45 104.615
R582 source.n280 source.n279 104.615
R583 source.n279 source.n149 104.615
R584 source.n272 source.n149 104.615
R585 source.n272 source.n271 104.615
R586 source.n271 source.n153 104.615
R587 source.n264 source.n153 104.615
R588 source.n264 source.n263 104.615
R589 source.n263 source.n157 104.615
R590 source.n161 source.n157 104.615
R591 source.n255 source.n161 104.615
R592 source.n255 source.n254 104.615
R593 source.n254 source.n162 104.615
R594 source.n247 source.n162 104.615
R595 source.n247 source.n246 104.615
R596 source.n246 source.n166 104.615
R597 source.n239 source.n166 104.615
R598 source.n239 source.n238 104.615
R599 source.n238 source.n170 104.615
R600 source.n231 source.n170 104.615
R601 source.n231 source.n230 104.615
R602 source.n230 source.n174 104.615
R603 source.n223 source.n174 104.615
R604 source.n223 source.n222 104.615
R605 source.n222 source.n178 104.615
R606 source.n215 source.n178 104.615
R607 source.n215 source.n214 104.615
R608 source.n214 source.n213 104.615
R609 source.n213 source.n182 104.615
R610 source.n206 source.n182 104.615
R611 source.n206 source.n205 104.615
R612 source.n205 source.n187 104.615
R613 source.n198 source.n187 104.615
R614 source.n198 source.n197 104.615
R615 source.n197 source.n191 104.615
R616 source.n420 source.n419 104.615
R617 source.n419 source.n289 104.615
R618 source.n412 source.n289 104.615
R619 source.n412 source.n411 104.615
R620 source.n411 source.n293 104.615
R621 source.n404 source.n293 104.615
R622 source.n404 source.n403 104.615
R623 source.n403 source.n297 104.615
R624 source.n301 source.n297 104.615
R625 source.n395 source.n301 104.615
R626 source.n395 source.n394 104.615
R627 source.n394 source.n302 104.615
R628 source.n387 source.n302 104.615
R629 source.n387 source.n386 104.615
R630 source.n386 source.n306 104.615
R631 source.n379 source.n306 104.615
R632 source.n379 source.n378 104.615
R633 source.n378 source.n310 104.615
R634 source.n371 source.n310 104.615
R635 source.n371 source.n370 104.615
R636 source.n370 source.n314 104.615
R637 source.n363 source.n314 104.615
R638 source.n363 source.n362 104.615
R639 source.n362 source.n318 104.615
R640 source.n355 source.n318 104.615
R641 source.n355 source.n354 104.615
R642 source.n354 source.n353 104.615
R643 source.n353 source.n322 104.615
R644 source.n346 source.n322 104.615
R645 source.n346 source.n345 104.615
R646 source.n345 source.n327 104.615
R647 source.n338 source.n327 104.615
R648 source.n338 source.n337 104.615
R649 source.n337 source.n331 104.615
R650 source.n566 source.n565 104.615
R651 source.n565 source.n435 104.615
R652 source.n558 source.n435 104.615
R653 source.n558 source.n557 104.615
R654 source.n557 source.n439 104.615
R655 source.n550 source.n439 104.615
R656 source.n550 source.n549 104.615
R657 source.n549 source.n443 104.615
R658 source.n447 source.n443 104.615
R659 source.n541 source.n447 104.615
R660 source.n541 source.n540 104.615
R661 source.n540 source.n448 104.615
R662 source.n533 source.n448 104.615
R663 source.n533 source.n532 104.615
R664 source.n532 source.n452 104.615
R665 source.n525 source.n452 104.615
R666 source.n525 source.n524 104.615
R667 source.n524 source.n456 104.615
R668 source.n517 source.n456 104.615
R669 source.n517 source.n516 104.615
R670 source.n516 source.n460 104.615
R671 source.n509 source.n460 104.615
R672 source.n509 source.n508 104.615
R673 source.n508 source.n464 104.615
R674 source.n501 source.n464 104.615
R675 source.n501 source.n500 104.615
R676 source.n500 source.n499 104.615
R677 source.n499 source.n468 104.615
R678 source.n492 source.n468 104.615
R679 source.n492 source.n491 104.615
R680 source.n491 source.n473 104.615
R681 source.n484 source.n473 104.615
R682 source.n484 source.n483 104.615
R683 source.n483 source.n477 104.615
R684 source.t13 source.n1047 52.3082
R685 source.t2 source.n901 52.3082
R686 source.t16 source.n761 52.3082
R687 source.t30 source.n615 52.3082
R688 source.t29 source.n45 52.3082
R689 source.t19 source.n191 52.3082
R690 source.t1 source.n331 52.3082
R691 source.t6 source.n477 52.3082
R692 source.n1003 source.n1002 42.0366
R693 source.n1001 source.n1000 42.0366
R694 source.n999 source.n998 42.0366
R695 source.n717 source.n716 42.0366
R696 source.n715 source.n714 42.0366
R697 source.n713 source.n712 42.0366
R698 source.n141 source.n140 42.0366
R699 source.n143 source.n142 42.0366
R700 source.n145 source.n144 42.0366
R701 source.n427 source.n426 42.0366
R702 source.n429 source.n428 42.0366
R703 source.n431 source.n430 42.0366
R704 source.n711 source.n571 31.9379
R705 source.n1143 source.n1142 30.6338
R706 source.n997 source.n996 30.6338
R707 source.n857 source.n856 30.6338
R708 source.n711 source.n710 30.6338
R709 source.n139 source.n138 30.6338
R710 source.n285 source.n284 30.6338
R711 source.n425 source.n424 30.6338
R712 source.n571 source.n570 30.6338
R713 source.n1144 source.n139 26.2741
R714 source.n1073 source.n1038 13.1884
R715 source.n1120 source.n1119 13.1884
R716 source.n927 source.n892 13.1884
R717 source.n974 source.n973 13.1884
R718 source.n787 source.n752 13.1884
R719 source.n834 source.n833 13.1884
R720 source.n641 source.n606 13.1884
R721 source.n688 source.n687 13.1884
R722 source.n116 source.n115 13.1884
R723 source.n70 source.n35 13.1884
R724 source.n262 source.n261 13.1884
R725 source.n216 source.n181 13.1884
R726 source.n402 source.n401 13.1884
R727 source.n356 source.n321 13.1884
R728 source.n548 source.n547 13.1884
R729 source.n502 source.n467 13.1884
R730 source.n1069 source.n1068 12.8005
R731 source.n1074 source.n1036 12.8005
R732 source.n1118 source.n1016 12.8005
R733 source.n1123 source.n1014 12.8005
R734 source.n923 source.n922 12.8005
R735 source.n928 source.n890 12.8005
R736 source.n972 source.n870 12.8005
R737 source.n977 source.n868 12.8005
R738 source.n783 source.n782 12.8005
R739 source.n788 source.n750 12.8005
R740 source.n832 source.n730 12.8005
R741 source.n837 source.n728 12.8005
R742 source.n637 source.n636 12.8005
R743 source.n642 source.n604 12.8005
R744 source.n686 source.n584 12.8005
R745 source.n691 source.n582 12.8005
R746 source.n119 source.n10 12.8005
R747 source.n114 source.n12 12.8005
R748 source.n71 source.n33 12.8005
R749 source.n66 source.n37 12.8005
R750 source.n265 source.n156 12.8005
R751 source.n260 source.n158 12.8005
R752 source.n217 source.n179 12.8005
R753 source.n212 source.n183 12.8005
R754 source.n405 source.n296 12.8005
R755 source.n400 source.n298 12.8005
R756 source.n357 source.n319 12.8005
R757 source.n352 source.n323 12.8005
R758 source.n551 source.n442 12.8005
R759 source.n546 source.n444 12.8005
R760 source.n503 source.n465 12.8005
R761 source.n498 source.n469 12.8005
R762 source.n1067 source.n1040 12.0247
R763 source.n1078 source.n1077 12.0247
R764 source.n1115 source.n1114 12.0247
R765 source.n1124 source.n1012 12.0247
R766 source.n921 source.n894 12.0247
R767 source.n932 source.n931 12.0247
R768 source.n969 source.n968 12.0247
R769 source.n978 source.n866 12.0247
R770 source.n781 source.n754 12.0247
R771 source.n792 source.n791 12.0247
R772 source.n829 source.n828 12.0247
R773 source.n838 source.n726 12.0247
R774 source.n635 source.n608 12.0247
R775 source.n646 source.n645 12.0247
R776 source.n683 source.n682 12.0247
R777 source.n692 source.n580 12.0247
R778 source.n120 source.n8 12.0247
R779 source.n111 source.n110 12.0247
R780 source.n75 source.n74 12.0247
R781 source.n65 source.n38 12.0247
R782 source.n266 source.n154 12.0247
R783 source.n257 source.n256 12.0247
R784 source.n221 source.n220 12.0247
R785 source.n211 source.n184 12.0247
R786 source.n406 source.n294 12.0247
R787 source.n397 source.n396 12.0247
R788 source.n361 source.n360 12.0247
R789 source.n351 source.n324 12.0247
R790 source.n552 source.n440 12.0247
R791 source.n543 source.n542 12.0247
R792 source.n507 source.n506 12.0247
R793 source.n497 source.n470 12.0247
R794 source.n1064 source.n1063 11.249
R795 source.n1081 source.n1034 11.249
R796 source.n1110 source.n1018 11.249
R797 source.n1128 source.n1127 11.249
R798 source.n918 source.n917 11.249
R799 source.n935 source.n888 11.249
R800 source.n964 source.n872 11.249
R801 source.n982 source.n981 11.249
R802 source.n778 source.n777 11.249
R803 source.n795 source.n748 11.249
R804 source.n824 source.n732 11.249
R805 source.n842 source.n841 11.249
R806 source.n632 source.n631 11.249
R807 source.n649 source.n602 11.249
R808 source.n678 source.n586 11.249
R809 source.n696 source.n695 11.249
R810 source.n124 source.n123 11.249
R811 source.n107 source.n14 11.249
R812 source.n78 source.n31 11.249
R813 source.n62 source.n61 11.249
R814 source.n270 source.n269 11.249
R815 source.n253 source.n160 11.249
R816 source.n224 source.n177 11.249
R817 source.n208 source.n207 11.249
R818 source.n410 source.n409 11.249
R819 source.n393 source.n300 11.249
R820 source.n364 source.n317 11.249
R821 source.n348 source.n347 11.249
R822 source.n556 source.n555 11.249
R823 source.n539 source.n446 11.249
R824 source.n510 source.n463 11.249
R825 source.n494 source.n493 11.249
R826 source.n1060 source.n1042 10.4732
R827 source.n1082 source.n1032 10.4732
R828 source.n1109 source.n1020 10.4732
R829 source.n1131 source.n1010 10.4732
R830 source.n914 source.n896 10.4732
R831 source.n936 source.n886 10.4732
R832 source.n963 source.n874 10.4732
R833 source.n985 source.n864 10.4732
R834 source.n774 source.n756 10.4732
R835 source.n796 source.n746 10.4732
R836 source.n823 source.n734 10.4732
R837 source.n845 source.n724 10.4732
R838 source.n628 source.n610 10.4732
R839 source.n650 source.n600 10.4732
R840 source.n677 source.n588 10.4732
R841 source.n699 source.n578 10.4732
R842 source.n127 source.n6 10.4732
R843 source.n106 source.n17 10.4732
R844 source.n79 source.n29 10.4732
R845 source.n58 source.n40 10.4732
R846 source.n273 source.n152 10.4732
R847 source.n252 source.n163 10.4732
R848 source.n225 source.n175 10.4732
R849 source.n204 source.n186 10.4732
R850 source.n413 source.n292 10.4732
R851 source.n392 source.n303 10.4732
R852 source.n365 source.n315 10.4732
R853 source.n344 source.n326 10.4732
R854 source.n559 source.n438 10.4732
R855 source.n538 source.n449 10.4732
R856 source.n511 source.n461 10.4732
R857 source.n490 source.n472 10.4732
R858 source.n1049 source.n1048 10.2747
R859 source.n903 source.n902 10.2747
R860 source.n763 source.n762 10.2747
R861 source.n617 source.n616 10.2747
R862 source.n47 source.n46 10.2747
R863 source.n193 source.n192 10.2747
R864 source.n333 source.n332 10.2747
R865 source.n479 source.n478 10.2747
R866 source.n1059 source.n1044 9.69747
R867 source.n1086 source.n1085 9.69747
R868 source.n1106 source.n1105 9.69747
R869 source.n1132 source.n1008 9.69747
R870 source.n913 source.n898 9.69747
R871 source.n940 source.n939 9.69747
R872 source.n960 source.n959 9.69747
R873 source.n986 source.n862 9.69747
R874 source.n773 source.n758 9.69747
R875 source.n800 source.n799 9.69747
R876 source.n820 source.n819 9.69747
R877 source.n846 source.n722 9.69747
R878 source.n627 source.n612 9.69747
R879 source.n654 source.n653 9.69747
R880 source.n674 source.n673 9.69747
R881 source.n700 source.n576 9.69747
R882 source.n128 source.n4 9.69747
R883 source.n103 source.n102 9.69747
R884 source.n83 source.n82 9.69747
R885 source.n57 source.n42 9.69747
R886 source.n274 source.n150 9.69747
R887 source.n249 source.n248 9.69747
R888 source.n229 source.n228 9.69747
R889 source.n203 source.n188 9.69747
R890 source.n414 source.n290 9.69747
R891 source.n389 source.n388 9.69747
R892 source.n369 source.n368 9.69747
R893 source.n343 source.n328 9.69747
R894 source.n560 source.n436 9.69747
R895 source.n535 source.n534 9.69747
R896 source.n515 source.n514 9.69747
R897 source.n489 source.n474 9.69747
R898 source.n1142 source.n1141 9.45567
R899 source.n996 source.n995 9.45567
R900 source.n856 source.n855 9.45567
R901 source.n710 source.n709 9.45567
R902 source.n138 source.n137 9.45567
R903 source.n284 source.n283 9.45567
R904 source.n424 source.n423 9.45567
R905 source.n570 source.n569 9.45567
R906 source.n1006 source.n1005 9.3005
R907 source.n1135 source.n1134 9.3005
R908 source.n1133 source.n1132 9.3005
R909 source.n1010 source.n1009 9.3005
R910 source.n1127 source.n1126 9.3005
R911 source.n1125 source.n1124 9.3005
R912 source.n1014 source.n1013 9.3005
R913 source.n1093 source.n1092 9.3005
R914 source.n1091 source.n1090 9.3005
R915 source.n1030 source.n1029 9.3005
R916 source.n1085 source.n1084 9.3005
R917 source.n1083 source.n1082 9.3005
R918 source.n1034 source.n1033 9.3005
R919 source.n1077 source.n1076 9.3005
R920 source.n1075 source.n1074 9.3005
R921 source.n1051 source.n1050 9.3005
R922 source.n1046 source.n1045 9.3005
R923 source.n1057 source.n1056 9.3005
R924 source.n1059 source.n1058 9.3005
R925 source.n1042 source.n1041 9.3005
R926 source.n1065 source.n1064 9.3005
R927 source.n1067 source.n1066 9.3005
R928 source.n1068 source.n1037 9.3005
R929 source.n1026 source.n1025 9.3005
R930 source.n1099 source.n1098 9.3005
R931 source.n1101 source.n1100 9.3005
R932 source.n1022 source.n1021 9.3005
R933 source.n1107 source.n1106 9.3005
R934 source.n1109 source.n1108 9.3005
R935 source.n1018 source.n1017 9.3005
R936 source.n1116 source.n1115 9.3005
R937 source.n1118 source.n1117 9.3005
R938 source.n1141 source.n1140 9.3005
R939 source.n860 source.n859 9.3005
R940 source.n989 source.n988 9.3005
R941 source.n987 source.n986 9.3005
R942 source.n864 source.n863 9.3005
R943 source.n981 source.n980 9.3005
R944 source.n979 source.n978 9.3005
R945 source.n868 source.n867 9.3005
R946 source.n947 source.n946 9.3005
R947 source.n945 source.n944 9.3005
R948 source.n884 source.n883 9.3005
R949 source.n939 source.n938 9.3005
R950 source.n937 source.n936 9.3005
R951 source.n888 source.n887 9.3005
R952 source.n931 source.n930 9.3005
R953 source.n929 source.n928 9.3005
R954 source.n905 source.n904 9.3005
R955 source.n900 source.n899 9.3005
R956 source.n911 source.n910 9.3005
R957 source.n913 source.n912 9.3005
R958 source.n896 source.n895 9.3005
R959 source.n919 source.n918 9.3005
R960 source.n921 source.n920 9.3005
R961 source.n922 source.n891 9.3005
R962 source.n880 source.n879 9.3005
R963 source.n953 source.n952 9.3005
R964 source.n955 source.n954 9.3005
R965 source.n876 source.n875 9.3005
R966 source.n961 source.n960 9.3005
R967 source.n963 source.n962 9.3005
R968 source.n872 source.n871 9.3005
R969 source.n970 source.n969 9.3005
R970 source.n972 source.n971 9.3005
R971 source.n995 source.n994 9.3005
R972 source.n720 source.n719 9.3005
R973 source.n849 source.n848 9.3005
R974 source.n847 source.n846 9.3005
R975 source.n724 source.n723 9.3005
R976 source.n841 source.n840 9.3005
R977 source.n839 source.n838 9.3005
R978 source.n728 source.n727 9.3005
R979 source.n807 source.n806 9.3005
R980 source.n805 source.n804 9.3005
R981 source.n744 source.n743 9.3005
R982 source.n799 source.n798 9.3005
R983 source.n797 source.n796 9.3005
R984 source.n748 source.n747 9.3005
R985 source.n791 source.n790 9.3005
R986 source.n789 source.n788 9.3005
R987 source.n765 source.n764 9.3005
R988 source.n760 source.n759 9.3005
R989 source.n771 source.n770 9.3005
R990 source.n773 source.n772 9.3005
R991 source.n756 source.n755 9.3005
R992 source.n779 source.n778 9.3005
R993 source.n781 source.n780 9.3005
R994 source.n782 source.n751 9.3005
R995 source.n740 source.n739 9.3005
R996 source.n813 source.n812 9.3005
R997 source.n815 source.n814 9.3005
R998 source.n736 source.n735 9.3005
R999 source.n821 source.n820 9.3005
R1000 source.n823 source.n822 9.3005
R1001 source.n732 source.n731 9.3005
R1002 source.n830 source.n829 9.3005
R1003 source.n832 source.n831 9.3005
R1004 source.n855 source.n854 9.3005
R1005 source.n574 source.n573 9.3005
R1006 source.n703 source.n702 9.3005
R1007 source.n701 source.n700 9.3005
R1008 source.n578 source.n577 9.3005
R1009 source.n695 source.n694 9.3005
R1010 source.n693 source.n692 9.3005
R1011 source.n582 source.n581 9.3005
R1012 source.n661 source.n660 9.3005
R1013 source.n659 source.n658 9.3005
R1014 source.n598 source.n597 9.3005
R1015 source.n653 source.n652 9.3005
R1016 source.n651 source.n650 9.3005
R1017 source.n602 source.n601 9.3005
R1018 source.n645 source.n644 9.3005
R1019 source.n643 source.n642 9.3005
R1020 source.n619 source.n618 9.3005
R1021 source.n614 source.n613 9.3005
R1022 source.n625 source.n624 9.3005
R1023 source.n627 source.n626 9.3005
R1024 source.n610 source.n609 9.3005
R1025 source.n633 source.n632 9.3005
R1026 source.n635 source.n634 9.3005
R1027 source.n636 source.n605 9.3005
R1028 source.n594 source.n593 9.3005
R1029 source.n667 source.n666 9.3005
R1030 source.n669 source.n668 9.3005
R1031 source.n590 source.n589 9.3005
R1032 source.n675 source.n674 9.3005
R1033 source.n677 source.n676 9.3005
R1034 source.n586 source.n585 9.3005
R1035 source.n684 source.n683 9.3005
R1036 source.n686 source.n685 9.3005
R1037 source.n709 source.n708 9.3005
R1038 source.n49 source.n48 9.3005
R1039 source.n44 source.n43 9.3005
R1040 source.n55 source.n54 9.3005
R1041 source.n57 source.n56 9.3005
R1042 source.n40 source.n39 9.3005
R1043 source.n63 source.n62 9.3005
R1044 source.n65 source.n64 9.3005
R1045 source.n37 source.n34 9.3005
R1046 source.n96 source.n95 9.3005
R1047 source.n98 source.n97 9.3005
R1048 source.n19 source.n18 9.3005
R1049 source.n104 source.n103 9.3005
R1050 source.n106 source.n105 9.3005
R1051 source.n14 source.n13 9.3005
R1052 source.n112 source.n111 9.3005
R1053 source.n114 source.n113 9.3005
R1054 source.n137 source.n136 9.3005
R1055 source.n2 source.n1 9.3005
R1056 source.n131 source.n130 9.3005
R1057 source.n129 source.n128 9.3005
R1058 source.n6 source.n5 9.3005
R1059 source.n123 source.n122 9.3005
R1060 source.n121 source.n120 9.3005
R1061 source.n10 source.n9 9.3005
R1062 source.n23 source.n22 9.3005
R1063 source.n90 source.n89 9.3005
R1064 source.n88 source.n87 9.3005
R1065 source.n27 source.n26 9.3005
R1066 source.n82 source.n81 9.3005
R1067 source.n80 source.n79 9.3005
R1068 source.n31 source.n30 9.3005
R1069 source.n74 source.n73 9.3005
R1070 source.n72 source.n71 9.3005
R1071 source.n195 source.n194 9.3005
R1072 source.n190 source.n189 9.3005
R1073 source.n201 source.n200 9.3005
R1074 source.n203 source.n202 9.3005
R1075 source.n186 source.n185 9.3005
R1076 source.n209 source.n208 9.3005
R1077 source.n211 source.n210 9.3005
R1078 source.n183 source.n180 9.3005
R1079 source.n242 source.n241 9.3005
R1080 source.n244 source.n243 9.3005
R1081 source.n165 source.n164 9.3005
R1082 source.n250 source.n249 9.3005
R1083 source.n252 source.n251 9.3005
R1084 source.n160 source.n159 9.3005
R1085 source.n258 source.n257 9.3005
R1086 source.n260 source.n259 9.3005
R1087 source.n283 source.n282 9.3005
R1088 source.n148 source.n147 9.3005
R1089 source.n277 source.n276 9.3005
R1090 source.n275 source.n274 9.3005
R1091 source.n152 source.n151 9.3005
R1092 source.n269 source.n268 9.3005
R1093 source.n267 source.n266 9.3005
R1094 source.n156 source.n155 9.3005
R1095 source.n169 source.n168 9.3005
R1096 source.n236 source.n235 9.3005
R1097 source.n234 source.n233 9.3005
R1098 source.n173 source.n172 9.3005
R1099 source.n228 source.n227 9.3005
R1100 source.n226 source.n225 9.3005
R1101 source.n177 source.n176 9.3005
R1102 source.n220 source.n219 9.3005
R1103 source.n218 source.n217 9.3005
R1104 source.n335 source.n334 9.3005
R1105 source.n330 source.n329 9.3005
R1106 source.n341 source.n340 9.3005
R1107 source.n343 source.n342 9.3005
R1108 source.n326 source.n325 9.3005
R1109 source.n349 source.n348 9.3005
R1110 source.n351 source.n350 9.3005
R1111 source.n323 source.n320 9.3005
R1112 source.n382 source.n381 9.3005
R1113 source.n384 source.n383 9.3005
R1114 source.n305 source.n304 9.3005
R1115 source.n390 source.n389 9.3005
R1116 source.n392 source.n391 9.3005
R1117 source.n300 source.n299 9.3005
R1118 source.n398 source.n397 9.3005
R1119 source.n400 source.n399 9.3005
R1120 source.n423 source.n422 9.3005
R1121 source.n288 source.n287 9.3005
R1122 source.n417 source.n416 9.3005
R1123 source.n415 source.n414 9.3005
R1124 source.n292 source.n291 9.3005
R1125 source.n409 source.n408 9.3005
R1126 source.n407 source.n406 9.3005
R1127 source.n296 source.n295 9.3005
R1128 source.n309 source.n308 9.3005
R1129 source.n376 source.n375 9.3005
R1130 source.n374 source.n373 9.3005
R1131 source.n313 source.n312 9.3005
R1132 source.n368 source.n367 9.3005
R1133 source.n366 source.n365 9.3005
R1134 source.n317 source.n316 9.3005
R1135 source.n360 source.n359 9.3005
R1136 source.n358 source.n357 9.3005
R1137 source.n481 source.n480 9.3005
R1138 source.n476 source.n475 9.3005
R1139 source.n487 source.n486 9.3005
R1140 source.n489 source.n488 9.3005
R1141 source.n472 source.n471 9.3005
R1142 source.n495 source.n494 9.3005
R1143 source.n497 source.n496 9.3005
R1144 source.n469 source.n466 9.3005
R1145 source.n528 source.n527 9.3005
R1146 source.n530 source.n529 9.3005
R1147 source.n451 source.n450 9.3005
R1148 source.n536 source.n535 9.3005
R1149 source.n538 source.n537 9.3005
R1150 source.n446 source.n445 9.3005
R1151 source.n544 source.n543 9.3005
R1152 source.n546 source.n545 9.3005
R1153 source.n569 source.n568 9.3005
R1154 source.n434 source.n433 9.3005
R1155 source.n563 source.n562 9.3005
R1156 source.n561 source.n560 9.3005
R1157 source.n438 source.n437 9.3005
R1158 source.n555 source.n554 9.3005
R1159 source.n553 source.n552 9.3005
R1160 source.n442 source.n441 9.3005
R1161 source.n455 source.n454 9.3005
R1162 source.n522 source.n521 9.3005
R1163 source.n520 source.n519 9.3005
R1164 source.n459 source.n458 9.3005
R1165 source.n514 source.n513 9.3005
R1166 source.n512 source.n511 9.3005
R1167 source.n463 source.n462 9.3005
R1168 source.n506 source.n505 9.3005
R1169 source.n504 source.n503 9.3005
R1170 source.n1056 source.n1055 8.92171
R1171 source.n1089 source.n1030 8.92171
R1172 source.n1102 source.n1022 8.92171
R1173 source.n1136 source.n1135 8.92171
R1174 source.n910 source.n909 8.92171
R1175 source.n943 source.n884 8.92171
R1176 source.n956 source.n876 8.92171
R1177 source.n990 source.n989 8.92171
R1178 source.n770 source.n769 8.92171
R1179 source.n803 source.n744 8.92171
R1180 source.n816 source.n736 8.92171
R1181 source.n850 source.n849 8.92171
R1182 source.n624 source.n623 8.92171
R1183 source.n657 source.n598 8.92171
R1184 source.n670 source.n590 8.92171
R1185 source.n704 source.n703 8.92171
R1186 source.n132 source.n131 8.92171
R1187 source.n99 source.n19 8.92171
R1188 source.n86 source.n27 8.92171
R1189 source.n54 source.n53 8.92171
R1190 source.n278 source.n277 8.92171
R1191 source.n245 source.n165 8.92171
R1192 source.n232 source.n173 8.92171
R1193 source.n200 source.n199 8.92171
R1194 source.n418 source.n417 8.92171
R1195 source.n385 source.n305 8.92171
R1196 source.n372 source.n313 8.92171
R1197 source.n340 source.n339 8.92171
R1198 source.n564 source.n563 8.92171
R1199 source.n531 source.n451 8.92171
R1200 source.n518 source.n459 8.92171
R1201 source.n486 source.n485 8.92171
R1202 source.n1052 source.n1046 8.14595
R1203 source.n1090 source.n1028 8.14595
R1204 source.n1101 source.n1024 8.14595
R1205 source.n1139 source.n1006 8.14595
R1206 source.n906 source.n900 8.14595
R1207 source.n944 source.n882 8.14595
R1208 source.n955 source.n878 8.14595
R1209 source.n993 source.n860 8.14595
R1210 source.n766 source.n760 8.14595
R1211 source.n804 source.n742 8.14595
R1212 source.n815 source.n738 8.14595
R1213 source.n853 source.n720 8.14595
R1214 source.n620 source.n614 8.14595
R1215 source.n658 source.n596 8.14595
R1216 source.n669 source.n592 8.14595
R1217 source.n707 source.n574 8.14595
R1218 source.n135 source.n2 8.14595
R1219 source.n98 source.n21 8.14595
R1220 source.n87 source.n25 8.14595
R1221 source.n50 source.n44 8.14595
R1222 source.n281 source.n148 8.14595
R1223 source.n244 source.n167 8.14595
R1224 source.n233 source.n171 8.14595
R1225 source.n196 source.n190 8.14595
R1226 source.n421 source.n288 8.14595
R1227 source.n384 source.n307 8.14595
R1228 source.n373 source.n311 8.14595
R1229 source.n336 source.n330 8.14595
R1230 source.n567 source.n434 8.14595
R1231 source.n530 source.n453 8.14595
R1232 source.n519 source.n457 8.14595
R1233 source.n482 source.n476 8.14595
R1234 source.n1051 source.n1048 7.3702
R1235 source.n1094 source.n1093 7.3702
R1236 source.n1098 source.n1097 7.3702
R1237 source.n1140 source.n1004 7.3702
R1238 source.n905 source.n902 7.3702
R1239 source.n948 source.n947 7.3702
R1240 source.n952 source.n951 7.3702
R1241 source.n994 source.n858 7.3702
R1242 source.n765 source.n762 7.3702
R1243 source.n808 source.n807 7.3702
R1244 source.n812 source.n811 7.3702
R1245 source.n854 source.n718 7.3702
R1246 source.n619 source.n616 7.3702
R1247 source.n662 source.n661 7.3702
R1248 source.n666 source.n665 7.3702
R1249 source.n708 source.n572 7.3702
R1250 source.n136 source.n0 7.3702
R1251 source.n95 source.n94 7.3702
R1252 source.n91 source.n90 7.3702
R1253 source.n49 source.n46 7.3702
R1254 source.n282 source.n146 7.3702
R1255 source.n241 source.n240 7.3702
R1256 source.n237 source.n236 7.3702
R1257 source.n195 source.n192 7.3702
R1258 source.n422 source.n286 7.3702
R1259 source.n381 source.n380 7.3702
R1260 source.n377 source.n376 7.3702
R1261 source.n335 source.n332 7.3702
R1262 source.n568 source.n432 7.3702
R1263 source.n527 source.n526 7.3702
R1264 source.n523 source.n522 7.3702
R1265 source.n481 source.n478 7.3702
R1266 source.n1094 source.n1026 6.59444
R1267 source.n1097 source.n1026 6.59444
R1268 source.n1142 source.n1004 6.59444
R1269 source.n948 source.n880 6.59444
R1270 source.n951 source.n880 6.59444
R1271 source.n996 source.n858 6.59444
R1272 source.n808 source.n740 6.59444
R1273 source.n811 source.n740 6.59444
R1274 source.n856 source.n718 6.59444
R1275 source.n662 source.n594 6.59444
R1276 source.n665 source.n594 6.59444
R1277 source.n710 source.n572 6.59444
R1278 source.n138 source.n0 6.59444
R1279 source.n94 source.n23 6.59444
R1280 source.n91 source.n23 6.59444
R1281 source.n284 source.n146 6.59444
R1282 source.n240 source.n169 6.59444
R1283 source.n237 source.n169 6.59444
R1284 source.n424 source.n286 6.59444
R1285 source.n380 source.n309 6.59444
R1286 source.n377 source.n309 6.59444
R1287 source.n570 source.n432 6.59444
R1288 source.n526 source.n455 6.59444
R1289 source.n523 source.n455 6.59444
R1290 source.n1052 source.n1051 5.81868
R1291 source.n1093 source.n1028 5.81868
R1292 source.n1098 source.n1024 5.81868
R1293 source.n1140 source.n1139 5.81868
R1294 source.n906 source.n905 5.81868
R1295 source.n947 source.n882 5.81868
R1296 source.n952 source.n878 5.81868
R1297 source.n994 source.n993 5.81868
R1298 source.n766 source.n765 5.81868
R1299 source.n807 source.n742 5.81868
R1300 source.n812 source.n738 5.81868
R1301 source.n854 source.n853 5.81868
R1302 source.n620 source.n619 5.81868
R1303 source.n661 source.n596 5.81868
R1304 source.n666 source.n592 5.81868
R1305 source.n708 source.n707 5.81868
R1306 source.n136 source.n135 5.81868
R1307 source.n95 source.n21 5.81868
R1308 source.n90 source.n25 5.81868
R1309 source.n50 source.n49 5.81868
R1310 source.n282 source.n281 5.81868
R1311 source.n241 source.n167 5.81868
R1312 source.n236 source.n171 5.81868
R1313 source.n196 source.n195 5.81868
R1314 source.n422 source.n421 5.81868
R1315 source.n381 source.n307 5.81868
R1316 source.n376 source.n311 5.81868
R1317 source.n336 source.n335 5.81868
R1318 source.n568 source.n567 5.81868
R1319 source.n527 source.n453 5.81868
R1320 source.n522 source.n457 5.81868
R1321 source.n482 source.n481 5.81868
R1322 source.n1144 source.n1143 5.66429
R1323 source.n1055 source.n1046 5.04292
R1324 source.n1090 source.n1089 5.04292
R1325 source.n1102 source.n1101 5.04292
R1326 source.n1136 source.n1006 5.04292
R1327 source.n909 source.n900 5.04292
R1328 source.n944 source.n943 5.04292
R1329 source.n956 source.n955 5.04292
R1330 source.n990 source.n860 5.04292
R1331 source.n769 source.n760 5.04292
R1332 source.n804 source.n803 5.04292
R1333 source.n816 source.n815 5.04292
R1334 source.n850 source.n720 5.04292
R1335 source.n623 source.n614 5.04292
R1336 source.n658 source.n657 5.04292
R1337 source.n670 source.n669 5.04292
R1338 source.n704 source.n574 5.04292
R1339 source.n132 source.n2 5.04292
R1340 source.n99 source.n98 5.04292
R1341 source.n87 source.n86 5.04292
R1342 source.n53 source.n44 5.04292
R1343 source.n278 source.n148 5.04292
R1344 source.n245 source.n244 5.04292
R1345 source.n233 source.n232 5.04292
R1346 source.n199 source.n190 5.04292
R1347 source.n418 source.n288 5.04292
R1348 source.n385 source.n384 5.04292
R1349 source.n373 source.n372 5.04292
R1350 source.n339 source.n330 5.04292
R1351 source.n564 source.n434 5.04292
R1352 source.n531 source.n530 5.04292
R1353 source.n519 source.n518 5.04292
R1354 source.n485 source.n476 5.04292
R1355 source.n1056 source.n1044 4.26717
R1356 source.n1086 source.n1030 4.26717
R1357 source.n1105 source.n1022 4.26717
R1358 source.n1135 source.n1008 4.26717
R1359 source.n910 source.n898 4.26717
R1360 source.n940 source.n884 4.26717
R1361 source.n959 source.n876 4.26717
R1362 source.n989 source.n862 4.26717
R1363 source.n770 source.n758 4.26717
R1364 source.n800 source.n744 4.26717
R1365 source.n819 source.n736 4.26717
R1366 source.n849 source.n722 4.26717
R1367 source.n624 source.n612 4.26717
R1368 source.n654 source.n598 4.26717
R1369 source.n673 source.n590 4.26717
R1370 source.n703 source.n576 4.26717
R1371 source.n131 source.n4 4.26717
R1372 source.n102 source.n19 4.26717
R1373 source.n83 source.n27 4.26717
R1374 source.n54 source.n42 4.26717
R1375 source.n277 source.n150 4.26717
R1376 source.n248 source.n165 4.26717
R1377 source.n229 source.n173 4.26717
R1378 source.n200 source.n188 4.26717
R1379 source.n417 source.n290 4.26717
R1380 source.n388 source.n305 4.26717
R1381 source.n369 source.n313 4.26717
R1382 source.n340 source.n328 4.26717
R1383 source.n563 source.n436 4.26717
R1384 source.n534 source.n451 4.26717
R1385 source.n515 source.n459 4.26717
R1386 source.n486 source.n474 4.26717
R1387 source.n1060 source.n1059 3.49141
R1388 source.n1085 source.n1032 3.49141
R1389 source.n1106 source.n1020 3.49141
R1390 source.n1132 source.n1131 3.49141
R1391 source.n914 source.n913 3.49141
R1392 source.n939 source.n886 3.49141
R1393 source.n960 source.n874 3.49141
R1394 source.n986 source.n985 3.49141
R1395 source.n774 source.n773 3.49141
R1396 source.n799 source.n746 3.49141
R1397 source.n820 source.n734 3.49141
R1398 source.n846 source.n845 3.49141
R1399 source.n628 source.n627 3.49141
R1400 source.n653 source.n600 3.49141
R1401 source.n674 source.n588 3.49141
R1402 source.n700 source.n699 3.49141
R1403 source.n128 source.n127 3.49141
R1404 source.n103 source.n17 3.49141
R1405 source.n82 source.n29 3.49141
R1406 source.n58 source.n57 3.49141
R1407 source.n274 source.n273 3.49141
R1408 source.n249 source.n163 3.49141
R1409 source.n228 source.n175 3.49141
R1410 source.n204 source.n203 3.49141
R1411 source.n414 source.n413 3.49141
R1412 source.n389 source.n303 3.49141
R1413 source.n368 source.n315 3.49141
R1414 source.n344 source.n343 3.49141
R1415 source.n560 source.n559 3.49141
R1416 source.n535 source.n449 3.49141
R1417 source.n514 source.n461 3.49141
R1418 source.n490 source.n489 3.49141
R1419 source.n48 source.n47 2.84303
R1420 source.n194 source.n193 2.84303
R1421 source.n334 source.n333 2.84303
R1422 source.n480 source.n479 2.84303
R1423 source.n1050 source.n1049 2.84303
R1424 source.n904 source.n903 2.84303
R1425 source.n764 source.n763 2.84303
R1426 source.n618 source.n617 2.84303
R1427 source.n1063 source.n1042 2.71565
R1428 source.n1082 source.n1081 2.71565
R1429 source.n1110 source.n1109 2.71565
R1430 source.n1128 source.n1010 2.71565
R1431 source.n917 source.n896 2.71565
R1432 source.n936 source.n935 2.71565
R1433 source.n964 source.n963 2.71565
R1434 source.n982 source.n864 2.71565
R1435 source.n777 source.n756 2.71565
R1436 source.n796 source.n795 2.71565
R1437 source.n824 source.n823 2.71565
R1438 source.n842 source.n724 2.71565
R1439 source.n631 source.n610 2.71565
R1440 source.n650 source.n649 2.71565
R1441 source.n678 source.n677 2.71565
R1442 source.n696 source.n578 2.71565
R1443 source.n124 source.n6 2.71565
R1444 source.n107 source.n106 2.71565
R1445 source.n79 source.n78 2.71565
R1446 source.n61 source.n40 2.71565
R1447 source.n270 source.n152 2.71565
R1448 source.n253 source.n252 2.71565
R1449 source.n225 source.n224 2.71565
R1450 source.n207 source.n186 2.71565
R1451 source.n410 source.n292 2.71565
R1452 source.n393 source.n392 2.71565
R1453 source.n365 source.n364 2.71565
R1454 source.n347 source.n326 2.71565
R1455 source.n556 source.n438 2.71565
R1456 source.n539 source.n538 2.71565
R1457 source.n511 source.n510 2.71565
R1458 source.n493 source.n472 2.71565
R1459 source.n1064 source.n1040 1.93989
R1460 source.n1078 source.n1034 1.93989
R1461 source.n1114 source.n1018 1.93989
R1462 source.n1127 source.n1012 1.93989
R1463 source.n918 source.n894 1.93989
R1464 source.n932 source.n888 1.93989
R1465 source.n968 source.n872 1.93989
R1466 source.n981 source.n866 1.93989
R1467 source.n778 source.n754 1.93989
R1468 source.n792 source.n748 1.93989
R1469 source.n828 source.n732 1.93989
R1470 source.n841 source.n726 1.93989
R1471 source.n632 source.n608 1.93989
R1472 source.n646 source.n602 1.93989
R1473 source.n682 source.n586 1.93989
R1474 source.n695 source.n580 1.93989
R1475 source.n123 source.n8 1.93989
R1476 source.n110 source.n14 1.93989
R1477 source.n75 source.n31 1.93989
R1478 source.n62 source.n38 1.93989
R1479 source.n269 source.n154 1.93989
R1480 source.n256 source.n160 1.93989
R1481 source.n221 source.n177 1.93989
R1482 source.n208 source.n184 1.93989
R1483 source.n409 source.n294 1.93989
R1484 source.n396 source.n300 1.93989
R1485 source.n361 source.n317 1.93989
R1486 source.n348 source.n324 1.93989
R1487 source.n555 source.n440 1.93989
R1488 source.n542 source.n446 1.93989
R1489 source.n507 source.n463 1.93989
R1490 source.n494 source.n470 1.93989
R1491 source.n1069 source.n1067 1.16414
R1492 source.n1077 source.n1036 1.16414
R1493 source.n1115 source.n1016 1.16414
R1494 source.n1124 source.n1123 1.16414
R1495 source.n923 source.n921 1.16414
R1496 source.n931 source.n890 1.16414
R1497 source.n969 source.n870 1.16414
R1498 source.n978 source.n977 1.16414
R1499 source.n783 source.n781 1.16414
R1500 source.n791 source.n750 1.16414
R1501 source.n829 source.n730 1.16414
R1502 source.n838 source.n837 1.16414
R1503 source.n637 source.n635 1.16414
R1504 source.n645 source.n604 1.16414
R1505 source.n683 source.n584 1.16414
R1506 source.n692 source.n691 1.16414
R1507 source.n120 source.n119 1.16414
R1508 source.n111 source.n12 1.16414
R1509 source.n74 source.n33 1.16414
R1510 source.n66 source.n65 1.16414
R1511 source.n266 source.n265 1.16414
R1512 source.n257 source.n158 1.16414
R1513 source.n220 source.n179 1.16414
R1514 source.n212 source.n211 1.16414
R1515 source.n406 source.n405 1.16414
R1516 source.n397 source.n298 1.16414
R1517 source.n360 source.n319 1.16414
R1518 source.n352 source.n351 1.16414
R1519 source.n552 source.n551 1.16414
R1520 source.n543 source.n444 1.16414
R1521 source.n506 source.n465 1.16414
R1522 source.n498 source.n497 1.16414
R1523 source.n571 source.n431 0.802224
R1524 source.n431 source.n429 0.802224
R1525 source.n429 source.n427 0.802224
R1526 source.n427 source.n425 0.802224
R1527 source.n285 source.n145 0.802224
R1528 source.n145 source.n143 0.802224
R1529 source.n143 source.n141 0.802224
R1530 source.n141 source.n139 0.802224
R1531 source.n713 source.n711 0.802224
R1532 source.n715 source.n713 0.802224
R1533 source.n717 source.n715 0.802224
R1534 source.n857 source.n717 0.802224
R1535 source.n999 source.n997 0.802224
R1536 source.n1001 source.n999 0.802224
R1537 source.n1003 source.n1001 0.802224
R1538 source.n1143 source.n1003 0.802224
R1539 source.n1002 source.t9 0.7925
R1540 source.n1002 source.t7 0.7925
R1541 source.n1000 source.t5 0.7925
R1542 source.n1000 source.t14 0.7925
R1543 source.n998 source.t15 0.7925
R1544 source.n998 source.t8 0.7925
R1545 source.n716 source.t18 0.7925
R1546 source.n716 source.t23 0.7925
R1547 source.n714 source.t26 0.7925
R1548 source.n714 source.t31 0.7925
R1549 source.n712 source.t17 0.7925
R1550 source.n712 source.t25 0.7925
R1551 source.n140 source.t27 0.7925
R1552 source.n140 source.t28 0.7925
R1553 source.n142 source.t22 0.7925
R1554 source.n142 source.t24 0.7925
R1555 source.n144 source.t20 0.7925
R1556 source.n144 source.t21 0.7925
R1557 source.n426 source.t0 0.7925
R1558 source.n426 source.t12 0.7925
R1559 source.n428 source.t3 0.7925
R1560 source.n428 source.t11 0.7925
R1561 source.n430 source.t10 0.7925
R1562 source.n430 source.t4 0.7925
R1563 source.n425 source.n285 0.470328
R1564 source.n997 source.n857 0.470328
R1565 source.n1068 source.n1038 0.388379
R1566 source.n1074 source.n1073 0.388379
R1567 source.n1119 source.n1118 0.388379
R1568 source.n1120 source.n1014 0.388379
R1569 source.n922 source.n892 0.388379
R1570 source.n928 source.n927 0.388379
R1571 source.n973 source.n972 0.388379
R1572 source.n974 source.n868 0.388379
R1573 source.n782 source.n752 0.388379
R1574 source.n788 source.n787 0.388379
R1575 source.n833 source.n832 0.388379
R1576 source.n834 source.n728 0.388379
R1577 source.n636 source.n606 0.388379
R1578 source.n642 source.n641 0.388379
R1579 source.n687 source.n686 0.388379
R1580 source.n688 source.n582 0.388379
R1581 source.n116 source.n10 0.388379
R1582 source.n115 source.n114 0.388379
R1583 source.n71 source.n70 0.388379
R1584 source.n37 source.n35 0.388379
R1585 source.n262 source.n156 0.388379
R1586 source.n261 source.n260 0.388379
R1587 source.n217 source.n216 0.388379
R1588 source.n183 source.n181 0.388379
R1589 source.n402 source.n296 0.388379
R1590 source.n401 source.n400 0.388379
R1591 source.n357 source.n356 0.388379
R1592 source.n323 source.n321 0.388379
R1593 source.n548 source.n442 0.388379
R1594 source.n547 source.n546 0.388379
R1595 source.n503 source.n502 0.388379
R1596 source.n469 source.n467 0.388379
R1597 source source.n1144 0.188
R1598 source.n1050 source.n1045 0.155672
R1599 source.n1057 source.n1045 0.155672
R1600 source.n1058 source.n1057 0.155672
R1601 source.n1058 source.n1041 0.155672
R1602 source.n1065 source.n1041 0.155672
R1603 source.n1066 source.n1065 0.155672
R1604 source.n1066 source.n1037 0.155672
R1605 source.n1075 source.n1037 0.155672
R1606 source.n1076 source.n1075 0.155672
R1607 source.n1076 source.n1033 0.155672
R1608 source.n1083 source.n1033 0.155672
R1609 source.n1084 source.n1083 0.155672
R1610 source.n1084 source.n1029 0.155672
R1611 source.n1091 source.n1029 0.155672
R1612 source.n1092 source.n1091 0.155672
R1613 source.n1092 source.n1025 0.155672
R1614 source.n1099 source.n1025 0.155672
R1615 source.n1100 source.n1099 0.155672
R1616 source.n1100 source.n1021 0.155672
R1617 source.n1107 source.n1021 0.155672
R1618 source.n1108 source.n1107 0.155672
R1619 source.n1108 source.n1017 0.155672
R1620 source.n1116 source.n1017 0.155672
R1621 source.n1117 source.n1116 0.155672
R1622 source.n1117 source.n1013 0.155672
R1623 source.n1125 source.n1013 0.155672
R1624 source.n1126 source.n1125 0.155672
R1625 source.n1126 source.n1009 0.155672
R1626 source.n1133 source.n1009 0.155672
R1627 source.n1134 source.n1133 0.155672
R1628 source.n1134 source.n1005 0.155672
R1629 source.n1141 source.n1005 0.155672
R1630 source.n904 source.n899 0.155672
R1631 source.n911 source.n899 0.155672
R1632 source.n912 source.n911 0.155672
R1633 source.n912 source.n895 0.155672
R1634 source.n919 source.n895 0.155672
R1635 source.n920 source.n919 0.155672
R1636 source.n920 source.n891 0.155672
R1637 source.n929 source.n891 0.155672
R1638 source.n930 source.n929 0.155672
R1639 source.n930 source.n887 0.155672
R1640 source.n937 source.n887 0.155672
R1641 source.n938 source.n937 0.155672
R1642 source.n938 source.n883 0.155672
R1643 source.n945 source.n883 0.155672
R1644 source.n946 source.n945 0.155672
R1645 source.n946 source.n879 0.155672
R1646 source.n953 source.n879 0.155672
R1647 source.n954 source.n953 0.155672
R1648 source.n954 source.n875 0.155672
R1649 source.n961 source.n875 0.155672
R1650 source.n962 source.n961 0.155672
R1651 source.n962 source.n871 0.155672
R1652 source.n970 source.n871 0.155672
R1653 source.n971 source.n970 0.155672
R1654 source.n971 source.n867 0.155672
R1655 source.n979 source.n867 0.155672
R1656 source.n980 source.n979 0.155672
R1657 source.n980 source.n863 0.155672
R1658 source.n987 source.n863 0.155672
R1659 source.n988 source.n987 0.155672
R1660 source.n988 source.n859 0.155672
R1661 source.n995 source.n859 0.155672
R1662 source.n764 source.n759 0.155672
R1663 source.n771 source.n759 0.155672
R1664 source.n772 source.n771 0.155672
R1665 source.n772 source.n755 0.155672
R1666 source.n779 source.n755 0.155672
R1667 source.n780 source.n779 0.155672
R1668 source.n780 source.n751 0.155672
R1669 source.n789 source.n751 0.155672
R1670 source.n790 source.n789 0.155672
R1671 source.n790 source.n747 0.155672
R1672 source.n797 source.n747 0.155672
R1673 source.n798 source.n797 0.155672
R1674 source.n798 source.n743 0.155672
R1675 source.n805 source.n743 0.155672
R1676 source.n806 source.n805 0.155672
R1677 source.n806 source.n739 0.155672
R1678 source.n813 source.n739 0.155672
R1679 source.n814 source.n813 0.155672
R1680 source.n814 source.n735 0.155672
R1681 source.n821 source.n735 0.155672
R1682 source.n822 source.n821 0.155672
R1683 source.n822 source.n731 0.155672
R1684 source.n830 source.n731 0.155672
R1685 source.n831 source.n830 0.155672
R1686 source.n831 source.n727 0.155672
R1687 source.n839 source.n727 0.155672
R1688 source.n840 source.n839 0.155672
R1689 source.n840 source.n723 0.155672
R1690 source.n847 source.n723 0.155672
R1691 source.n848 source.n847 0.155672
R1692 source.n848 source.n719 0.155672
R1693 source.n855 source.n719 0.155672
R1694 source.n618 source.n613 0.155672
R1695 source.n625 source.n613 0.155672
R1696 source.n626 source.n625 0.155672
R1697 source.n626 source.n609 0.155672
R1698 source.n633 source.n609 0.155672
R1699 source.n634 source.n633 0.155672
R1700 source.n634 source.n605 0.155672
R1701 source.n643 source.n605 0.155672
R1702 source.n644 source.n643 0.155672
R1703 source.n644 source.n601 0.155672
R1704 source.n651 source.n601 0.155672
R1705 source.n652 source.n651 0.155672
R1706 source.n652 source.n597 0.155672
R1707 source.n659 source.n597 0.155672
R1708 source.n660 source.n659 0.155672
R1709 source.n660 source.n593 0.155672
R1710 source.n667 source.n593 0.155672
R1711 source.n668 source.n667 0.155672
R1712 source.n668 source.n589 0.155672
R1713 source.n675 source.n589 0.155672
R1714 source.n676 source.n675 0.155672
R1715 source.n676 source.n585 0.155672
R1716 source.n684 source.n585 0.155672
R1717 source.n685 source.n684 0.155672
R1718 source.n685 source.n581 0.155672
R1719 source.n693 source.n581 0.155672
R1720 source.n694 source.n693 0.155672
R1721 source.n694 source.n577 0.155672
R1722 source.n701 source.n577 0.155672
R1723 source.n702 source.n701 0.155672
R1724 source.n702 source.n573 0.155672
R1725 source.n709 source.n573 0.155672
R1726 source.n137 source.n1 0.155672
R1727 source.n130 source.n1 0.155672
R1728 source.n130 source.n129 0.155672
R1729 source.n129 source.n5 0.155672
R1730 source.n122 source.n5 0.155672
R1731 source.n122 source.n121 0.155672
R1732 source.n121 source.n9 0.155672
R1733 source.n113 source.n9 0.155672
R1734 source.n113 source.n112 0.155672
R1735 source.n112 source.n13 0.155672
R1736 source.n105 source.n13 0.155672
R1737 source.n105 source.n104 0.155672
R1738 source.n104 source.n18 0.155672
R1739 source.n97 source.n18 0.155672
R1740 source.n97 source.n96 0.155672
R1741 source.n96 source.n22 0.155672
R1742 source.n89 source.n22 0.155672
R1743 source.n89 source.n88 0.155672
R1744 source.n88 source.n26 0.155672
R1745 source.n81 source.n26 0.155672
R1746 source.n81 source.n80 0.155672
R1747 source.n80 source.n30 0.155672
R1748 source.n73 source.n30 0.155672
R1749 source.n73 source.n72 0.155672
R1750 source.n72 source.n34 0.155672
R1751 source.n64 source.n34 0.155672
R1752 source.n64 source.n63 0.155672
R1753 source.n63 source.n39 0.155672
R1754 source.n56 source.n39 0.155672
R1755 source.n56 source.n55 0.155672
R1756 source.n55 source.n43 0.155672
R1757 source.n48 source.n43 0.155672
R1758 source.n283 source.n147 0.155672
R1759 source.n276 source.n147 0.155672
R1760 source.n276 source.n275 0.155672
R1761 source.n275 source.n151 0.155672
R1762 source.n268 source.n151 0.155672
R1763 source.n268 source.n267 0.155672
R1764 source.n267 source.n155 0.155672
R1765 source.n259 source.n155 0.155672
R1766 source.n259 source.n258 0.155672
R1767 source.n258 source.n159 0.155672
R1768 source.n251 source.n159 0.155672
R1769 source.n251 source.n250 0.155672
R1770 source.n250 source.n164 0.155672
R1771 source.n243 source.n164 0.155672
R1772 source.n243 source.n242 0.155672
R1773 source.n242 source.n168 0.155672
R1774 source.n235 source.n168 0.155672
R1775 source.n235 source.n234 0.155672
R1776 source.n234 source.n172 0.155672
R1777 source.n227 source.n172 0.155672
R1778 source.n227 source.n226 0.155672
R1779 source.n226 source.n176 0.155672
R1780 source.n219 source.n176 0.155672
R1781 source.n219 source.n218 0.155672
R1782 source.n218 source.n180 0.155672
R1783 source.n210 source.n180 0.155672
R1784 source.n210 source.n209 0.155672
R1785 source.n209 source.n185 0.155672
R1786 source.n202 source.n185 0.155672
R1787 source.n202 source.n201 0.155672
R1788 source.n201 source.n189 0.155672
R1789 source.n194 source.n189 0.155672
R1790 source.n423 source.n287 0.155672
R1791 source.n416 source.n287 0.155672
R1792 source.n416 source.n415 0.155672
R1793 source.n415 source.n291 0.155672
R1794 source.n408 source.n291 0.155672
R1795 source.n408 source.n407 0.155672
R1796 source.n407 source.n295 0.155672
R1797 source.n399 source.n295 0.155672
R1798 source.n399 source.n398 0.155672
R1799 source.n398 source.n299 0.155672
R1800 source.n391 source.n299 0.155672
R1801 source.n391 source.n390 0.155672
R1802 source.n390 source.n304 0.155672
R1803 source.n383 source.n304 0.155672
R1804 source.n383 source.n382 0.155672
R1805 source.n382 source.n308 0.155672
R1806 source.n375 source.n308 0.155672
R1807 source.n375 source.n374 0.155672
R1808 source.n374 source.n312 0.155672
R1809 source.n367 source.n312 0.155672
R1810 source.n367 source.n366 0.155672
R1811 source.n366 source.n316 0.155672
R1812 source.n359 source.n316 0.155672
R1813 source.n359 source.n358 0.155672
R1814 source.n358 source.n320 0.155672
R1815 source.n350 source.n320 0.155672
R1816 source.n350 source.n349 0.155672
R1817 source.n349 source.n325 0.155672
R1818 source.n342 source.n325 0.155672
R1819 source.n342 source.n341 0.155672
R1820 source.n341 source.n329 0.155672
R1821 source.n334 source.n329 0.155672
R1822 source.n569 source.n433 0.155672
R1823 source.n562 source.n433 0.155672
R1824 source.n562 source.n561 0.155672
R1825 source.n561 source.n437 0.155672
R1826 source.n554 source.n437 0.155672
R1827 source.n554 source.n553 0.155672
R1828 source.n553 source.n441 0.155672
R1829 source.n545 source.n441 0.155672
R1830 source.n545 source.n544 0.155672
R1831 source.n544 source.n445 0.155672
R1832 source.n537 source.n445 0.155672
R1833 source.n537 source.n536 0.155672
R1834 source.n536 source.n450 0.155672
R1835 source.n529 source.n450 0.155672
R1836 source.n529 source.n528 0.155672
R1837 source.n528 source.n454 0.155672
R1838 source.n521 source.n454 0.155672
R1839 source.n521 source.n520 0.155672
R1840 source.n520 source.n458 0.155672
R1841 source.n513 source.n458 0.155672
R1842 source.n513 source.n512 0.155672
R1843 source.n512 source.n462 0.155672
R1844 source.n505 source.n462 0.155672
R1845 source.n505 source.n504 0.155672
R1846 source.n504 source.n466 0.155672
R1847 source.n496 source.n466 0.155672
R1848 source.n496 source.n495 0.155672
R1849 source.n495 source.n471 0.155672
R1850 source.n488 source.n471 0.155672
R1851 source.n488 source.n487 0.155672
R1852 source.n487 source.n475 0.155672
R1853 source.n480 source.n475 0.155672
R1854 minus.n6 minus.t11 1090.62
R1855 minus.n30 minus.t13 1090.62
R1856 minus.n5 minus.t10 1069.64
R1857 minus.n9 minus.t9 1069.64
R1858 minus.n3 minus.t8 1069.64
R1859 minus.n15 minus.t4 1069.64
R1860 minus.n1 minus.t6 1069.64
R1861 minus.n21 minus.t5 1069.64
R1862 minus.n22 minus.t1 1069.64
R1863 minus.n29 minus.t3 1069.64
R1864 minus.n33 minus.t7 1069.64
R1865 minus.n27 minus.t15 1069.64
R1866 minus.n39 minus.t2 1069.64
R1867 minus.n25 minus.t0 1069.64
R1868 minus.n45 minus.t12 1069.64
R1869 minus.n46 minus.t14 1069.64
R1870 minus.n23 minus.n22 161.3
R1871 minus.n21 minus.n0 161.3
R1872 minus.n20 minus.n19 161.3
R1873 minus.n18 minus.n1 161.3
R1874 minus.n17 minus.n16 161.3
R1875 minus.n15 minus.n2 161.3
R1876 minus.n14 minus.n13 161.3
R1877 minus.n12 minus.n3 161.3
R1878 minus.n11 minus.n10 161.3
R1879 minus.n9 minus.n4 161.3
R1880 minus.n8 minus.n7 161.3
R1881 minus.n47 minus.n46 161.3
R1882 minus.n45 minus.n24 161.3
R1883 minus.n44 minus.n43 161.3
R1884 minus.n42 minus.n25 161.3
R1885 minus.n41 minus.n40 161.3
R1886 minus.n39 minus.n26 161.3
R1887 minus.n38 minus.n37 161.3
R1888 minus.n36 minus.n27 161.3
R1889 minus.n35 minus.n34 161.3
R1890 minus.n33 minus.n28 161.3
R1891 minus.n32 minus.n31 161.3
R1892 minus.n7 minus.n6 70.4033
R1893 minus.n31 minus.n30 70.4033
R1894 minus.n22 minus.n21 48.2005
R1895 minus.n46 minus.n45 48.2005
R1896 minus.n48 minus.n23 48.1785
R1897 minus.n9 minus.n8 44.549
R1898 minus.n20 minus.n1 44.549
R1899 minus.n33 minus.n32 44.549
R1900 minus.n44 minus.n25 44.549
R1901 minus.n10 minus.n3 34.3247
R1902 minus.n16 minus.n15 34.3247
R1903 minus.n34 minus.n27 34.3247
R1904 minus.n40 minus.n39 34.3247
R1905 minus.n15 minus.n14 24.1005
R1906 minus.n14 minus.n3 24.1005
R1907 minus.n38 minus.n27 24.1005
R1908 minus.n39 minus.n38 24.1005
R1909 minus.n6 minus.n5 20.9576
R1910 minus.n30 minus.n29 20.9576
R1911 minus.n10 minus.n9 13.8763
R1912 minus.n16 minus.n1 13.8763
R1913 minus.n34 minus.n33 13.8763
R1914 minus.n40 minus.n25 13.8763
R1915 minus.n48 minus.n47 6.6558
R1916 minus.n8 minus.n5 3.65202
R1917 minus.n21 minus.n20 3.65202
R1918 minus.n32 minus.n29 3.65202
R1919 minus.n45 minus.n44 3.65202
R1920 minus.n23 minus.n0 0.189894
R1921 minus.n19 minus.n0 0.189894
R1922 minus.n19 minus.n18 0.189894
R1923 minus.n18 minus.n17 0.189894
R1924 minus.n17 minus.n2 0.189894
R1925 minus.n13 minus.n2 0.189894
R1926 minus.n13 minus.n12 0.189894
R1927 minus.n12 minus.n11 0.189894
R1928 minus.n11 minus.n4 0.189894
R1929 minus.n7 minus.n4 0.189894
R1930 minus.n31 minus.n28 0.189894
R1931 minus.n35 minus.n28 0.189894
R1932 minus.n36 minus.n35 0.189894
R1933 minus.n37 minus.n36 0.189894
R1934 minus.n37 minus.n26 0.189894
R1935 minus.n41 minus.n26 0.189894
R1936 minus.n42 minus.n41 0.189894
R1937 minus.n43 minus.n42 0.189894
R1938 minus.n43 minus.n24 0.189894
R1939 minus.n47 minus.n24 0.189894
R1940 minus minus.n48 0.188
R1941 drain_right.n5 drain_right.n3 59.5172
R1942 drain_right.n2 drain_right.n0 59.5172
R1943 drain_right.n9 drain_right.n7 59.517
R1944 drain_right.n5 drain_right.n4 58.7154
R1945 drain_right.n2 drain_right.n1 58.7154
R1946 drain_right.n9 drain_right.n8 58.7154
R1947 drain_right.n11 drain_right.n10 58.7154
R1948 drain_right.n13 drain_right.n12 58.7154
R1949 drain_right drain_right.n6 41.8735
R1950 drain_right drain_right.n13 6.45494
R1951 drain_right.n13 drain_right.n11 0.802224
R1952 drain_right.n11 drain_right.n9 0.802224
R1953 drain_right.n3 drain_right.t3 0.7925
R1954 drain_right.n3 drain_right.t1 0.7925
R1955 drain_right.n4 drain_right.t13 0.7925
R1956 drain_right.n4 drain_right.t15 0.7925
R1957 drain_right.n1 drain_right.t8 0.7925
R1958 drain_right.n1 drain_right.t0 0.7925
R1959 drain_right.n0 drain_right.t2 0.7925
R1960 drain_right.n0 drain_right.t12 0.7925
R1961 drain_right.n7 drain_right.t5 0.7925
R1962 drain_right.n7 drain_right.t4 0.7925
R1963 drain_right.n8 drain_right.t7 0.7925
R1964 drain_right.n8 drain_right.t6 0.7925
R1965 drain_right.n10 drain_right.t9 0.7925
R1966 drain_right.n10 drain_right.t11 0.7925
R1967 drain_right.n12 drain_right.t14 0.7925
R1968 drain_right.n12 drain_right.t10 0.7925
R1969 drain_right.n6 drain_right.n5 0.346016
R1970 drain_right.n6 drain_right.n2 0.346016
C0 minus plus 8.531651f
C1 drain_left plus 19.1241f
C2 minus drain_left 0.172752f
C3 source drain_right 41.0365f
C4 drain_right plus 0.391974f
C5 minus drain_right 18.888199f
C6 drain_left drain_right 1.24373f
C7 source plus 18.357698f
C8 minus source 18.3437f
C9 source drain_left 41.034798f
C10 drain_right a_n2390_n5888# 9.07189f
C11 drain_left a_n2390_n5888# 9.41079f
C12 source a_n2390_n5888# 16.398415f
C13 minus a_n2390_n5888# 10.359813f
C14 plus a_n2390_n5888# 12.85349f
C15 drain_right.t2 a_n2390_n5888# 0.5564f
C16 drain_right.t12 a_n2390_n5888# 0.5564f
C17 drain_right.n0 a_n2390_n5888# 5.13315f
C18 drain_right.t8 a_n2390_n5888# 0.5564f
C19 drain_right.t0 a_n2390_n5888# 0.5564f
C20 drain_right.n1 a_n2390_n5888# 5.12783f
C21 drain_right.n2 a_n2390_n5888# 0.733675f
C22 drain_right.t3 a_n2390_n5888# 0.5564f
C23 drain_right.t1 a_n2390_n5888# 0.5564f
C24 drain_right.n3 a_n2390_n5888# 5.13315f
C25 drain_right.t13 a_n2390_n5888# 0.5564f
C26 drain_right.t15 a_n2390_n5888# 0.5564f
C27 drain_right.n4 a_n2390_n5888# 5.12783f
C28 drain_right.n5 a_n2390_n5888# 0.733675f
C29 drain_right.n6 a_n2390_n5888# 2.42265f
C30 drain_right.t5 a_n2390_n5888# 0.5564f
C31 drain_right.t4 a_n2390_n5888# 0.5564f
C32 drain_right.n7 a_n2390_n5888# 5.13314f
C33 drain_right.t7 a_n2390_n5888# 0.5564f
C34 drain_right.t6 a_n2390_n5888# 0.5564f
C35 drain_right.n8 a_n2390_n5888# 5.12783f
C36 drain_right.n9 a_n2390_n5888# 0.773196f
C37 drain_right.t9 a_n2390_n5888# 0.5564f
C38 drain_right.t11 a_n2390_n5888# 0.5564f
C39 drain_right.n10 a_n2390_n5888# 5.12783f
C40 drain_right.n11 a_n2390_n5888# 0.38358f
C41 drain_right.t14 a_n2390_n5888# 0.5564f
C42 drain_right.t10 a_n2390_n5888# 0.5564f
C43 drain_right.n12 a_n2390_n5888# 5.12783f
C44 drain_right.n13 a_n2390_n5888# 0.629167f
C45 minus.n0 a_n2390_n5888# 0.042353f
C46 minus.t6 a_n2390_n5888# 1.79536f
C47 minus.n1 a_n2390_n5888# 0.659267f
C48 minus.n2 a_n2390_n5888# 0.042353f
C49 minus.t8 a_n2390_n5888# 1.79536f
C50 minus.n3 a_n2390_n5888# 0.659267f
C51 minus.n4 a_n2390_n5888# 0.042353f
C52 minus.t10 a_n2390_n5888# 1.79536f
C53 minus.n5 a_n2390_n5888# 0.658092f
C54 minus.t11 a_n2390_n5888# 1.80801f
C55 minus.n6 a_n2390_n5888# 0.645129f
C56 minus.n7 a_n2390_n5888# 0.142649f
C57 minus.n8 a_n2390_n5888# 0.009611f
C58 minus.t9 a_n2390_n5888# 1.79536f
C59 minus.n9 a_n2390_n5888# 0.659267f
C60 minus.n10 a_n2390_n5888# 0.009611f
C61 minus.n11 a_n2390_n5888# 0.042353f
C62 minus.n12 a_n2390_n5888# 0.042353f
C63 minus.n13 a_n2390_n5888# 0.042353f
C64 minus.n14 a_n2390_n5888# 0.009611f
C65 minus.t4 a_n2390_n5888# 1.79536f
C66 minus.n15 a_n2390_n5888# 0.659267f
C67 minus.n16 a_n2390_n5888# 0.009611f
C68 minus.n17 a_n2390_n5888# 0.042353f
C69 minus.n18 a_n2390_n5888# 0.042353f
C70 minus.n19 a_n2390_n5888# 0.042353f
C71 minus.n20 a_n2390_n5888# 0.009611f
C72 minus.t5 a_n2390_n5888# 1.79536f
C73 minus.n21 a_n2390_n5888# 0.658092f
C74 minus.t1 a_n2390_n5888# 1.79536f
C75 minus.n22 a_n2390_n5888# 0.65744f
C76 minus.n23 a_n2390_n5888# 2.28832f
C77 minus.n24 a_n2390_n5888# 0.042353f
C78 minus.t0 a_n2390_n5888# 1.79536f
C79 minus.n25 a_n2390_n5888# 0.659267f
C80 minus.n26 a_n2390_n5888# 0.042353f
C81 minus.t15 a_n2390_n5888# 1.79536f
C82 minus.n27 a_n2390_n5888# 0.659267f
C83 minus.n28 a_n2390_n5888# 0.042353f
C84 minus.t3 a_n2390_n5888# 1.79536f
C85 minus.n29 a_n2390_n5888# 0.658092f
C86 minus.t13 a_n2390_n5888# 1.80801f
C87 minus.n30 a_n2390_n5888# 0.645129f
C88 minus.n31 a_n2390_n5888# 0.142649f
C89 minus.n32 a_n2390_n5888# 0.009611f
C90 minus.t7 a_n2390_n5888# 1.79536f
C91 minus.n33 a_n2390_n5888# 0.659267f
C92 minus.n34 a_n2390_n5888# 0.009611f
C93 minus.n35 a_n2390_n5888# 0.042353f
C94 minus.n36 a_n2390_n5888# 0.042353f
C95 minus.n37 a_n2390_n5888# 0.042353f
C96 minus.n38 a_n2390_n5888# 0.009611f
C97 minus.t2 a_n2390_n5888# 1.79536f
C98 minus.n39 a_n2390_n5888# 0.659267f
C99 minus.n40 a_n2390_n5888# 0.009611f
C100 minus.n41 a_n2390_n5888# 0.042353f
C101 minus.n42 a_n2390_n5888# 0.042353f
C102 minus.n43 a_n2390_n5888# 0.042353f
C103 minus.n44 a_n2390_n5888# 0.009611f
C104 minus.t12 a_n2390_n5888# 1.79536f
C105 minus.n45 a_n2390_n5888# 0.658092f
C106 minus.t14 a_n2390_n5888# 1.79536f
C107 minus.n46 a_n2390_n5888# 0.65744f
C108 minus.n47 a_n2390_n5888# 0.292328f
C109 minus.n48 a_n2390_n5888# 2.68512f
C110 source.n0 a_n2390_n5888# 0.031706f
C111 source.n1 a_n2390_n5888# 0.022999f
C112 source.n2 a_n2390_n5888# 0.012359f
C113 source.n3 a_n2390_n5888# 0.029211f
C114 source.n4 a_n2390_n5888# 0.013086f
C115 source.n5 a_n2390_n5888# 0.022999f
C116 source.n6 a_n2390_n5888# 0.012359f
C117 source.n7 a_n2390_n5888# 0.029211f
C118 source.n8 a_n2390_n5888# 0.013086f
C119 source.n9 a_n2390_n5888# 0.022999f
C120 source.n10 a_n2390_n5888# 0.012359f
C121 source.n11 a_n2390_n5888# 0.029211f
C122 source.n12 a_n2390_n5888# 0.013086f
C123 source.n13 a_n2390_n5888# 0.022999f
C124 source.n14 a_n2390_n5888# 0.012359f
C125 source.n15 a_n2390_n5888# 0.029211f
C126 source.n16 a_n2390_n5888# 0.029211f
C127 source.n17 a_n2390_n5888# 0.013086f
C128 source.n18 a_n2390_n5888# 0.022999f
C129 source.n19 a_n2390_n5888# 0.012359f
C130 source.n20 a_n2390_n5888# 0.029211f
C131 source.n21 a_n2390_n5888# 0.013086f
C132 source.n22 a_n2390_n5888# 0.022999f
C133 source.n23 a_n2390_n5888# 0.012359f
C134 source.n24 a_n2390_n5888# 0.029211f
C135 source.n25 a_n2390_n5888# 0.013086f
C136 source.n26 a_n2390_n5888# 0.022999f
C137 source.n27 a_n2390_n5888# 0.012359f
C138 source.n28 a_n2390_n5888# 0.029211f
C139 source.n29 a_n2390_n5888# 0.013086f
C140 source.n30 a_n2390_n5888# 0.022999f
C141 source.n31 a_n2390_n5888# 0.012359f
C142 source.n32 a_n2390_n5888# 0.029211f
C143 source.n33 a_n2390_n5888# 0.013086f
C144 source.n34 a_n2390_n5888# 0.022999f
C145 source.n35 a_n2390_n5888# 0.012722f
C146 source.n36 a_n2390_n5888# 0.029211f
C147 source.n37 a_n2390_n5888# 0.012359f
C148 source.n38 a_n2390_n5888# 0.013086f
C149 source.n39 a_n2390_n5888# 0.022999f
C150 source.n40 a_n2390_n5888# 0.012359f
C151 source.n41 a_n2390_n5888# 0.029211f
C152 source.n42 a_n2390_n5888# 0.013086f
C153 source.n43 a_n2390_n5888# 0.022999f
C154 source.n44 a_n2390_n5888# 0.012359f
C155 source.n45 a_n2390_n5888# 0.021909f
C156 source.n46 a_n2390_n5888# 0.02065f
C157 source.t29 a_n2390_n5888# 0.050946f
C158 source.n47 a_n2390_n5888# 0.280606f
C159 source.n48 a_n2390_n5888# 2.49011f
C160 source.n49 a_n2390_n5888# 0.012359f
C161 source.n50 a_n2390_n5888# 0.013086f
C162 source.n51 a_n2390_n5888# 0.029211f
C163 source.n52 a_n2390_n5888# 0.029211f
C164 source.n53 a_n2390_n5888# 0.013086f
C165 source.n54 a_n2390_n5888# 0.012359f
C166 source.n55 a_n2390_n5888# 0.022999f
C167 source.n56 a_n2390_n5888# 0.022999f
C168 source.n57 a_n2390_n5888# 0.012359f
C169 source.n58 a_n2390_n5888# 0.013086f
C170 source.n59 a_n2390_n5888# 0.029211f
C171 source.n60 a_n2390_n5888# 0.029211f
C172 source.n61 a_n2390_n5888# 0.013086f
C173 source.n62 a_n2390_n5888# 0.012359f
C174 source.n63 a_n2390_n5888# 0.022999f
C175 source.n64 a_n2390_n5888# 0.022999f
C176 source.n65 a_n2390_n5888# 0.012359f
C177 source.n66 a_n2390_n5888# 0.013086f
C178 source.n67 a_n2390_n5888# 0.029211f
C179 source.n68 a_n2390_n5888# 0.029211f
C180 source.n69 a_n2390_n5888# 0.029211f
C181 source.n70 a_n2390_n5888# 0.012722f
C182 source.n71 a_n2390_n5888# 0.012359f
C183 source.n72 a_n2390_n5888# 0.022999f
C184 source.n73 a_n2390_n5888# 0.022999f
C185 source.n74 a_n2390_n5888# 0.012359f
C186 source.n75 a_n2390_n5888# 0.013086f
C187 source.n76 a_n2390_n5888# 0.029211f
C188 source.n77 a_n2390_n5888# 0.029211f
C189 source.n78 a_n2390_n5888# 0.013086f
C190 source.n79 a_n2390_n5888# 0.012359f
C191 source.n80 a_n2390_n5888# 0.022999f
C192 source.n81 a_n2390_n5888# 0.022999f
C193 source.n82 a_n2390_n5888# 0.012359f
C194 source.n83 a_n2390_n5888# 0.013086f
C195 source.n84 a_n2390_n5888# 0.029211f
C196 source.n85 a_n2390_n5888# 0.029211f
C197 source.n86 a_n2390_n5888# 0.013086f
C198 source.n87 a_n2390_n5888# 0.012359f
C199 source.n88 a_n2390_n5888# 0.022999f
C200 source.n89 a_n2390_n5888# 0.022999f
C201 source.n90 a_n2390_n5888# 0.012359f
C202 source.n91 a_n2390_n5888# 0.013086f
C203 source.n92 a_n2390_n5888# 0.029211f
C204 source.n93 a_n2390_n5888# 0.029211f
C205 source.n94 a_n2390_n5888# 0.013086f
C206 source.n95 a_n2390_n5888# 0.012359f
C207 source.n96 a_n2390_n5888# 0.022999f
C208 source.n97 a_n2390_n5888# 0.022999f
C209 source.n98 a_n2390_n5888# 0.012359f
C210 source.n99 a_n2390_n5888# 0.013086f
C211 source.n100 a_n2390_n5888# 0.029211f
C212 source.n101 a_n2390_n5888# 0.029211f
C213 source.n102 a_n2390_n5888# 0.013086f
C214 source.n103 a_n2390_n5888# 0.012359f
C215 source.n104 a_n2390_n5888# 0.022999f
C216 source.n105 a_n2390_n5888# 0.022999f
C217 source.n106 a_n2390_n5888# 0.012359f
C218 source.n107 a_n2390_n5888# 0.013086f
C219 source.n108 a_n2390_n5888# 0.029211f
C220 source.n109 a_n2390_n5888# 0.029211f
C221 source.n110 a_n2390_n5888# 0.013086f
C222 source.n111 a_n2390_n5888# 0.012359f
C223 source.n112 a_n2390_n5888# 0.022999f
C224 source.n113 a_n2390_n5888# 0.022999f
C225 source.n114 a_n2390_n5888# 0.012359f
C226 source.n115 a_n2390_n5888# 0.012722f
C227 source.n116 a_n2390_n5888# 0.012722f
C228 source.n117 a_n2390_n5888# 0.029211f
C229 source.n118 a_n2390_n5888# 0.029211f
C230 source.n119 a_n2390_n5888# 0.013086f
C231 source.n120 a_n2390_n5888# 0.012359f
C232 source.n121 a_n2390_n5888# 0.022999f
C233 source.n122 a_n2390_n5888# 0.022999f
C234 source.n123 a_n2390_n5888# 0.012359f
C235 source.n124 a_n2390_n5888# 0.013086f
C236 source.n125 a_n2390_n5888# 0.029211f
C237 source.n126 a_n2390_n5888# 0.029211f
C238 source.n127 a_n2390_n5888# 0.013086f
C239 source.n128 a_n2390_n5888# 0.012359f
C240 source.n129 a_n2390_n5888# 0.022999f
C241 source.n130 a_n2390_n5888# 0.022999f
C242 source.n131 a_n2390_n5888# 0.012359f
C243 source.n132 a_n2390_n5888# 0.013086f
C244 source.n133 a_n2390_n5888# 0.029211f
C245 source.n134 a_n2390_n5888# 0.06214f
C246 source.n135 a_n2390_n5888# 0.013086f
C247 source.n136 a_n2390_n5888# 0.012359f
C248 source.n137 a_n2390_n5888# 0.050647f
C249 source.n138 a_n2390_n5888# 0.034578f
C250 source.n139 a_n2390_n5888# 1.83721f
C251 source.t27 a_n2390_n5888# 0.454361f
C252 source.t28 a_n2390_n5888# 0.454361f
C253 source.n140 a_n2390_n5888# 4.11203f
C254 source.n141 a_n2390_n5888# 0.357372f
C255 source.t22 a_n2390_n5888# 0.454361f
C256 source.t24 a_n2390_n5888# 0.454361f
C257 source.n142 a_n2390_n5888# 4.11203f
C258 source.n143 a_n2390_n5888# 0.357372f
C259 source.t20 a_n2390_n5888# 0.454361f
C260 source.t21 a_n2390_n5888# 0.454361f
C261 source.n144 a_n2390_n5888# 4.11203f
C262 source.n145 a_n2390_n5888# 0.357372f
C263 source.n146 a_n2390_n5888# 0.031706f
C264 source.n147 a_n2390_n5888# 0.022999f
C265 source.n148 a_n2390_n5888# 0.012359f
C266 source.n149 a_n2390_n5888# 0.029211f
C267 source.n150 a_n2390_n5888# 0.013086f
C268 source.n151 a_n2390_n5888# 0.022999f
C269 source.n152 a_n2390_n5888# 0.012359f
C270 source.n153 a_n2390_n5888# 0.029211f
C271 source.n154 a_n2390_n5888# 0.013086f
C272 source.n155 a_n2390_n5888# 0.022999f
C273 source.n156 a_n2390_n5888# 0.012359f
C274 source.n157 a_n2390_n5888# 0.029211f
C275 source.n158 a_n2390_n5888# 0.013086f
C276 source.n159 a_n2390_n5888# 0.022999f
C277 source.n160 a_n2390_n5888# 0.012359f
C278 source.n161 a_n2390_n5888# 0.029211f
C279 source.n162 a_n2390_n5888# 0.029211f
C280 source.n163 a_n2390_n5888# 0.013086f
C281 source.n164 a_n2390_n5888# 0.022999f
C282 source.n165 a_n2390_n5888# 0.012359f
C283 source.n166 a_n2390_n5888# 0.029211f
C284 source.n167 a_n2390_n5888# 0.013086f
C285 source.n168 a_n2390_n5888# 0.022999f
C286 source.n169 a_n2390_n5888# 0.012359f
C287 source.n170 a_n2390_n5888# 0.029211f
C288 source.n171 a_n2390_n5888# 0.013086f
C289 source.n172 a_n2390_n5888# 0.022999f
C290 source.n173 a_n2390_n5888# 0.012359f
C291 source.n174 a_n2390_n5888# 0.029211f
C292 source.n175 a_n2390_n5888# 0.013086f
C293 source.n176 a_n2390_n5888# 0.022999f
C294 source.n177 a_n2390_n5888# 0.012359f
C295 source.n178 a_n2390_n5888# 0.029211f
C296 source.n179 a_n2390_n5888# 0.013086f
C297 source.n180 a_n2390_n5888# 0.022999f
C298 source.n181 a_n2390_n5888# 0.012722f
C299 source.n182 a_n2390_n5888# 0.029211f
C300 source.n183 a_n2390_n5888# 0.012359f
C301 source.n184 a_n2390_n5888# 0.013086f
C302 source.n185 a_n2390_n5888# 0.022999f
C303 source.n186 a_n2390_n5888# 0.012359f
C304 source.n187 a_n2390_n5888# 0.029211f
C305 source.n188 a_n2390_n5888# 0.013086f
C306 source.n189 a_n2390_n5888# 0.022999f
C307 source.n190 a_n2390_n5888# 0.012359f
C308 source.n191 a_n2390_n5888# 0.021909f
C309 source.n192 a_n2390_n5888# 0.02065f
C310 source.t19 a_n2390_n5888# 0.050946f
C311 source.n193 a_n2390_n5888# 0.280606f
C312 source.n194 a_n2390_n5888# 2.49011f
C313 source.n195 a_n2390_n5888# 0.012359f
C314 source.n196 a_n2390_n5888# 0.013086f
C315 source.n197 a_n2390_n5888# 0.029211f
C316 source.n198 a_n2390_n5888# 0.029211f
C317 source.n199 a_n2390_n5888# 0.013086f
C318 source.n200 a_n2390_n5888# 0.012359f
C319 source.n201 a_n2390_n5888# 0.022999f
C320 source.n202 a_n2390_n5888# 0.022999f
C321 source.n203 a_n2390_n5888# 0.012359f
C322 source.n204 a_n2390_n5888# 0.013086f
C323 source.n205 a_n2390_n5888# 0.029211f
C324 source.n206 a_n2390_n5888# 0.029211f
C325 source.n207 a_n2390_n5888# 0.013086f
C326 source.n208 a_n2390_n5888# 0.012359f
C327 source.n209 a_n2390_n5888# 0.022999f
C328 source.n210 a_n2390_n5888# 0.022999f
C329 source.n211 a_n2390_n5888# 0.012359f
C330 source.n212 a_n2390_n5888# 0.013086f
C331 source.n213 a_n2390_n5888# 0.029211f
C332 source.n214 a_n2390_n5888# 0.029211f
C333 source.n215 a_n2390_n5888# 0.029211f
C334 source.n216 a_n2390_n5888# 0.012722f
C335 source.n217 a_n2390_n5888# 0.012359f
C336 source.n218 a_n2390_n5888# 0.022999f
C337 source.n219 a_n2390_n5888# 0.022999f
C338 source.n220 a_n2390_n5888# 0.012359f
C339 source.n221 a_n2390_n5888# 0.013086f
C340 source.n222 a_n2390_n5888# 0.029211f
C341 source.n223 a_n2390_n5888# 0.029211f
C342 source.n224 a_n2390_n5888# 0.013086f
C343 source.n225 a_n2390_n5888# 0.012359f
C344 source.n226 a_n2390_n5888# 0.022999f
C345 source.n227 a_n2390_n5888# 0.022999f
C346 source.n228 a_n2390_n5888# 0.012359f
C347 source.n229 a_n2390_n5888# 0.013086f
C348 source.n230 a_n2390_n5888# 0.029211f
C349 source.n231 a_n2390_n5888# 0.029211f
C350 source.n232 a_n2390_n5888# 0.013086f
C351 source.n233 a_n2390_n5888# 0.012359f
C352 source.n234 a_n2390_n5888# 0.022999f
C353 source.n235 a_n2390_n5888# 0.022999f
C354 source.n236 a_n2390_n5888# 0.012359f
C355 source.n237 a_n2390_n5888# 0.013086f
C356 source.n238 a_n2390_n5888# 0.029211f
C357 source.n239 a_n2390_n5888# 0.029211f
C358 source.n240 a_n2390_n5888# 0.013086f
C359 source.n241 a_n2390_n5888# 0.012359f
C360 source.n242 a_n2390_n5888# 0.022999f
C361 source.n243 a_n2390_n5888# 0.022999f
C362 source.n244 a_n2390_n5888# 0.012359f
C363 source.n245 a_n2390_n5888# 0.013086f
C364 source.n246 a_n2390_n5888# 0.029211f
C365 source.n247 a_n2390_n5888# 0.029211f
C366 source.n248 a_n2390_n5888# 0.013086f
C367 source.n249 a_n2390_n5888# 0.012359f
C368 source.n250 a_n2390_n5888# 0.022999f
C369 source.n251 a_n2390_n5888# 0.022999f
C370 source.n252 a_n2390_n5888# 0.012359f
C371 source.n253 a_n2390_n5888# 0.013086f
C372 source.n254 a_n2390_n5888# 0.029211f
C373 source.n255 a_n2390_n5888# 0.029211f
C374 source.n256 a_n2390_n5888# 0.013086f
C375 source.n257 a_n2390_n5888# 0.012359f
C376 source.n258 a_n2390_n5888# 0.022999f
C377 source.n259 a_n2390_n5888# 0.022999f
C378 source.n260 a_n2390_n5888# 0.012359f
C379 source.n261 a_n2390_n5888# 0.012722f
C380 source.n262 a_n2390_n5888# 0.012722f
C381 source.n263 a_n2390_n5888# 0.029211f
C382 source.n264 a_n2390_n5888# 0.029211f
C383 source.n265 a_n2390_n5888# 0.013086f
C384 source.n266 a_n2390_n5888# 0.012359f
C385 source.n267 a_n2390_n5888# 0.022999f
C386 source.n268 a_n2390_n5888# 0.022999f
C387 source.n269 a_n2390_n5888# 0.012359f
C388 source.n270 a_n2390_n5888# 0.013086f
C389 source.n271 a_n2390_n5888# 0.029211f
C390 source.n272 a_n2390_n5888# 0.029211f
C391 source.n273 a_n2390_n5888# 0.013086f
C392 source.n274 a_n2390_n5888# 0.012359f
C393 source.n275 a_n2390_n5888# 0.022999f
C394 source.n276 a_n2390_n5888# 0.022999f
C395 source.n277 a_n2390_n5888# 0.012359f
C396 source.n278 a_n2390_n5888# 0.013086f
C397 source.n279 a_n2390_n5888# 0.029211f
C398 source.n280 a_n2390_n5888# 0.06214f
C399 source.n281 a_n2390_n5888# 0.013086f
C400 source.n282 a_n2390_n5888# 0.012359f
C401 source.n283 a_n2390_n5888# 0.050647f
C402 source.n284 a_n2390_n5888# 0.034578f
C403 source.n285 a_n2390_n5888# 0.112458f
C404 source.n286 a_n2390_n5888# 0.031706f
C405 source.n287 a_n2390_n5888# 0.022999f
C406 source.n288 a_n2390_n5888# 0.012359f
C407 source.n289 a_n2390_n5888# 0.029211f
C408 source.n290 a_n2390_n5888# 0.013086f
C409 source.n291 a_n2390_n5888# 0.022999f
C410 source.n292 a_n2390_n5888# 0.012359f
C411 source.n293 a_n2390_n5888# 0.029211f
C412 source.n294 a_n2390_n5888# 0.013086f
C413 source.n295 a_n2390_n5888# 0.022999f
C414 source.n296 a_n2390_n5888# 0.012359f
C415 source.n297 a_n2390_n5888# 0.029211f
C416 source.n298 a_n2390_n5888# 0.013086f
C417 source.n299 a_n2390_n5888# 0.022999f
C418 source.n300 a_n2390_n5888# 0.012359f
C419 source.n301 a_n2390_n5888# 0.029211f
C420 source.n302 a_n2390_n5888# 0.029211f
C421 source.n303 a_n2390_n5888# 0.013086f
C422 source.n304 a_n2390_n5888# 0.022999f
C423 source.n305 a_n2390_n5888# 0.012359f
C424 source.n306 a_n2390_n5888# 0.029211f
C425 source.n307 a_n2390_n5888# 0.013086f
C426 source.n308 a_n2390_n5888# 0.022999f
C427 source.n309 a_n2390_n5888# 0.012359f
C428 source.n310 a_n2390_n5888# 0.029211f
C429 source.n311 a_n2390_n5888# 0.013086f
C430 source.n312 a_n2390_n5888# 0.022999f
C431 source.n313 a_n2390_n5888# 0.012359f
C432 source.n314 a_n2390_n5888# 0.029211f
C433 source.n315 a_n2390_n5888# 0.013086f
C434 source.n316 a_n2390_n5888# 0.022999f
C435 source.n317 a_n2390_n5888# 0.012359f
C436 source.n318 a_n2390_n5888# 0.029211f
C437 source.n319 a_n2390_n5888# 0.013086f
C438 source.n320 a_n2390_n5888# 0.022999f
C439 source.n321 a_n2390_n5888# 0.012722f
C440 source.n322 a_n2390_n5888# 0.029211f
C441 source.n323 a_n2390_n5888# 0.012359f
C442 source.n324 a_n2390_n5888# 0.013086f
C443 source.n325 a_n2390_n5888# 0.022999f
C444 source.n326 a_n2390_n5888# 0.012359f
C445 source.n327 a_n2390_n5888# 0.029211f
C446 source.n328 a_n2390_n5888# 0.013086f
C447 source.n329 a_n2390_n5888# 0.022999f
C448 source.n330 a_n2390_n5888# 0.012359f
C449 source.n331 a_n2390_n5888# 0.021909f
C450 source.n332 a_n2390_n5888# 0.02065f
C451 source.t1 a_n2390_n5888# 0.050946f
C452 source.n333 a_n2390_n5888# 0.280606f
C453 source.n334 a_n2390_n5888# 2.49011f
C454 source.n335 a_n2390_n5888# 0.012359f
C455 source.n336 a_n2390_n5888# 0.013086f
C456 source.n337 a_n2390_n5888# 0.029211f
C457 source.n338 a_n2390_n5888# 0.029211f
C458 source.n339 a_n2390_n5888# 0.013086f
C459 source.n340 a_n2390_n5888# 0.012359f
C460 source.n341 a_n2390_n5888# 0.022999f
C461 source.n342 a_n2390_n5888# 0.022999f
C462 source.n343 a_n2390_n5888# 0.012359f
C463 source.n344 a_n2390_n5888# 0.013086f
C464 source.n345 a_n2390_n5888# 0.029211f
C465 source.n346 a_n2390_n5888# 0.029211f
C466 source.n347 a_n2390_n5888# 0.013086f
C467 source.n348 a_n2390_n5888# 0.012359f
C468 source.n349 a_n2390_n5888# 0.022999f
C469 source.n350 a_n2390_n5888# 0.022999f
C470 source.n351 a_n2390_n5888# 0.012359f
C471 source.n352 a_n2390_n5888# 0.013086f
C472 source.n353 a_n2390_n5888# 0.029211f
C473 source.n354 a_n2390_n5888# 0.029211f
C474 source.n355 a_n2390_n5888# 0.029211f
C475 source.n356 a_n2390_n5888# 0.012722f
C476 source.n357 a_n2390_n5888# 0.012359f
C477 source.n358 a_n2390_n5888# 0.022999f
C478 source.n359 a_n2390_n5888# 0.022999f
C479 source.n360 a_n2390_n5888# 0.012359f
C480 source.n361 a_n2390_n5888# 0.013086f
C481 source.n362 a_n2390_n5888# 0.029211f
C482 source.n363 a_n2390_n5888# 0.029211f
C483 source.n364 a_n2390_n5888# 0.013086f
C484 source.n365 a_n2390_n5888# 0.012359f
C485 source.n366 a_n2390_n5888# 0.022999f
C486 source.n367 a_n2390_n5888# 0.022999f
C487 source.n368 a_n2390_n5888# 0.012359f
C488 source.n369 a_n2390_n5888# 0.013086f
C489 source.n370 a_n2390_n5888# 0.029211f
C490 source.n371 a_n2390_n5888# 0.029211f
C491 source.n372 a_n2390_n5888# 0.013086f
C492 source.n373 a_n2390_n5888# 0.012359f
C493 source.n374 a_n2390_n5888# 0.022999f
C494 source.n375 a_n2390_n5888# 0.022999f
C495 source.n376 a_n2390_n5888# 0.012359f
C496 source.n377 a_n2390_n5888# 0.013086f
C497 source.n378 a_n2390_n5888# 0.029211f
C498 source.n379 a_n2390_n5888# 0.029211f
C499 source.n380 a_n2390_n5888# 0.013086f
C500 source.n381 a_n2390_n5888# 0.012359f
C501 source.n382 a_n2390_n5888# 0.022999f
C502 source.n383 a_n2390_n5888# 0.022999f
C503 source.n384 a_n2390_n5888# 0.012359f
C504 source.n385 a_n2390_n5888# 0.013086f
C505 source.n386 a_n2390_n5888# 0.029211f
C506 source.n387 a_n2390_n5888# 0.029211f
C507 source.n388 a_n2390_n5888# 0.013086f
C508 source.n389 a_n2390_n5888# 0.012359f
C509 source.n390 a_n2390_n5888# 0.022999f
C510 source.n391 a_n2390_n5888# 0.022999f
C511 source.n392 a_n2390_n5888# 0.012359f
C512 source.n393 a_n2390_n5888# 0.013086f
C513 source.n394 a_n2390_n5888# 0.029211f
C514 source.n395 a_n2390_n5888# 0.029211f
C515 source.n396 a_n2390_n5888# 0.013086f
C516 source.n397 a_n2390_n5888# 0.012359f
C517 source.n398 a_n2390_n5888# 0.022999f
C518 source.n399 a_n2390_n5888# 0.022999f
C519 source.n400 a_n2390_n5888# 0.012359f
C520 source.n401 a_n2390_n5888# 0.012722f
C521 source.n402 a_n2390_n5888# 0.012722f
C522 source.n403 a_n2390_n5888# 0.029211f
C523 source.n404 a_n2390_n5888# 0.029211f
C524 source.n405 a_n2390_n5888# 0.013086f
C525 source.n406 a_n2390_n5888# 0.012359f
C526 source.n407 a_n2390_n5888# 0.022999f
C527 source.n408 a_n2390_n5888# 0.022999f
C528 source.n409 a_n2390_n5888# 0.012359f
C529 source.n410 a_n2390_n5888# 0.013086f
C530 source.n411 a_n2390_n5888# 0.029211f
C531 source.n412 a_n2390_n5888# 0.029211f
C532 source.n413 a_n2390_n5888# 0.013086f
C533 source.n414 a_n2390_n5888# 0.012359f
C534 source.n415 a_n2390_n5888# 0.022999f
C535 source.n416 a_n2390_n5888# 0.022999f
C536 source.n417 a_n2390_n5888# 0.012359f
C537 source.n418 a_n2390_n5888# 0.013086f
C538 source.n419 a_n2390_n5888# 0.029211f
C539 source.n420 a_n2390_n5888# 0.06214f
C540 source.n421 a_n2390_n5888# 0.013086f
C541 source.n422 a_n2390_n5888# 0.012359f
C542 source.n423 a_n2390_n5888# 0.050647f
C543 source.n424 a_n2390_n5888# 0.034578f
C544 source.n425 a_n2390_n5888# 0.112458f
C545 source.t0 a_n2390_n5888# 0.454361f
C546 source.t12 a_n2390_n5888# 0.454361f
C547 source.n426 a_n2390_n5888# 4.11203f
C548 source.n427 a_n2390_n5888# 0.357372f
C549 source.t3 a_n2390_n5888# 0.454361f
C550 source.t11 a_n2390_n5888# 0.454361f
C551 source.n428 a_n2390_n5888# 4.11203f
C552 source.n429 a_n2390_n5888# 0.357372f
C553 source.t10 a_n2390_n5888# 0.454361f
C554 source.t4 a_n2390_n5888# 0.454361f
C555 source.n430 a_n2390_n5888# 4.11203f
C556 source.n431 a_n2390_n5888# 0.357372f
C557 source.n432 a_n2390_n5888# 0.031706f
C558 source.n433 a_n2390_n5888# 0.022999f
C559 source.n434 a_n2390_n5888# 0.012359f
C560 source.n435 a_n2390_n5888# 0.029211f
C561 source.n436 a_n2390_n5888# 0.013086f
C562 source.n437 a_n2390_n5888# 0.022999f
C563 source.n438 a_n2390_n5888# 0.012359f
C564 source.n439 a_n2390_n5888# 0.029211f
C565 source.n440 a_n2390_n5888# 0.013086f
C566 source.n441 a_n2390_n5888# 0.022999f
C567 source.n442 a_n2390_n5888# 0.012359f
C568 source.n443 a_n2390_n5888# 0.029211f
C569 source.n444 a_n2390_n5888# 0.013086f
C570 source.n445 a_n2390_n5888# 0.022999f
C571 source.n446 a_n2390_n5888# 0.012359f
C572 source.n447 a_n2390_n5888# 0.029211f
C573 source.n448 a_n2390_n5888# 0.029211f
C574 source.n449 a_n2390_n5888# 0.013086f
C575 source.n450 a_n2390_n5888# 0.022999f
C576 source.n451 a_n2390_n5888# 0.012359f
C577 source.n452 a_n2390_n5888# 0.029211f
C578 source.n453 a_n2390_n5888# 0.013086f
C579 source.n454 a_n2390_n5888# 0.022999f
C580 source.n455 a_n2390_n5888# 0.012359f
C581 source.n456 a_n2390_n5888# 0.029211f
C582 source.n457 a_n2390_n5888# 0.013086f
C583 source.n458 a_n2390_n5888# 0.022999f
C584 source.n459 a_n2390_n5888# 0.012359f
C585 source.n460 a_n2390_n5888# 0.029211f
C586 source.n461 a_n2390_n5888# 0.013086f
C587 source.n462 a_n2390_n5888# 0.022999f
C588 source.n463 a_n2390_n5888# 0.012359f
C589 source.n464 a_n2390_n5888# 0.029211f
C590 source.n465 a_n2390_n5888# 0.013086f
C591 source.n466 a_n2390_n5888# 0.022999f
C592 source.n467 a_n2390_n5888# 0.012722f
C593 source.n468 a_n2390_n5888# 0.029211f
C594 source.n469 a_n2390_n5888# 0.012359f
C595 source.n470 a_n2390_n5888# 0.013086f
C596 source.n471 a_n2390_n5888# 0.022999f
C597 source.n472 a_n2390_n5888# 0.012359f
C598 source.n473 a_n2390_n5888# 0.029211f
C599 source.n474 a_n2390_n5888# 0.013086f
C600 source.n475 a_n2390_n5888# 0.022999f
C601 source.n476 a_n2390_n5888# 0.012359f
C602 source.n477 a_n2390_n5888# 0.021909f
C603 source.n478 a_n2390_n5888# 0.02065f
C604 source.t6 a_n2390_n5888# 0.050946f
C605 source.n479 a_n2390_n5888# 0.280606f
C606 source.n480 a_n2390_n5888# 2.49011f
C607 source.n481 a_n2390_n5888# 0.012359f
C608 source.n482 a_n2390_n5888# 0.013086f
C609 source.n483 a_n2390_n5888# 0.029211f
C610 source.n484 a_n2390_n5888# 0.029211f
C611 source.n485 a_n2390_n5888# 0.013086f
C612 source.n486 a_n2390_n5888# 0.012359f
C613 source.n487 a_n2390_n5888# 0.022999f
C614 source.n488 a_n2390_n5888# 0.022999f
C615 source.n489 a_n2390_n5888# 0.012359f
C616 source.n490 a_n2390_n5888# 0.013086f
C617 source.n491 a_n2390_n5888# 0.029211f
C618 source.n492 a_n2390_n5888# 0.029211f
C619 source.n493 a_n2390_n5888# 0.013086f
C620 source.n494 a_n2390_n5888# 0.012359f
C621 source.n495 a_n2390_n5888# 0.022999f
C622 source.n496 a_n2390_n5888# 0.022999f
C623 source.n497 a_n2390_n5888# 0.012359f
C624 source.n498 a_n2390_n5888# 0.013086f
C625 source.n499 a_n2390_n5888# 0.029211f
C626 source.n500 a_n2390_n5888# 0.029211f
C627 source.n501 a_n2390_n5888# 0.029211f
C628 source.n502 a_n2390_n5888# 0.012722f
C629 source.n503 a_n2390_n5888# 0.012359f
C630 source.n504 a_n2390_n5888# 0.022999f
C631 source.n505 a_n2390_n5888# 0.022999f
C632 source.n506 a_n2390_n5888# 0.012359f
C633 source.n507 a_n2390_n5888# 0.013086f
C634 source.n508 a_n2390_n5888# 0.029211f
C635 source.n509 a_n2390_n5888# 0.029211f
C636 source.n510 a_n2390_n5888# 0.013086f
C637 source.n511 a_n2390_n5888# 0.012359f
C638 source.n512 a_n2390_n5888# 0.022999f
C639 source.n513 a_n2390_n5888# 0.022999f
C640 source.n514 a_n2390_n5888# 0.012359f
C641 source.n515 a_n2390_n5888# 0.013086f
C642 source.n516 a_n2390_n5888# 0.029211f
C643 source.n517 a_n2390_n5888# 0.029211f
C644 source.n518 a_n2390_n5888# 0.013086f
C645 source.n519 a_n2390_n5888# 0.012359f
C646 source.n520 a_n2390_n5888# 0.022999f
C647 source.n521 a_n2390_n5888# 0.022999f
C648 source.n522 a_n2390_n5888# 0.012359f
C649 source.n523 a_n2390_n5888# 0.013086f
C650 source.n524 a_n2390_n5888# 0.029211f
C651 source.n525 a_n2390_n5888# 0.029211f
C652 source.n526 a_n2390_n5888# 0.013086f
C653 source.n527 a_n2390_n5888# 0.012359f
C654 source.n528 a_n2390_n5888# 0.022999f
C655 source.n529 a_n2390_n5888# 0.022999f
C656 source.n530 a_n2390_n5888# 0.012359f
C657 source.n531 a_n2390_n5888# 0.013086f
C658 source.n532 a_n2390_n5888# 0.029211f
C659 source.n533 a_n2390_n5888# 0.029211f
C660 source.n534 a_n2390_n5888# 0.013086f
C661 source.n535 a_n2390_n5888# 0.012359f
C662 source.n536 a_n2390_n5888# 0.022999f
C663 source.n537 a_n2390_n5888# 0.022999f
C664 source.n538 a_n2390_n5888# 0.012359f
C665 source.n539 a_n2390_n5888# 0.013086f
C666 source.n540 a_n2390_n5888# 0.029211f
C667 source.n541 a_n2390_n5888# 0.029211f
C668 source.n542 a_n2390_n5888# 0.013086f
C669 source.n543 a_n2390_n5888# 0.012359f
C670 source.n544 a_n2390_n5888# 0.022999f
C671 source.n545 a_n2390_n5888# 0.022999f
C672 source.n546 a_n2390_n5888# 0.012359f
C673 source.n547 a_n2390_n5888# 0.012722f
C674 source.n548 a_n2390_n5888# 0.012722f
C675 source.n549 a_n2390_n5888# 0.029211f
C676 source.n550 a_n2390_n5888# 0.029211f
C677 source.n551 a_n2390_n5888# 0.013086f
C678 source.n552 a_n2390_n5888# 0.012359f
C679 source.n553 a_n2390_n5888# 0.022999f
C680 source.n554 a_n2390_n5888# 0.022999f
C681 source.n555 a_n2390_n5888# 0.012359f
C682 source.n556 a_n2390_n5888# 0.013086f
C683 source.n557 a_n2390_n5888# 0.029211f
C684 source.n558 a_n2390_n5888# 0.029211f
C685 source.n559 a_n2390_n5888# 0.013086f
C686 source.n560 a_n2390_n5888# 0.012359f
C687 source.n561 a_n2390_n5888# 0.022999f
C688 source.n562 a_n2390_n5888# 0.022999f
C689 source.n563 a_n2390_n5888# 0.012359f
C690 source.n564 a_n2390_n5888# 0.013086f
C691 source.n565 a_n2390_n5888# 0.029211f
C692 source.n566 a_n2390_n5888# 0.06214f
C693 source.n567 a_n2390_n5888# 0.013086f
C694 source.n568 a_n2390_n5888# 0.012359f
C695 source.n569 a_n2390_n5888# 0.050647f
C696 source.n570 a_n2390_n5888# 0.034578f
C697 source.n571 a_n2390_n5888# 2.27134f
C698 source.n572 a_n2390_n5888# 0.031706f
C699 source.n573 a_n2390_n5888# 0.022999f
C700 source.n574 a_n2390_n5888# 0.012359f
C701 source.n575 a_n2390_n5888# 0.029211f
C702 source.n576 a_n2390_n5888# 0.013086f
C703 source.n577 a_n2390_n5888# 0.022999f
C704 source.n578 a_n2390_n5888# 0.012359f
C705 source.n579 a_n2390_n5888# 0.029211f
C706 source.n580 a_n2390_n5888# 0.013086f
C707 source.n581 a_n2390_n5888# 0.022999f
C708 source.n582 a_n2390_n5888# 0.012359f
C709 source.n583 a_n2390_n5888# 0.029211f
C710 source.n584 a_n2390_n5888# 0.013086f
C711 source.n585 a_n2390_n5888# 0.022999f
C712 source.n586 a_n2390_n5888# 0.012359f
C713 source.n587 a_n2390_n5888# 0.029211f
C714 source.n588 a_n2390_n5888# 0.013086f
C715 source.n589 a_n2390_n5888# 0.022999f
C716 source.n590 a_n2390_n5888# 0.012359f
C717 source.n591 a_n2390_n5888# 0.029211f
C718 source.n592 a_n2390_n5888# 0.013086f
C719 source.n593 a_n2390_n5888# 0.022999f
C720 source.n594 a_n2390_n5888# 0.012359f
C721 source.n595 a_n2390_n5888# 0.029211f
C722 source.n596 a_n2390_n5888# 0.013086f
C723 source.n597 a_n2390_n5888# 0.022999f
C724 source.n598 a_n2390_n5888# 0.012359f
C725 source.n599 a_n2390_n5888# 0.029211f
C726 source.n600 a_n2390_n5888# 0.013086f
C727 source.n601 a_n2390_n5888# 0.022999f
C728 source.n602 a_n2390_n5888# 0.012359f
C729 source.n603 a_n2390_n5888# 0.029211f
C730 source.n604 a_n2390_n5888# 0.013086f
C731 source.n605 a_n2390_n5888# 0.022999f
C732 source.n606 a_n2390_n5888# 0.012722f
C733 source.n607 a_n2390_n5888# 0.029211f
C734 source.n608 a_n2390_n5888# 0.013086f
C735 source.n609 a_n2390_n5888# 0.022999f
C736 source.n610 a_n2390_n5888# 0.012359f
C737 source.n611 a_n2390_n5888# 0.029211f
C738 source.n612 a_n2390_n5888# 0.013086f
C739 source.n613 a_n2390_n5888# 0.022999f
C740 source.n614 a_n2390_n5888# 0.012359f
C741 source.n615 a_n2390_n5888# 0.021909f
C742 source.n616 a_n2390_n5888# 0.02065f
C743 source.t30 a_n2390_n5888# 0.050946f
C744 source.n617 a_n2390_n5888# 0.280606f
C745 source.n618 a_n2390_n5888# 2.49011f
C746 source.n619 a_n2390_n5888# 0.012359f
C747 source.n620 a_n2390_n5888# 0.013086f
C748 source.n621 a_n2390_n5888# 0.029211f
C749 source.n622 a_n2390_n5888# 0.029211f
C750 source.n623 a_n2390_n5888# 0.013086f
C751 source.n624 a_n2390_n5888# 0.012359f
C752 source.n625 a_n2390_n5888# 0.022999f
C753 source.n626 a_n2390_n5888# 0.022999f
C754 source.n627 a_n2390_n5888# 0.012359f
C755 source.n628 a_n2390_n5888# 0.013086f
C756 source.n629 a_n2390_n5888# 0.029211f
C757 source.n630 a_n2390_n5888# 0.029211f
C758 source.n631 a_n2390_n5888# 0.013086f
C759 source.n632 a_n2390_n5888# 0.012359f
C760 source.n633 a_n2390_n5888# 0.022999f
C761 source.n634 a_n2390_n5888# 0.022999f
C762 source.n635 a_n2390_n5888# 0.012359f
C763 source.n636 a_n2390_n5888# 0.012359f
C764 source.n637 a_n2390_n5888# 0.013086f
C765 source.n638 a_n2390_n5888# 0.029211f
C766 source.n639 a_n2390_n5888# 0.029211f
C767 source.n640 a_n2390_n5888# 0.029211f
C768 source.n641 a_n2390_n5888# 0.012722f
C769 source.n642 a_n2390_n5888# 0.012359f
C770 source.n643 a_n2390_n5888# 0.022999f
C771 source.n644 a_n2390_n5888# 0.022999f
C772 source.n645 a_n2390_n5888# 0.012359f
C773 source.n646 a_n2390_n5888# 0.013086f
C774 source.n647 a_n2390_n5888# 0.029211f
C775 source.n648 a_n2390_n5888# 0.029211f
C776 source.n649 a_n2390_n5888# 0.013086f
C777 source.n650 a_n2390_n5888# 0.012359f
C778 source.n651 a_n2390_n5888# 0.022999f
C779 source.n652 a_n2390_n5888# 0.022999f
C780 source.n653 a_n2390_n5888# 0.012359f
C781 source.n654 a_n2390_n5888# 0.013086f
C782 source.n655 a_n2390_n5888# 0.029211f
C783 source.n656 a_n2390_n5888# 0.029211f
C784 source.n657 a_n2390_n5888# 0.013086f
C785 source.n658 a_n2390_n5888# 0.012359f
C786 source.n659 a_n2390_n5888# 0.022999f
C787 source.n660 a_n2390_n5888# 0.022999f
C788 source.n661 a_n2390_n5888# 0.012359f
C789 source.n662 a_n2390_n5888# 0.013086f
C790 source.n663 a_n2390_n5888# 0.029211f
C791 source.n664 a_n2390_n5888# 0.029211f
C792 source.n665 a_n2390_n5888# 0.013086f
C793 source.n666 a_n2390_n5888# 0.012359f
C794 source.n667 a_n2390_n5888# 0.022999f
C795 source.n668 a_n2390_n5888# 0.022999f
C796 source.n669 a_n2390_n5888# 0.012359f
C797 source.n670 a_n2390_n5888# 0.013086f
C798 source.n671 a_n2390_n5888# 0.029211f
C799 source.n672 a_n2390_n5888# 0.029211f
C800 source.n673 a_n2390_n5888# 0.013086f
C801 source.n674 a_n2390_n5888# 0.012359f
C802 source.n675 a_n2390_n5888# 0.022999f
C803 source.n676 a_n2390_n5888# 0.022999f
C804 source.n677 a_n2390_n5888# 0.012359f
C805 source.n678 a_n2390_n5888# 0.013086f
C806 source.n679 a_n2390_n5888# 0.029211f
C807 source.n680 a_n2390_n5888# 0.029211f
C808 source.n681 a_n2390_n5888# 0.029211f
C809 source.n682 a_n2390_n5888# 0.013086f
C810 source.n683 a_n2390_n5888# 0.012359f
C811 source.n684 a_n2390_n5888# 0.022999f
C812 source.n685 a_n2390_n5888# 0.022999f
C813 source.n686 a_n2390_n5888# 0.012359f
C814 source.n687 a_n2390_n5888# 0.012722f
C815 source.n688 a_n2390_n5888# 0.012722f
C816 source.n689 a_n2390_n5888# 0.029211f
C817 source.n690 a_n2390_n5888# 0.029211f
C818 source.n691 a_n2390_n5888# 0.013086f
C819 source.n692 a_n2390_n5888# 0.012359f
C820 source.n693 a_n2390_n5888# 0.022999f
C821 source.n694 a_n2390_n5888# 0.022999f
C822 source.n695 a_n2390_n5888# 0.012359f
C823 source.n696 a_n2390_n5888# 0.013086f
C824 source.n697 a_n2390_n5888# 0.029211f
C825 source.n698 a_n2390_n5888# 0.029211f
C826 source.n699 a_n2390_n5888# 0.013086f
C827 source.n700 a_n2390_n5888# 0.012359f
C828 source.n701 a_n2390_n5888# 0.022999f
C829 source.n702 a_n2390_n5888# 0.022999f
C830 source.n703 a_n2390_n5888# 0.012359f
C831 source.n704 a_n2390_n5888# 0.013086f
C832 source.n705 a_n2390_n5888# 0.029211f
C833 source.n706 a_n2390_n5888# 0.06214f
C834 source.n707 a_n2390_n5888# 0.013086f
C835 source.n708 a_n2390_n5888# 0.012359f
C836 source.n709 a_n2390_n5888# 0.050647f
C837 source.n710 a_n2390_n5888# 0.034578f
C838 source.n711 a_n2390_n5888# 2.27134f
C839 source.t17 a_n2390_n5888# 0.454361f
C840 source.t25 a_n2390_n5888# 0.454361f
C841 source.n712 a_n2390_n5888# 4.11203f
C842 source.n713 a_n2390_n5888# 0.357374f
C843 source.t26 a_n2390_n5888# 0.454361f
C844 source.t31 a_n2390_n5888# 0.454361f
C845 source.n714 a_n2390_n5888# 4.11203f
C846 source.n715 a_n2390_n5888# 0.357374f
C847 source.t18 a_n2390_n5888# 0.454361f
C848 source.t23 a_n2390_n5888# 0.454361f
C849 source.n716 a_n2390_n5888# 4.11203f
C850 source.n717 a_n2390_n5888# 0.357374f
C851 source.n718 a_n2390_n5888# 0.031706f
C852 source.n719 a_n2390_n5888# 0.022999f
C853 source.n720 a_n2390_n5888# 0.012359f
C854 source.n721 a_n2390_n5888# 0.029211f
C855 source.n722 a_n2390_n5888# 0.013086f
C856 source.n723 a_n2390_n5888# 0.022999f
C857 source.n724 a_n2390_n5888# 0.012359f
C858 source.n725 a_n2390_n5888# 0.029211f
C859 source.n726 a_n2390_n5888# 0.013086f
C860 source.n727 a_n2390_n5888# 0.022999f
C861 source.n728 a_n2390_n5888# 0.012359f
C862 source.n729 a_n2390_n5888# 0.029211f
C863 source.n730 a_n2390_n5888# 0.013086f
C864 source.n731 a_n2390_n5888# 0.022999f
C865 source.n732 a_n2390_n5888# 0.012359f
C866 source.n733 a_n2390_n5888# 0.029211f
C867 source.n734 a_n2390_n5888# 0.013086f
C868 source.n735 a_n2390_n5888# 0.022999f
C869 source.n736 a_n2390_n5888# 0.012359f
C870 source.n737 a_n2390_n5888# 0.029211f
C871 source.n738 a_n2390_n5888# 0.013086f
C872 source.n739 a_n2390_n5888# 0.022999f
C873 source.n740 a_n2390_n5888# 0.012359f
C874 source.n741 a_n2390_n5888# 0.029211f
C875 source.n742 a_n2390_n5888# 0.013086f
C876 source.n743 a_n2390_n5888# 0.022999f
C877 source.n744 a_n2390_n5888# 0.012359f
C878 source.n745 a_n2390_n5888# 0.029211f
C879 source.n746 a_n2390_n5888# 0.013086f
C880 source.n747 a_n2390_n5888# 0.022999f
C881 source.n748 a_n2390_n5888# 0.012359f
C882 source.n749 a_n2390_n5888# 0.029211f
C883 source.n750 a_n2390_n5888# 0.013086f
C884 source.n751 a_n2390_n5888# 0.022999f
C885 source.n752 a_n2390_n5888# 0.012722f
C886 source.n753 a_n2390_n5888# 0.029211f
C887 source.n754 a_n2390_n5888# 0.013086f
C888 source.n755 a_n2390_n5888# 0.022999f
C889 source.n756 a_n2390_n5888# 0.012359f
C890 source.n757 a_n2390_n5888# 0.029211f
C891 source.n758 a_n2390_n5888# 0.013086f
C892 source.n759 a_n2390_n5888# 0.022999f
C893 source.n760 a_n2390_n5888# 0.012359f
C894 source.n761 a_n2390_n5888# 0.021909f
C895 source.n762 a_n2390_n5888# 0.02065f
C896 source.t16 a_n2390_n5888# 0.050946f
C897 source.n763 a_n2390_n5888# 0.280606f
C898 source.n764 a_n2390_n5888# 2.49011f
C899 source.n765 a_n2390_n5888# 0.012359f
C900 source.n766 a_n2390_n5888# 0.013086f
C901 source.n767 a_n2390_n5888# 0.029211f
C902 source.n768 a_n2390_n5888# 0.029211f
C903 source.n769 a_n2390_n5888# 0.013086f
C904 source.n770 a_n2390_n5888# 0.012359f
C905 source.n771 a_n2390_n5888# 0.022999f
C906 source.n772 a_n2390_n5888# 0.022999f
C907 source.n773 a_n2390_n5888# 0.012359f
C908 source.n774 a_n2390_n5888# 0.013086f
C909 source.n775 a_n2390_n5888# 0.029211f
C910 source.n776 a_n2390_n5888# 0.029211f
C911 source.n777 a_n2390_n5888# 0.013086f
C912 source.n778 a_n2390_n5888# 0.012359f
C913 source.n779 a_n2390_n5888# 0.022999f
C914 source.n780 a_n2390_n5888# 0.022999f
C915 source.n781 a_n2390_n5888# 0.012359f
C916 source.n782 a_n2390_n5888# 0.012359f
C917 source.n783 a_n2390_n5888# 0.013086f
C918 source.n784 a_n2390_n5888# 0.029211f
C919 source.n785 a_n2390_n5888# 0.029211f
C920 source.n786 a_n2390_n5888# 0.029211f
C921 source.n787 a_n2390_n5888# 0.012722f
C922 source.n788 a_n2390_n5888# 0.012359f
C923 source.n789 a_n2390_n5888# 0.022999f
C924 source.n790 a_n2390_n5888# 0.022999f
C925 source.n791 a_n2390_n5888# 0.012359f
C926 source.n792 a_n2390_n5888# 0.013086f
C927 source.n793 a_n2390_n5888# 0.029211f
C928 source.n794 a_n2390_n5888# 0.029211f
C929 source.n795 a_n2390_n5888# 0.013086f
C930 source.n796 a_n2390_n5888# 0.012359f
C931 source.n797 a_n2390_n5888# 0.022999f
C932 source.n798 a_n2390_n5888# 0.022999f
C933 source.n799 a_n2390_n5888# 0.012359f
C934 source.n800 a_n2390_n5888# 0.013086f
C935 source.n801 a_n2390_n5888# 0.029211f
C936 source.n802 a_n2390_n5888# 0.029211f
C937 source.n803 a_n2390_n5888# 0.013086f
C938 source.n804 a_n2390_n5888# 0.012359f
C939 source.n805 a_n2390_n5888# 0.022999f
C940 source.n806 a_n2390_n5888# 0.022999f
C941 source.n807 a_n2390_n5888# 0.012359f
C942 source.n808 a_n2390_n5888# 0.013086f
C943 source.n809 a_n2390_n5888# 0.029211f
C944 source.n810 a_n2390_n5888# 0.029211f
C945 source.n811 a_n2390_n5888# 0.013086f
C946 source.n812 a_n2390_n5888# 0.012359f
C947 source.n813 a_n2390_n5888# 0.022999f
C948 source.n814 a_n2390_n5888# 0.022999f
C949 source.n815 a_n2390_n5888# 0.012359f
C950 source.n816 a_n2390_n5888# 0.013086f
C951 source.n817 a_n2390_n5888# 0.029211f
C952 source.n818 a_n2390_n5888# 0.029211f
C953 source.n819 a_n2390_n5888# 0.013086f
C954 source.n820 a_n2390_n5888# 0.012359f
C955 source.n821 a_n2390_n5888# 0.022999f
C956 source.n822 a_n2390_n5888# 0.022999f
C957 source.n823 a_n2390_n5888# 0.012359f
C958 source.n824 a_n2390_n5888# 0.013086f
C959 source.n825 a_n2390_n5888# 0.029211f
C960 source.n826 a_n2390_n5888# 0.029211f
C961 source.n827 a_n2390_n5888# 0.029211f
C962 source.n828 a_n2390_n5888# 0.013086f
C963 source.n829 a_n2390_n5888# 0.012359f
C964 source.n830 a_n2390_n5888# 0.022999f
C965 source.n831 a_n2390_n5888# 0.022999f
C966 source.n832 a_n2390_n5888# 0.012359f
C967 source.n833 a_n2390_n5888# 0.012722f
C968 source.n834 a_n2390_n5888# 0.012722f
C969 source.n835 a_n2390_n5888# 0.029211f
C970 source.n836 a_n2390_n5888# 0.029211f
C971 source.n837 a_n2390_n5888# 0.013086f
C972 source.n838 a_n2390_n5888# 0.012359f
C973 source.n839 a_n2390_n5888# 0.022999f
C974 source.n840 a_n2390_n5888# 0.022999f
C975 source.n841 a_n2390_n5888# 0.012359f
C976 source.n842 a_n2390_n5888# 0.013086f
C977 source.n843 a_n2390_n5888# 0.029211f
C978 source.n844 a_n2390_n5888# 0.029211f
C979 source.n845 a_n2390_n5888# 0.013086f
C980 source.n846 a_n2390_n5888# 0.012359f
C981 source.n847 a_n2390_n5888# 0.022999f
C982 source.n848 a_n2390_n5888# 0.022999f
C983 source.n849 a_n2390_n5888# 0.012359f
C984 source.n850 a_n2390_n5888# 0.013086f
C985 source.n851 a_n2390_n5888# 0.029211f
C986 source.n852 a_n2390_n5888# 0.06214f
C987 source.n853 a_n2390_n5888# 0.013086f
C988 source.n854 a_n2390_n5888# 0.012359f
C989 source.n855 a_n2390_n5888# 0.050647f
C990 source.n856 a_n2390_n5888# 0.034578f
C991 source.n857 a_n2390_n5888# 0.112458f
C992 source.n858 a_n2390_n5888# 0.031706f
C993 source.n859 a_n2390_n5888# 0.022999f
C994 source.n860 a_n2390_n5888# 0.012359f
C995 source.n861 a_n2390_n5888# 0.029211f
C996 source.n862 a_n2390_n5888# 0.013086f
C997 source.n863 a_n2390_n5888# 0.022999f
C998 source.n864 a_n2390_n5888# 0.012359f
C999 source.n865 a_n2390_n5888# 0.029211f
C1000 source.n866 a_n2390_n5888# 0.013086f
C1001 source.n867 a_n2390_n5888# 0.022999f
C1002 source.n868 a_n2390_n5888# 0.012359f
C1003 source.n869 a_n2390_n5888# 0.029211f
C1004 source.n870 a_n2390_n5888# 0.013086f
C1005 source.n871 a_n2390_n5888# 0.022999f
C1006 source.n872 a_n2390_n5888# 0.012359f
C1007 source.n873 a_n2390_n5888# 0.029211f
C1008 source.n874 a_n2390_n5888# 0.013086f
C1009 source.n875 a_n2390_n5888# 0.022999f
C1010 source.n876 a_n2390_n5888# 0.012359f
C1011 source.n877 a_n2390_n5888# 0.029211f
C1012 source.n878 a_n2390_n5888# 0.013086f
C1013 source.n879 a_n2390_n5888# 0.022999f
C1014 source.n880 a_n2390_n5888# 0.012359f
C1015 source.n881 a_n2390_n5888# 0.029211f
C1016 source.n882 a_n2390_n5888# 0.013086f
C1017 source.n883 a_n2390_n5888# 0.022999f
C1018 source.n884 a_n2390_n5888# 0.012359f
C1019 source.n885 a_n2390_n5888# 0.029211f
C1020 source.n886 a_n2390_n5888# 0.013086f
C1021 source.n887 a_n2390_n5888# 0.022999f
C1022 source.n888 a_n2390_n5888# 0.012359f
C1023 source.n889 a_n2390_n5888# 0.029211f
C1024 source.n890 a_n2390_n5888# 0.013086f
C1025 source.n891 a_n2390_n5888# 0.022999f
C1026 source.n892 a_n2390_n5888# 0.012722f
C1027 source.n893 a_n2390_n5888# 0.029211f
C1028 source.n894 a_n2390_n5888# 0.013086f
C1029 source.n895 a_n2390_n5888# 0.022999f
C1030 source.n896 a_n2390_n5888# 0.012359f
C1031 source.n897 a_n2390_n5888# 0.029211f
C1032 source.n898 a_n2390_n5888# 0.013086f
C1033 source.n899 a_n2390_n5888# 0.022999f
C1034 source.n900 a_n2390_n5888# 0.012359f
C1035 source.n901 a_n2390_n5888# 0.021909f
C1036 source.n902 a_n2390_n5888# 0.02065f
C1037 source.t2 a_n2390_n5888# 0.050946f
C1038 source.n903 a_n2390_n5888# 0.280606f
C1039 source.n904 a_n2390_n5888# 2.49011f
C1040 source.n905 a_n2390_n5888# 0.012359f
C1041 source.n906 a_n2390_n5888# 0.013086f
C1042 source.n907 a_n2390_n5888# 0.029211f
C1043 source.n908 a_n2390_n5888# 0.029211f
C1044 source.n909 a_n2390_n5888# 0.013086f
C1045 source.n910 a_n2390_n5888# 0.012359f
C1046 source.n911 a_n2390_n5888# 0.022999f
C1047 source.n912 a_n2390_n5888# 0.022999f
C1048 source.n913 a_n2390_n5888# 0.012359f
C1049 source.n914 a_n2390_n5888# 0.013086f
C1050 source.n915 a_n2390_n5888# 0.029211f
C1051 source.n916 a_n2390_n5888# 0.029211f
C1052 source.n917 a_n2390_n5888# 0.013086f
C1053 source.n918 a_n2390_n5888# 0.012359f
C1054 source.n919 a_n2390_n5888# 0.022999f
C1055 source.n920 a_n2390_n5888# 0.022999f
C1056 source.n921 a_n2390_n5888# 0.012359f
C1057 source.n922 a_n2390_n5888# 0.012359f
C1058 source.n923 a_n2390_n5888# 0.013086f
C1059 source.n924 a_n2390_n5888# 0.029211f
C1060 source.n925 a_n2390_n5888# 0.029211f
C1061 source.n926 a_n2390_n5888# 0.029211f
C1062 source.n927 a_n2390_n5888# 0.012722f
C1063 source.n928 a_n2390_n5888# 0.012359f
C1064 source.n929 a_n2390_n5888# 0.022999f
C1065 source.n930 a_n2390_n5888# 0.022999f
C1066 source.n931 a_n2390_n5888# 0.012359f
C1067 source.n932 a_n2390_n5888# 0.013086f
C1068 source.n933 a_n2390_n5888# 0.029211f
C1069 source.n934 a_n2390_n5888# 0.029211f
C1070 source.n935 a_n2390_n5888# 0.013086f
C1071 source.n936 a_n2390_n5888# 0.012359f
C1072 source.n937 a_n2390_n5888# 0.022999f
C1073 source.n938 a_n2390_n5888# 0.022999f
C1074 source.n939 a_n2390_n5888# 0.012359f
C1075 source.n940 a_n2390_n5888# 0.013086f
C1076 source.n941 a_n2390_n5888# 0.029211f
C1077 source.n942 a_n2390_n5888# 0.029211f
C1078 source.n943 a_n2390_n5888# 0.013086f
C1079 source.n944 a_n2390_n5888# 0.012359f
C1080 source.n945 a_n2390_n5888# 0.022999f
C1081 source.n946 a_n2390_n5888# 0.022999f
C1082 source.n947 a_n2390_n5888# 0.012359f
C1083 source.n948 a_n2390_n5888# 0.013086f
C1084 source.n949 a_n2390_n5888# 0.029211f
C1085 source.n950 a_n2390_n5888# 0.029211f
C1086 source.n951 a_n2390_n5888# 0.013086f
C1087 source.n952 a_n2390_n5888# 0.012359f
C1088 source.n953 a_n2390_n5888# 0.022999f
C1089 source.n954 a_n2390_n5888# 0.022999f
C1090 source.n955 a_n2390_n5888# 0.012359f
C1091 source.n956 a_n2390_n5888# 0.013086f
C1092 source.n957 a_n2390_n5888# 0.029211f
C1093 source.n958 a_n2390_n5888# 0.029211f
C1094 source.n959 a_n2390_n5888# 0.013086f
C1095 source.n960 a_n2390_n5888# 0.012359f
C1096 source.n961 a_n2390_n5888# 0.022999f
C1097 source.n962 a_n2390_n5888# 0.022999f
C1098 source.n963 a_n2390_n5888# 0.012359f
C1099 source.n964 a_n2390_n5888# 0.013086f
C1100 source.n965 a_n2390_n5888# 0.029211f
C1101 source.n966 a_n2390_n5888# 0.029211f
C1102 source.n967 a_n2390_n5888# 0.029211f
C1103 source.n968 a_n2390_n5888# 0.013086f
C1104 source.n969 a_n2390_n5888# 0.012359f
C1105 source.n970 a_n2390_n5888# 0.022999f
C1106 source.n971 a_n2390_n5888# 0.022999f
C1107 source.n972 a_n2390_n5888# 0.012359f
C1108 source.n973 a_n2390_n5888# 0.012722f
C1109 source.n974 a_n2390_n5888# 0.012722f
C1110 source.n975 a_n2390_n5888# 0.029211f
C1111 source.n976 a_n2390_n5888# 0.029211f
C1112 source.n977 a_n2390_n5888# 0.013086f
C1113 source.n978 a_n2390_n5888# 0.012359f
C1114 source.n979 a_n2390_n5888# 0.022999f
C1115 source.n980 a_n2390_n5888# 0.022999f
C1116 source.n981 a_n2390_n5888# 0.012359f
C1117 source.n982 a_n2390_n5888# 0.013086f
C1118 source.n983 a_n2390_n5888# 0.029211f
C1119 source.n984 a_n2390_n5888# 0.029211f
C1120 source.n985 a_n2390_n5888# 0.013086f
C1121 source.n986 a_n2390_n5888# 0.012359f
C1122 source.n987 a_n2390_n5888# 0.022999f
C1123 source.n988 a_n2390_n5888# 0.022999f
C1124 source.n989 a_n2390_n5888# 0.012359f
C1125 source.n990 a_n2390_n5888# 0.013086f
C1126 source.n991 a_n2390_n5888# 0.029211f
C1127 source.n992 a_n2390_n5888# 0.06214f
C1128 source.n993 a_n2390_n5888# 0.013086f
C1129 source.n994 a_n2390_n5888# 0.012359f
C1130 source.n995 a_n2390_n5888# 0.050647f
C1131 source.n996 a_n2390_n5888# 0.034578f
C1132 source.n997 a_n2390_n5888# 0.112458f
C1133 source.t15 a_n2390_n5888# 0.454361f
C1134 source.t8 a_n2390_n5888# 0.454361f
C1135 source.n998 a_n2390_n5888# 4.11203f
C1136 source.n999 a_n2390_n5888# 0.357374f
C1137 source.t5 a_n2390_n5888# 0.454361f
C1138 source.t14 a_n2390_n5888# 0.454361f
C1139 source.n1000 a_n2390_n5888# 4.11203f
C1140 source.n1001 a_n2390_n5888# 0.357374f
C1141 source.t9 a_n2390_n5888# 0.454361f
C1142 source.t7 a_n2390_n5888# 0.454361f
C1143 source.n1002 a_n2390_n5888# 4.11203f
C1144 source.n1003 a_n2390_n5888# 0.357374f
C1145 source.n1004 a_n2390_n5888# 0.031706f
C1146 source.n1005 a_n2390_n5888# 0.022999f
C1147 source.n1006 a_n2390_n5888# 0.012359f
C1148 source.n1007 a_n2390_n5888# 0.029211f
C1149 source.n1008 a_n2390_n5888# 0.013086f
C1150 source.n1009 a_n2390_n5888# 0.022999f
C1151 source.n1010 a_n2390_n5888# 0.012359f
C1152 source.n1011 a_n2390_n5888# 0.029211f
C1153 source.n1012 a_n2390_n5888# 0.013086f
C1154 source.n1013 a_n2390_n5888# 0.022999f
C1155 source.n1014 a_n2390_n5888# 0.012359f
C1156 source.n1015 a_n2390_n5888# 0.029211f
C1157 source.n1016 a_n2390_n5888# 0.013086f
C1158 source.n1017 a_n2390_n5888# 0.022999f
C1159 source.n1018 a_n2390_n5888# 0.012359f
C1160 source.n1019 a_n2390_n5888# 0.029211f
C1161 source.n1020 a_n2390_n5888# 0.013086f
C1162 source.n1021 a_n2390_n5888# 0.022999f
C1163 source.n1022 a_n2390_n5888# 0.012359f
C1164 source.n1023 a_n2390_n5888# 0.029211f
C1165 source.n1024 a_n2390_n5888# 0.013086f
C1166 source.n1025 a_n2390_n5888# 0.022999f
C1167 source.n1026 a_n2390_n5888# 0.012359f
C1168 source.n1027 a_n2390_n5888# 0.029211f
C1169 source.n1028 a_n2390_n5888# 0.013086f
C1170 source.n1029 a_n2390_n5888# 0.022999f
C1171 source.n1030 a_n2390_n5888# 0.012359f
C1172 source.n1031 a_n2390_n5888# 0.029211f
C1173 source.n1032 a_n2390_n5888# 0.013086f
C1174 source.n1033 a_n2390_n5888# 0.022999f
C1175 source.n1034 a_n2390_n5888# 0.012359f
C1176 source.n1035 a_n2390_n5888# 0.029211f
C1177 source.n1036 a_n2390_n5888# 0.013086f
C1178 source.n1037 a_n2390_n5888# 0.022999f
C1179 source.n1038 a_n2390_n5888# 0.012722f
C1180 source.n1039 a_n2390_n5888# 0.029211f
C1181 source.n1040 a_n2390_n5888# 0.013086f
C1182 source.n1041 a_n2390_n5888# 0.022999f
C1183 source.n1042 a_n2390_n5888# 0.012359f
C1184 source.n1043 a_n2390_n5888# 0.029211f
C1185 source.n1044 a_n2390_n5888# 0.013086f
C1186 source.n1045 a_n2390_n5888# 0.022999f
C1187 source.n1046 a_n2390_n5888# 0.012359f
C1188 source.n1047 a_n2390_n5888# 0.021909f
C1189 source.n1048 a_n2390_n5888# 0.02065f
C1190 source.t13 a_n2390_n5888# 0.050946f
C1191 source.n1049 a_n2390_n5888# 0.280606f
C1192 source.n1050 a_n2390_n5888# 2.49011f
C1193 source.n1051 a_n2390_n5888# 0.012359f
C1194 source.n1052 a_n2390_n5888# 0.013086f
C1195 source.n1053 a_n2390_n5888# 0.029211f
C1196 source.n1054 a_n2390_n5888# 0.029211f
C1197 source.n1055 a_n2390_n5888# 0.013086f
C1198 source.n1056 a_n2390_n5888# 0.012359f
C1199 source.n1057 a_n2390_n5888# 0.022999f
C1200 source.n1058 a_n2390_n5888# 0.022999f
C1201 source.n1059 a_n2390_n5888# 0.012359f
C1202 source.n1060 a_n2390_n5888# 0.013086f
C1203 source.n1061 a_n2390_n5888# 0.029211f
C1204 source.n1062 a_n2390_n5888# 0.029211f
C1205 source.n1063 a_n2390_n5888# 0.013086f
C1206 source.n1064 a_n2390_n5888# 0.012359f
C1207 source.n1065 a_n2390_n5888# 0.022999f
C1208 source.n1066 a_n2390_n5888# 0.022999f
C1209 source.n1067 a_n2390_n5888# 0.012359f
C1210 source.n1068 a_n2390_n5888# 0.012359f
C1211 source.n1069 a_n2390_n5888# 0.013086f
C1212 source.n1070 a_n2390_n5888# 0.029211f
C1213 source.n1071 a_n2390_n5888# 0.029211f
C1214 source.n1072 a_n2390_n5888# 0.029211f
C1215 source.n1073 a_n2390_n5888# 0.012722f
C1216 source.n1074 a_n2390_n5888# 0.012359f
C1217 source.n1075 a_n2390_n5888# 0.022999f
C1218 source.n1076 a_n2390_n5888# 0.022999f
C1219 source.n1077 a_n2390_n5888# 0.012359f
C1220 source.n1078 a_n2390_n5888# 0.013086f
C1221 source.n1079 a_n2390_n5888# 0.029211f
C1222 source.n1080 a_n2390_n5888# 0.029211f
C1223 source.n1081 a_n2390_n5888# 0.013086f
C1224 source.n1082 a_n2390_n5888# 0.012359f
C1225 source.n1083 a_n2390_n5888# 0.022999f
C1226 source.n1084 a_n2390_n5888# 0.022999f
C1227 source.n1085 a_n2390_n5888# 0.012359f
C1228 source.n1086 a_n2390_n5888# 0.013086f
C1229 source.n1087 a_n2390_n5888# 0.029211f
C1230 source.n1088 a_n2390_n5888# 0.029211f
C1231 source.n1089 a_n2390_n5888# 0.013086f
C1232 source.n1090 a_n2390_n5888# 0.012359f
C1233 source.n1091 a_n2390_n5888# 0.022999f
C1234 source.n1092 a_n2390_n5888# 0.022999f
C1235 source.n1093 a_n2390_n5888# 0.012359f
C1236 source.n1094 a_n2390_n5888# 0.013086f
C1237 source.n1095 a_n2390_n5888# 0.029211f
C1238 source.n1096 a_n2390_n5888# 0.029211f
C1239 source.n1097 a_n2390_n5888# 0.013086f
C1240 source.n1098 a_n2390_n5888# 0.012359f
C1241 source.n1099 a_n2390_n5888# 0.022999f
C1242 source.n1100 a_n2390_n5888# 0.022999f
C1243 source.n1101 a_n2390_n5888# 0.012359f
C1244 source.n1102 a_n2390_n5888# 0.013086f
C1245 source.n1103 a_n2390_n5888# 0.029211f
C1246 source.n1104 a_n2390_n5888# 0.029211f
C1247 source.n1105 a_n2390_n5888# 0.013086f
C1248 source.n1106 a_n2390_n5888# 0.012359f
C1249 source.n1107 a_n2390_n5888# 0.022999f
C1250 source.n1108 a_n2390_n5888# 0.022999f
C1251 source.n1109 a_n2390_n5888# 0.012359f
C1252 source.n1110 a_n2390_n5888# 0.013086f
C1253 source.n1111 a_n2390_n5888# 0.029211f
C1254 source.n1112 a_n2390_n5888# 0.029211f
C1255 source.n1113 a_n2390_n5888# 0.029211f
C1256 source.n1114 a_n2390_n5888# 0.013086f
C1257 source.n1115 a_n2390_n5888# 0.012359f
C1258 source.n1116 a_n2390_n5888# 0.022999f
C1259 source.n1117 a_n2390_n5888# 0.022999f
C1260 source.n1118 a_n2390_n5888# 0.012359f
C1261 source.n1119 a_n2390_n5888# 0.012722f
C1262 source.n1120 a_n2390_n5888# 0.012722f
C1263 source.n1121 a_n2390_n5888# 0.029211f
C1264 source.n1122 a_n2390_n5888# 0.029211f
C1265 source.n1123 a_n2390_n5888# 0.013086f
C1266 source.n1124 a_n2390_n5888# 0.012359f
C1267 source.n1125 a_n2390_n5888# 0.022999f
C1268 source.n1126 a_n2390_n5888# 0.022999f
C1269 source.n1127 a_n2390_n5888# 0.012359f
C1270 source.n1128 a_n2390_n5888# 0.013086f
C1271 source.n1129 a_n2390_n5888# 0.029211f
C1272 source.n1130 a_n2390_n5888# 0.029211f
C1273 source.n1131 a_n2390_n5888# 0.013086f
C1274 source.n1132 a_n2390_n5888# 0.012359f
C1275 source.n1133 a_n2390_n5888# 0.022999f
C1276 source.n1134 a_n2390_n5888# 0.022999f
C1277 source.n1135 a_n2390_n5888# 0.012359f
C1278 source.n1136 a_n2390_n5888# 0.013086f
C1279 source.n1137 a_n2390_n5888# 0.029211f
C1280 source.n1138 a_n2390_n5888# 0.06214f
C1281 source.n1139 a_n2390_n5888# 0.013086f
C1282 source.n1140 a_n2390_n5888# 0.012359f
C1283 source.n1141 a_n2390_n5888# 0.050647f
C1284 source.n1142 a_n2390_n5888# 0.034578f
C1285 source.n1143 a_n2390_n5888# 0.257474f
C1286 source.n1144 a_n2390_n5888# 2.46435f
C1287 drain_left.t10 a_n2390_n5888# 0.557233f
C1288 drain_left.t7 a_n2390_n5888# 0.557233f
C1289 drain_left.n0 a_n2390_n5888# 5.14083f
C1290 drain_left.t13 a_n2390_n5888# 0.557233f
C1291 drain_left.t14 a_n2390_n5888# 0.557233f
C1292 drain_left.n1 a_n2390_n5888# 5.1355f
C1293 drain_left.n2 a_n2390_n5888# 0.734773f
C1294 drain_left.t1 a_n2390_n5888# 0.557233f
C1295 drain_left.t6 a_n2390_n5888# 0.557233f
C1296 drain_left.n3 a_n2390_n5888# 5.14083f
C1297 drain_left.t11 a_n2390_n5888# 0.557233f
C1298 drain_left.t8 a_n2390_n5888# 0.557233f
C1299 drain_left.n4 a_n2390_n5888# 5.1355f
C1300 drain_left.n5 a_n2390_n5888# 0.734773f
C1301 drain_left.n6 a_n2390_n5888# 2.48436f
C1302 drain_left.t9 a_n2390_n5888# 0.557233f
C1303 drain_left.t2 a_n2390_n5888# 0.557233f
C1304 drain_left.n7 a_n2390_n5888# 5.14083f
C1305 drain_left.t3 a_n2390_n5888# 0.557233f
C1306 drain_left.t0 a_n2390_n5888# 0.557233f
C1307 drain_left.n8 a_n2390_n5888# 5.1355f
C1308 drain_left.n9 a_n2390_n5888# 0.774341f
C1309 drain_left.t12 a_n2390_n5888# 0.557233f
C1310 drain_left.t15 a_n2390_n5888# 0.557233f
C1311 drain_left.n10 a_n2390_n5888# 5.1355f
C1312 drain_left.n11 a_n2390_n5888# 0.384154f
C1313 drain_left.t4 a_n2390_n5888# 0.557233f
C1314 drain_left.t5 a_n2390_n5888# 0.557233f
C1315 drain_left.n12 a_n2390_n5888# 5.13549f
C1316 drain_left.n13 a_n2390_n5888# 0.630122f
C1317 plus.n0 a_n2390_n5888# 0.042711f
C1318 plus.t2 a_n2390_n5888# 1.81054f
C1319 plus.t3 a_n2390_n5888# 1.81054f
C1320 plus.t4 a_n2390_n5888# 1.81054f
C1321 plus.n1 a_n2390_n5888# 0.664841f
C1322 plus.n2 a_n2390_n5888# 0.042711f
C1323 plus.t7 a_n2390_n5888# 1.81054f
C1324 plus.t9 a_n2390_n5888# 1.81054f
C1325 plus.n3 a_n2390_n5888# 0.664841f
C1326 plus.n4 a_n2390_n5888# 0.042711f
C1327 plus.t10 a_n2390_n5888# 1.81054f
C1328 plus.t11 a_n2390_n5888# 1.81054f
C1329 plus.n5 a_n2390_n5888# 0.663656f
C1330 plus.t12 a_n2390_n5888# 1.82329f
C1331 plus.n6 a_n2390_n5888# 0.650583f
C1332 plus.n7 a_n2390_n5888# 0.143855f
C1333 plus.n8 a_n2390_n5888# 0.009692f
C1334 plus.n9 a_n2390_n5888# 0.664841f
C1335 plus.n10 a_n2390_n5888# 0.009692f
C1336 plus.n11 a_n2390_n5888# 0.042711f
C1337 plus.n12 a_n2390_n5888# 0.042711f
C1338 plus.n13 a_n2390_n5888# 0.042711f
C1339 plus.n14 a_n2390_n5888# 0.009692f
C1340 plus.n15 a_n2390_n5888# 0.664841f
C1341 plus.n16 a_n2390_n5888# 0.009692f
C1342 plus.n17 a_n2390_n5888# 0.042711f
C1343 plus.n18 a_n2390_n5888# 0.042711f
C1344 plus.n19 a_n2390_n5888# 0.042711f
C1345 plus.n20 a_n2390_n5888# 0.009692f
C1346 plus.n21 a_n2390_n5888# 0.663656f
C1347 plus.n22 a_n2390_n5888# 0.662998f
C1348 plus.n23 a_n2390_n5888# 0.777357f
C1349 plus.n24 a_n2390_n5888# 0.042711f
C1350 plus.t1 a_n2390_n5888# 1.81054f
C1351 plus.t14 a_n2390_n5888# 1.81054f
C1352 plus.t6 a_n2390_n5888# 1.81054f
C1353 plus.n25 a_n2390_n5888# 0.664841f
C1354 plus.n26 a_n2390_n5888# 0.042711f
C1355 plus.t5 a_n2390_n5888# 1.81054f
C1356 plus.t0 a_n2390_n5888# 1.81054f
C1357 plus.n27 a_n2390_n5888# 0.664841f
C1358 plus.n28 a_n2390_n5888# 0.042711f
C1359 plus.t13 a_n2390_n5888# 1.81054f
C1360 plus.t8 a_n2390_n5888# 1.81054f
C1361 plus.n29 a_n2390_n5888# 0.663656f
C1362 plus.t15 a_n2390_n5888# 1.82329f
C1363 plus.n30 a_n2390_n5888# 0.650583f
C1364 plus.n31 a_n2390_n5888# 0.143855f
C1365 plus.n32 a_n2390_n5888# 0.009692f
C1366 plus.n33 a_n2390_n5888# 0.664841f
C1367 plus.n34 a_n2390_n5888# 0.009692f
C1368 plus.n35 a_n2390_n5888# 0.042711f
C1369 plus.n36 a_n2390_n5888# 0.042711f
C1370 plus.n37 a_n2390_n5888# 0.042711f
C1371 plus.n38 a_n2390_n5888# 0.009692f
C1372 plus.n39 a_n2390_n5888# 0.664841f
C1373 plus.n40 a_n2390_n5888# 0.009692f
C1374 plus.n41 a_n2390_n5888# 0.042711f
C1375 plus.n42 a_n2390_n5888# 0.042711f
C1376 plus.n43 a_n2390_n5888# 0.042711f
C1377 plus.n44 a_n2390_n5888# 0.009692f
C1378 plus.n45 a_n2390_n5888# 0.663656f
C1379 plus.n46 a_n2390_n5888# 0.662998f
C1380 plus.n47 a_n2390_n5888# 1.78521f
.ends

