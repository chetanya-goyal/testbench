* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t25 minus.t0 drain_right.t5 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X1 source.t24 minus.t1 drain_right.t3 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X2 a_n2524_n1288# a_n2524_n1288# a_n2524_n1288# a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.8
X3 source.t23 minus.t2 drain_right.t13 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X4 source.t4 plus.t0 drain_left.t13 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X5 a_n2524_n1288# a_n2524_n1288# a_n2524_n1288# a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X6 source.t7 plus.t1 drain_left.t12 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X7 source.t10 plus.t2 drain_left.t11 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X8 drain_right.t12 minus.t3 source.t22 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X9 a_n2524_n1288# a_n2524_n1288# a_n2524_n1288# a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X10 source.t21 minus.t4 drain_right.t9 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X11 drain_right.t7 minus.t5 source.t20 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X12 drain_right.t10 minus.t6 source.t19 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X13 drain_right.t11 minus.t7 source.t18 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X14 source.t17 minus.t8 drain_right.t0 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X15 drain_right.t4 minus.t9 source.t16 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X16 drain_left.t10 plus.t3 source.t3 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X17 source.t15 minus.t10 drain_right.t1 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X18 drain_left.t9 plus.t4 source.t8 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X19 drain_right.t2 minus.t11 source.t14 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X20 drain_left.t8 plus.t5 source.t9 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X21 source.t0 plus.t6 drain_left.t7 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X22 source.t1 plus.t7 drain_left.t6 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X23 drain_right.t8 minus.t12 source.t13 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X24 drain_left.t5 plus.t8 source.t2 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X25 a_n2524_n1288# a_n2524_n1288# a_n2524_n1288# a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X26 drain_right.t6 minus.t13 source.t12 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X27 drain_left.t4 plus.t9 source.t11 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X28 source.t26 plus.t10 drain_left.t3 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X29 drain_left.t2 plus.t11 source.t27 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X30 drain_left.t1 plus.t12 source.t6 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X31 drain_left.t0 plus.t13 source.t5 a_n2524_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
R0 minus.n17 minus.n16 161.3
R1 minus.n15 minus.n0 161.3
R2 minus.n14 minus.n13 161.3
R3 minus.n12 minus.n1 161.3
R4 minus.n6 minus.n3 161.3
R5 minus.n35 minus.n34 161.3
R6 minus.n33 minus.n18 161.3
R7 minus.n32 minus.n31 161.3
R8 minus.n30 minus.n19 161.3
R9 minus.n24 minus.n21 161.3
R10 minus.n5 minus.t6 133.201
R11 minus.n23 minus.t12 133.201
R12 minus.n4 minus.t4 109.355
R13 minus.n8 minus.t3 109.355
R14 minus.n9 minus.t10 109.355
R15 minus.n10 minus.t11 109.355
R16 minus.n14 minus.t8 109.355
R17 minus.n16 minus.t5 109.355
R18 minus.n22 minus.t0 109.355
R19 minus.n26 minus.t13 109.355
R20 minus.n27 minus.t1 109.355
R21 minus.n28 minus.t7 109.355
R22 minus.n32 minus.t2 109.355
R23 minus.n34 minus.t9 109.355
R24 minus.n11 minus.n10 80.6037
R25 minus.n9 minus.n2 80.6037
R26 minus.n8 minus.n7 80.6037
R27 minus.n29 minus.n28 80.6037
R28 minus.n27 minus.n20 80.6037
R29 minus.n26 minus.n25 80.6037
R30 minus.n9 minus.n8 48.2005
R31 minus.n10 minus.n9 48.2005
R32 minus.n27 minus.n26 48.2005
R33 minus.n28 minus.n27 48.2005
R34 minus.n6 minus.n5 44.9119
R35 minus.n24 minus.n23 44.9119
R36 minus.n16 minus.n15 35.055
R37 minus.n34 minus.n33 35.055
R38 minus.n8 minus.n3 32.1338
R39 minus.n10 minus.n1 32.1338
R40 minus.n26 minus.n21 32.1338
R41 minus.n28 minus.n19 32.1338
R42 minus.n36 minus.n17 31.3319
R43 minus.n5 minus.n4 17.739
R44 minus.n23 minus.n22 17.739
R45 minus.n4 minus.n3 16.0672
R46 minus.n14 minus.n1 16.0672
R47 minus.n22 minus.n21 16.0672
R48 minus.n32 minus.n19 16.0672
R49 minus.n15 minus.n14 13.146
R50 minus.n33 minus.n32 13.146
R51 minus.n36 minus.n35 6.72588
R52 minus.n11 minus.n2 0.380177
R53 minus.n7 minus.n2 0.380177
R54 minus.n25 minus.n20 0.380177
R55 minus.n29 minus.n20 0.380177
R56 minus.n12 minus.n11 0.285035
R57 minus.n7 minus.n6 0.285035
R58 minus.n25 minus.n24 0.285035
R59 minus.n30 minus.n29 0.285035
R60 minus.n17 minus.n0 0.189894
R61 minus.n13 minus.n0 0.189894
R62 minus.n13 minus.n12 0.189894
R63 minus.n31 minus.n30 0.189894
R64 minus.n31 minus.n18 0.189894
R65 minus.n35 minus.n18 0.189894
R66 minus minus.n36 0.188
R67 drain_right.n2 drain_right.n0 289.615
R68 drain_right.n20 drain_right.n18 289.615
R69 drain_right.n3 drain_right.n2 185
R70 drain_right.n21 drain_right.n20 185
R71 drain_right.t8 drain_right.n1 167.117
R72 drain_right.t7 drain_right.n19 167.117
R73 drain_right.n15 drain_right.n13 101.769
R74 drain_right.n11 drain_right.n9 101.769
R75 drain_right.n15 drain_right.n14 100.796
R76 drain_right.n17 drain_right.n16 100.796
R77 drain_right.n11 drain_right.n10 100.796
R78 drain_right.n8 drain_right.n7 100.796
R79 drain_right.n2 drain_right.t8 52.3082
R80 drain_right.n20 drain_right.t7 52.3082
R81 drain_right.n8 drain_right.n6 49.0625
R82 drain_right.n25 drain_right.n24 48.0884
R83 drain_right drain_right.n12 24.8394
R84 drain_right.n9 drain_right.t13 9.9005
R85 drain_right.n9 drain_right.t4 9.9005
R86 drain_right.n10 drain_right.t3 9.9005
R87 drain_right.n10 drain_right.t11 9.9005
R88 drain_right.n7 drain_right.t5 9.9005
R89 drain_right.n7 drain_right.t6 9.9005
R90 drain_right.n13 drain_right.t9 9.9005
R91 drain_right.n13 drain_right.t10 9.9005
R92 drain_right.n14 drain_right.t1 9.9005
R93 drain_right.n14 drain_right.t12 9.9005
R94 drain_right.n16 drain_right.t0 9.9005
R95 drain_right.n16 drain_right.t2 9.9005
R96 drain_right.n3 drain_right.n1 9.71174
R97 drain_right.n21 drain_right.n19 9.71174
R98 drain_right.n6 drain_right.n5 9.45567
R99 drain_right.n24 drain_right.n23 9.45567
R100 drain_right.n5 drain_right.n4 9.3005
R101 drain_right.n23 drain_right.n22 9.3005
R102 drain_right.n6 drain_right.n0 8.14595
R103 drain_right.n24 drain_right.n18 8.14595
R104 drain_right.n4 drain_right.n3 7.3702
R105 drain_right.n22 drain_right.n21 7.3702
R106 drain_right drain_right.n25 6.14028
R107 drain_right.n4 drain_right.n0 5.81868
R108 drain_right.n22 drain_right.n18 5.81868
R109 drain_right.n5 drain_right.n1 3.44771
R110 drain_right.n23 drain_right.n19 3.44771
R111 drain_right.n25 drain_right.n17 0.974638
R112 drain_right.n17 drain_right.n15 0.974638
R113 drain_right.n12 drain_right.n8 0.675757
R114 drain_right.n12 drain_right.n11 0.188688
R115 source.n50 source.n48 289.615
R116 source.n36 source.n34 289.615
R117 source.n2 source.n0 289.615
R118 source.n16 source.n14 289.615
R119 source.n51 source.n50 185
R120 source.n37 source.n36 185
R121 source.n3 source.n2 185
R122 source.n17 source.n16 185
R123 source.t16 source.n49 167.117
R124 source.t27 source.n35 167.117
R125 source.t9 source.n1 167.117
R126 source.t19 source.n15 167.117
R127 source.n9 source.n8 84.1169
R128 source.n11 source.n10 84.1169
R129 source.n13 source.n12 84.1169
R130 source.n23 source.n22 84.1169
R131 source.n25 source.n24 84.1169
R132 source.n27 source.n26 84.1169
R133 source.n47 source.n46 84.1168
R134 source.n45 source.n44 84.1168
R135 source.n43 source.n42 84.1168
R136 source.n33 source.n32 84.1168
R137 source.n31 source.n30 84.1168
R138 source.n29 source.n28 84.1168
R139 source.n50 source.t16 52.3082
R140 source.n36 source.t27 52.3082
R141 source.n2 source.t9 52.3082
R142 source.n16 source.t19 52.3082
R143 source.n55 source.n54 31.4096
R144 source.n41 source.n40 31.4096
R145 source.n7 source.n6 31.4096
R146 source.n21 source.n20 31.4096
R147 source.n29 source.n27 15.6602
R148 source.n46 source.t18 9.9005
R149 source.n46 source.t23 9.9005
R150 source.n44 source.t12 9.9005
R151 source.n44 source.t24 9.9005
R152 source.n42 source.t13 9.9005
R153 source.n42 source.t25 9.9005
R154 source.n32 source.t5 9.9005
R155 source.n32 source.t4 9.9005
R156 source.n30 source.t3 9.9005
R157 source.n30 source.t7 9.9005
R158 source.n28 source.t8 9.9005
R159 source.n28 source.t10 9.9005
R160 source.n8 source.t11 9.9005
R161 source.n8 source.t0 9.9005
R162 source.n10 source.t2 9.9005
R163 source.n10 source.t1 9.9005
R164 source.n12 source.t6 9.9005
R165 source.n12 source.t26 9.9005
R166 source.n22 source.t22 9.9005
R167 source.n22 source.t21 9.9005
R168 source.n24 source.t14 9.9005
R169 source.n24 source.t15 9.9005
R170 source.n26 source.t20 9.9005
R171 source.n26 source.t17 9.9005
R172 source.n51 source.n49 9.71174
R173 source.n37 source.n35 9.71174
R174 source.n3 source.n1 9.71174
R175 source.n17 source.n15 9.71174
R176 source.n54 source.n53 9.45567
R177 source.n40 source.n39 9.45567
R178 source.n6 source.n5 9.45567
R179 source.n20 source.n19 9.45567
R180 source.n53 source.n52 9.3005
R181 source.n39 source.n38 9.3005
R182 source.n5 source.n4 9.3005
R183 source.n19 source.n18 9.3005
R184 source.n56 source.n7 8.93611
R185 source.n54 source.n48 8.14595
R186 source.n40 source.n34 8.14595
R187 source.n6 source.n0 8.14595
R188 source.n20 source.n14 8.14595
R189 source.n52 source.n51 7.3702
R190 source.n38 source.n37 7.3702
R191 source.n4 source.n3 7.3702
R192 source.n18 source.n17 7.3702
R193 source.n52 source.n48 5.81868
R194 source.n38 source.n34 5.81868
R195 source.n4 source.n0 5.81868
R196 source.n18 source.n14 5.81868
R197 source.n56 source.n55 5.7505
R198 source.n53 source.n49 3.44771
R199 source.n39 source.n35 3.44771
R200 source.n5 source.n1 3.44771
R201 source.n19 source.n15 3.44771
R202 source.n27 source.n25 0.974638
R203 source.n25 source.n23 0.974638
R204 source.n23 source.n21 0.974638
R205 source.n13 source.n11 0.974638
R206 source.n11 source.n9 0.974638
R207 source.n9 source.n7 0.974638
R208 source.n31 source.n29 0.974638
R209 source.n33 source.n31 0.974638
R210 source.n41 source.n33 0.974638
R211 source.n45 source.n43 0.974638
R212 source.n47 source.n45 0.974638
R213 source.n55 source.n47 0.974638
R214 source.n21 source.n13 0.957397
R215 source.n43 source.n41 0.957397
R216 source source.n56 0.188
R217 plus.n7 plus.n6 161.3
R218 plus.n13 plus.n12 161.3
R219 plus.n14 plus.n1 161.3
R220 plus.n15 plus.n0 161.3
R221 plus.n17 plus.n16 161.3
R222 plus.n25 plus.n24 161.3
R223 plus.n31 plus.n30 161.3
R224 plus.n32 plus.n19 161.3
R225 plus.n33 plus.n18 161.3
R226 plus.n35 plus.n34 161.3
R227 plus.n5 plus.t12 133.201
R228 plus.n23 plus.t11 133.201
R229 plus.n16 plus.t5 109.355
R230 plus.n14 plus.t6 109.355
R231 plus.n2 plus.t9 109.355
R232 plus.n9 plus.t7 109.355
R233 plus.n8 plus.t8 109.355
R234 plus.n4 plus.t10 109.355
R235 plus.n34 plus.t4 109.355
R236 plus.n32 plus.t2 109.355
R237 plus.n20 plus.t3 109.355
R238 plus.n27 plus.t1 109.355
R239 plus.n26 plus.t13 109.355
R240 plus.n22 plus.t0 109.355
R241 plus.n8 plus.n3 80.6037
R242 plus.n10 plus.n9 80.6037
R243 plus.n11 plus.n2 80.6037
R244 plus.n26 plus.n21 80.6037
R245 plus.n28 plus.n27 80.6037
R246 plus.n29 plus.n20 80.6037
R247 plus.n9 plus.n2 48.2005
R248 plus.n9 plus.n8 48.2005
R249 plus.n27 plus.n20 48.2005
R250 plus.n27 plus.n26 48.2005
R251 plus.n24 plus.n23 44.9119
R252 plus.n6 plus.n5 44.9119
R253 plus.n16 plus.n15 35.055
R254 plus.n34 plus.n33 35.055
R255 plus.n13 plus.n2 32.1338
R256 plus.n8 plus.n7 32.1338
R257 plus.n31 plus.n20 32.1338
R258 plus.n26 plus.n25 32.1338
R259 plus plus.n35 29.0009
R260 plus.n23 plus.n22 17.739
R261 plus.n5 plus.n4 17.739
R262 plus.n14 plus.n13 16.0672
R263 plus.n7 plus.n4 16.0672
R264 plus.n32 plus.n31 16.0672
R265 plus.n25 plus.n22 16.0672
R266 plus.n15 plus.n14 13.146
R267 plus.n33 plus.n32 13.146
R268 plus plus.n17 8.58194
R269 plus.n10 plus.n3 0.380177
R270 plus.n11 plus.n10 0.380177
R271 plus.n29 plus.n28 0.380177
R272 plus.n28 plus.n21 0.380177
R273 plus.n6 plus.n3 0.285035
R274 plus.n12 plus.n11 0.285035
R275 plus.n30 plus.n29 0.285035
R276 plus.n24 plus.n21 0.285035
R277 plus.n12 plus.n1 0.189894
R278 plus.n1 plus.n0 0.189894
R279 plus.n17 plus.n0 0.189894
R280 plus.n35 plus.n18 0.189894
R281 plus.n19 plus.n18 0.189894
R282 plus.n30 plus.n19 0.189894
R283 drain_left.n2 drain_left.n0 289.615
R284 drain_left.n15 drain_left.n13 289.615
R285 drain_left.n3 drain_left.n2 185
R286 drain_left.n16 drain_left.n15 185
R287 drain_left.t9 drain_left.n1 167.117
R288 drain_left.t1 drain_left.n14 167.117
R289 drain_left.n11 drain_left.n9 101.769
R290 drain_left.n25 drain_left.n24 100.796
R291 drain_left.n23 drain_left.n22 100.796
R292 drain_left.n21 drain_left.n20 100.796
R293 drain_left.n11 drain_left.n10 100.796
R294 drain_left.n8 drain_left.n7 100.796
R295 drain_left.n2 drain_left.t9 52.3082
R296 drain_left.n15 drain_left.t1 52.3082
R297 drain_left.n8 drain_left.n6 49.0625
R298 drain_left.n21 drain_left.n19 49.0625
R299 drain_left drain_left.n12 25.3926
R300 drain_left.n9 drain_left.t13 9.9005
R301 drain_left.n9 drain_left.t2 9.9005
R302 drain_left.n10 drain_left.t12 9.9005
R303 drain_left.n10 drain_left.t0 9.9005
R304 drain_left.n7 drain_left.t11 9.9005
R305 drain_left.n7 drain_left.t10 9.9005
R306 drain_left.n24 drain_left.t7 9.9005
R307 drain_left.n24 drain_left.t8 9.9005
R308 drain_left.n22 drain_left.t6 9.9005
R309 drain_left.n22 drain_left.t4 9.9005
R310 drain_left.n20 drain_left.t3 9.9005
R311 drain_left.n20 drain_left.t5 9.9005
R312 drain_left.n3 drain_left.n1 9.71174
R313 drain_left.n16 drain_left.n14 9.71174
R314 drain_left.n6 drain_left.n5 9.45567
R315 drain_left.n19 drain_left.n18 9.45567
R316 drain_left.n5 drain_left.n4 9.3005
R317 drain_left.n18 drain_left.n17 9.3005
R318 drain_left.n6 drain_left.n0 8.14595
R319 drain_left.n19 drain_left.n13 8.14595
R320 drain_left.n4 drain_left.n3 7.3702
R321 drain_left.n17 drain_left.n16 7.3702
R322 drain_left drain_left.n25 6.62735
R323 drain_left.n4 drain_left.n0 5.81868
R324 drain_left.n17 drain_left.n13 5.81868
R325 drain_left.n5 drain_left.n1 3.44771
R326 drain_left.n18 drain_left.n14 3.44771
R327 drain_left.n23 drain_left.n21 0.974638
R328 drain_left.n25 drain_left.n23 0.974638
R329 drain_left.n12 drain_left.n8 0.675757
R330 drain_left.n12 drain_left.n11 0.188688
C0 minus drain_right 2.07761f
C1 minus plus 4.44261f
C2 source drain_right 5.73694f
C3 source plus 2.68183f
C4 minus drain_left 0.179749f
C5 source drain_left 5.7363f
C6 drain_right plus 0.414177f
C7 minus source 2.66778f
C8 drain_right drain_left 1.31403f
C9 drain_left plus 2.32692f
C10 drain_right a_n2524_n1288# 4.87615f
C11 drain_left a_n2524_n1288# 5.2597f
C12 source a_n2524_n1288# 2.843657f
C13 minus a_n2524_n1288# 9.204286f
C14 plus a_n2524_n1288# 10.459149f
C15 drain_left.n0 a_n2524_n1288# 0.036604f
C16 drain_left.n1 a_n2524_n1288# 0.080992f
C17 drain_left.t9 a_n2524_n1288# 0.06078f
C18 drain_left.n2 a_n2524_n1288# 0.063387f
C19 drain_left.n3 a_n2524_n1288# 0.020434f
C20 drain_left.n4 a_n2524_n1288# 0.013476f
C21 drain_left.n5 a_n2524_n1288# 0.178526f
C22 drain_left.n6 a_n2524_n1288# 0.059961f
C23 drain_left.t11 a_n2524_n1288# 0.039637f
C24 drain_left.t10 a_n2524_n1288# 0.039637f
C25 drain_left.n7 a_n2524_n1288# 0.249009f
C26 drain_left.n8 a_n2524_n1288# 0.449824f
C27 drain_left.t13 a_n2524_n1288# 0.039637f
C28 drain_left.t2 a_n2524_n1288# 0.039637f
C29 drain_left.n9 a_n2524_n1288# 0.25245f
C30 drain_left.t12 a_n2524_n1288# 0.039637f
C31 drain_left.t0 a_n2524_n1288# 0.039637f
C32 drain_left.n10 a_n2524_n1288# 0.249009f
C33 drain_left.n11 a_n2524_n1288# 0.645025f
C34 drain_left.n12 a_n2524_n1288# 0.911513f
C35 drain_left.n13 a_n2524_n1288# 0.036604f
C36 drain_left.n14 a_n2524_n1288# 0.080992f
C37 drain_left.t1 a_n2524_n1288# 0.06078f
C38 drain_left.n15 a_n2524_n1288# 0.063387f
C39 drain_left.n16 a_n2524_n1288# 0.020434f
C40 drain_left.n17 a_n2524_n1288# 0.013476f
C41 drain_left.n18 a_n2524_n1288# 0.178526f
C42 drain_left.n19 a_n2524_n1288# 0.059961f
C43 drain_left.t3 a_n2524_n1288# 0.039637f
C44 drain_left.t5 a_n2524_n1288# 0.039637f
C45 drain_left.n20 a_n2524_n1288# 0.24901f
C46 drain_left.n21 a_n2524_n1288# 0.473115f
C47 drain_left.t6 a_n2524_n1288# 0.039637f
C48 drain_left.t4 a_n2524_n1288# 0.039637f
C49 drain_left.n22 a_n2524_n1288# 0.24901f
C50 drain_left.n23 a_n2524_n1288# 0.349393f
C51 drain_left.t7 a_n2524_n1288# 0.039637f
C52 drain_left.t8 a_n2524_n1288# 0.039637f
C53 drain_left.n24 a_n2524_n1288# 0.24901f
C54 drain_left.n25 a_n2524_n1288# 0.574275f
C55 plus.n0 a_n2524_n1288# 0.04375f
C56 plus.t5 a_n2524_n1288# 0.216771f
C57 plus.t6 a_n2524_n1288# 0.216771f
C58 plus.n1 a_n2524_n1288# 0.04375f
C59 plus.t9 a_n2524_n1288# 0.216771f
C60 plus.n2 a_n2524_n1288# 0.157152f
C61 plus.n3 a_n2524_n1288# 0.072871f
C62 plus.t7 a_n2524_n1288# 0.216771f
C63 plus.t8 a_n2524_n1288# 0.216771f
C64 plus.t10 a_n2524_n1288# 0.216771f
C65 plus.n4 a_n2524_n1288# 0.152104f
C66 plus.t12 a_n2524_n1288# 0.243525f
C67 plus.n5 a_n2524_n1288# 0.126474f
C68 plus.n6 a_n2524_n1288# 0.204319f
C69 plus.n7 a_n2524_n1288# 0.009928f
C70 plus.n8 a_n2524_n1288# 0.157152f
C71 plus.n9 a_n2524_n1288# 0.160119f
C72 plus.n10 a_n2524_n1288# 0.0875f
C73 plus.n11 a_n2524_n1288# 0.072871f
C74 plus.n12 a_n2524_n1288# 0.058379f
C75 plus.n13 a_n2524_n1288# 0.009928f
C76 plus.n14 a_n2524_n1288# 0.146685f
C77 plus.n15 a_n2524_n1288# 0.009928f
C78 plus.n16 a_n2524_n1288# 0.147764f
C79 plus.n17 a_n2524_n1288# 0.337075f
C80 plus.n18 a_n2524_n1288# 0.04375f
C81 plus.t4 a_n2524_n1288# 0.216771f
C82 plus.n19 a_n2524_n1288# 0.04375f
C83 plus.t2 a_n2524_n1288# 0.216771f
C84 plus.t3 a_n2524_n1288# 0.216771f
C85 plus.n20 a_n2524_n1288# 0.157152f
C86 plus.n21 a_n2524_n1288# 0.072871f
C87 plus.t1 a_n2524_n1288# 0.216771f
C88 plus.t13 a_n2524_n1288# 0.216771f
C89 plus.t0 a_n2524_n1288# 0.216771f
C90 plus.n22 a_n2524_n1288# 0.152104f
C91 plus.t11 a_n2524_n1288# 0.243525f
C92 plus.n23 a_n2524_n1288# 0.126474f
C93 plus.n24 a_n2524_n1288# 0.204319f
C94 plus.n25 a_n2524_n1288# 0.009928f
C95 plus.n26 a_n2524_n1288# 0.157152f
C96 plus.n27 a_n2524_n1288# 0.160119f
C97 plus.n28 a_n2524_n1288# 0.0875f
C98 plus.n29 a_n2524_n1288# 0.072871f
C99 plus.n30 a_n2524_n1288# 0.058379f
C100 plus.n31 a_n2524_n1288# 0.009928f
C101 plus.n32 a_n2524_n1288# 0.146685f
C102 plus.n33 a_n2524_n1288# 0.009928f
C103 plus.n34 a_n2524_n1288# 0.147764f
C104 plus.n35 a_n2524_n1288# 1.17413f
C105 source.n0 a_n2524_n1288# 0.048648f
C106 source.n1 a_n2524_n1288# 0.107641f
C107 source.t9 a_n2524_n1288# 0.080779f
C108 source.n2 a_n2524_n1288# 0.084244f
C109 source.n3 a_n2524_n1288# 0.027157f
C110 source.n4 a_n2524_n1288# 0.017911f
C111 source.n5 a_n2524_n1288# 0.237266f
C112 source.n6 a_n2524_n1288# 0.05333f
C113 source.n7 a_n2524_n1288# 0.5852f
C114 source.t11 a_n2524_n1288# 0.052678f
C115 source.t0 a_n2524_n1288# 0.052678f
C116 source.n8 a_n2524_n1288# 0.281615f
C117 source.n9 a_n2524_n1288# 0.468375f
C118 source.t2 a_n2524_n1288# 0.052678f
C119 source.t1 a_n2524_n1288# 0.052678f
C120 source.n10 a_n2524_n1288# 0.281615f
C121 source.n11 a_n2524_n1288# 0.468375f
C122 source.t6 a_n2524_n1288# 0.052678f
C123 source.t26 a_n2524_n1288# 0.052678f
C124 source.n12 a_n2524_n1288# 0.281615f
C125 source.n13 a_n2524_n1288# 0.466524f
C126 source.n14 a_n2524_n1288# 0.048648f
C127 source.n15 a_n2524_n1288# 0.107641f
C128 source.t19 a_n2524_n1288# 0.080779f
C129 source.n16 a_n2524_n1288# 0.084244f
C130 source.n17 a_n2524_n1288# 0.027157f
C131 source.n18 a_n2524_n1288# 0.017911f
C132 source.n19 a_n2524_n1288# 0.237266f
C133 source.n20 a_n2524_n1288# 0.05333f
C134 source.n21 a_n2524_n1288# 0.234831f
C135 source.t22 a_n2524_n1288# 0.052678f
C136 source.t21 a_n2524_n1288# 0.052678f
C137 source.n22 a_n2524_n1288# 0.281615f
C138 source.n23 a_n2524_n1288# 0.468375f
C139 source.t14 a_n2524_n1288# 0.052678f
C140 source.t15 a_n2524_n1288# 0.052678f
C141 source.n24 a_n2524_n1288# 0.281615f
C142 source.n25 a_n2524_n1288# 0.468375f
C143 source.t20 a_n2524_n1288# 0.052678f
C144 source.t17 a_n2524_n1288# 0.052678f
C145 source.n26 a_n2524_n1288# 0.281615f
C146 source.n27 a_n2524_n1288# 1.24289f
C147 source.t8 a_n2524_n1288# 0.052678f
C148 source.t10 a_n2524_n1288# 0.052678f
C149 source.n28 a_n2524_n1288# 0.281614f
C150 source.n29 a_n2524_n1288# 1.24289f
C151 source.t3 a_n2524_n1288# 0.052678f
C152 source.t7 a_n2524_n1288# 0.052678f
C153 source.n30 a_n2524_n1288# 0.281614f
C154 source.n31 a_n2524_n1288# 0.468377f
C155 source.t5 a_n2524_n1288# 0.052678f
C156 source.t4 a_n2524_n1288# 0.052678f
C157 source.n32 a_n2524_n1288# 0.281614f
C158 source.n33 a_n2524_n1288# 0.468377f
C159 source.n34 a_n2524_n1288# 0.048648f
C160 source.n35 a_n2524_n1288# 0.107641f
C161 source.t27 a_n2524_n1288# 0.080779f
C162 source.n36 a_n2524_n1288# 0.084244f
C163 source.n37 a_n2524_n1288# 0.027157f
C164 source.n38 a_n2524_n1288# 0.017911f
C165 source.n39 a_n2524_n1288# 0.237266f
C166 source.n40 a_n2524_n1288# 0.05333f
C167 source.n41 a_n2524_n1288# 0.234831f
C168 source.t13 a_n2524_n1288# 0.052678f
C169 source.t25 a_n2524_n1288# 0.052678f
C170 source.n42 a_n2524_n1288# 0.281614f
C171 source.n43 a_n2524_n1288# 0.466525f
C172 source.t12 a_n2524_n1288# 0.052678f
C173 source.t24 a_n2524_n1288# 0.052678f
C174 source.n44 a_n2524_n1288# 0.281614f
C175 source.n45 a_n2524_n1288# 0.468377f
C176 source.t18 a_n2524_n1288# 0.052678f
C177 source.t23 a_n2524_n1288# 0.052678f
C178 source.n46 a_n2524_n1288# 0.281614f
C179 source.n47 a_n2524_n1288# 0.468377f
C180 source.n48 a_n2524_n1288# 0.048648f
C181 source.n49 a_n2524_n1288# 0.107641f
C182 source.t16 a_n2524_n1288# 0.080779f
C183 source.n50 a_n2524_n1288# 0.084244f
C184 source.n51 a_n2524_n1288# 0.027157f
C185 source.n52 a_n2524_n1288# 0.017911f
C186 source.n53 a_n2524_n1288# 0.237266f
C187 source.n54 a_n2524_n1288# 0.05333f
C188 source.n55 a_n2524_n1288# 0.407154f
C189 source.n56 a_n2524_n1288# 0.844496f
C190 drain_right.n0 a_n2524_n1288# 0.036132f
C191 drain_right.n1 a_n2524_n1288# 0.079948f
C192 drain_right.t8 a_n2524_n1288# 0.059997f
C193 drain_right.n2 a_n2524_n1288# 0.06257f
C194 drain_right.n3 a_n2524_n1288# 0.02017f
C195 drain_right.n4 a_n2524_n1288# 0.013303f
C196 drain_right.n5 a_n2524_n1288# 0.176224f
C197 drain_right.n6 a_n2524_n1288# 0.059188f
C198 drain_right.t5 a_n2524_n1288# 0.039125f
C199 drain_right.t6 a_n2524_n1288# 0.039125f
C200 drain_right.n7 a_n2524_n1288# 0.245798f
C201 drain_right.n8 a_n2524_n1288# 0.444023f
C202 drain_right.t13 a_n2524_n1288# 0.039125f
C203 drain_right.t4 a_n2524_n1288# 0.039125f
C204 drain_right.n9 a_n2524_n1288# 0.249194f
C205 drain_right.t3 a_n2524_n1288# 0.039125f
C206 drain_right.t11 a_n2524_n1288# 0.039125f
C207 drain_right.n10 a_n2524_n1288# 0.245798f
C208 drain_right.n11 a_n2524_n1288# 0.636707f
C209 drain_right.n12 a_n2524_n1288# 0.851571f
C210 drain_right.t9 a_n2524_n1288# 0.039125f
C211 drain_right.t10 a_n2524_n1288# 0.039125f
C212 drain_right.n13 a_n2524_n1288# 0.249196f
C213 drain_right.t1 a_n2524_n1288# 0.039125f
C214 drain_right.t12 a_n2524_n1288# 0.039125f
C215 drain_right.n14 a_n2524_n1288# 0.245799f
C216 drain_right.n15 a_n2524_n1288# 0.69635f
C217 drain_right.t0 a_n2524_n1288# 0.039125f
C218 drain_right.t2 a_n2524_n1288# 0.039125f
C219 drain_right.n16 a_n2524_n1288# 0.245799f
C220 drain_right.n17 a_n2524_n1288# 0.344888f
C221 drain_right.n18 a_n2524_n1288# 0.036132f
C222 drain_right.n19 a_n2524_n1288# 0.079948f
C223 drain_right.t7 a_n2524_n1288# 0.059997f
C224 drain_right.n20 a_n2524_n1288# 0.06257f
C225 drain_right.n21 a_n2524_n1288# 0.02017f
C226 drain_right.n22 a_n2524_n1288# 0.013303f
C227 drain_right.n23 a_n2524_n1288# 0.176224f
C228 drain_right.n24 a_n2524_n1288# 0.056714f
C229 drain_right.n25 a_n2524_n1288# 0.357304f
C230 minus.n0 a_n2524_n1288# 0.04242f
C231 minus.n1 a_n2524_n1288# 0.009626f
C232 minus.t8 a_n2524_n1288# 0.210181f
C233 minus.n2 a_n2524_n1288# 0.08484f
C234 minus.n3 a_n2524_n1288# 0.009626f
C235 minus.t3 a_n2524_n1288# 0.210181f
C236 minus.t6 a_n2524_n1288# 0.236121f
C237 minus.t4 a_n2524_n1288# 0.210181f
C238 minus.n4 a_n2524_n1288# 0.14748f
C239 minus.n5 a_n2524_n1288# 0.122628f
C240 minus.n6 a_n2524_n1288# 0.198107f
C241 minus.n7 a_n2524_n1288# 0.070656f
C242 minus.n8 a_n2524_n1288# 0.152374f
C243 minus.t10 a_n2524_n1288# 0.210181f
C244 minus.n9 a_n2524_n1288# 0.155251f
C245 minus.t11 a_n2524_n1288# 0.210181f
C246 minus.n10 a_n2524_n1288# 0.152374f
C247 minus.n11 a_n2524_n1288# 0.070656f
C248 minus.n12 a_n2524_n1288# 0.056604f
C249 minus.n13 a_n2524_n1288# 0.04242f
C250 minus.n14 a_n2524_n1288# 0.142225f
C251 minus.n15 a_n2524_n1288# 0.009626f
C252 minus.t5 a_n2524_n1288# 0.210181f
C253 minus.n16 a_n2524_n1288# 0.143271f
C254 minus.n17 a_n2524_n1288# 1.19607f
C255 minus.n18 a_n2524_n1288# 0.04242f
C256 minus.n19 a_n2524_n1288# 0.009626f
C257 minus.n20 a_n2524_n1288# 0.08484f
C258 minus.n21 a_n2524_n1288# 0.009626f
C259 minus.t12 a_n2524_n1288# 0.236121f
C260 minus.t0 a_n2524_n1288# 0.210181f
C261 minus.n22 a_n2524_n1288# 0.14748f
C262 minus.n23 a_n2524_n1288# 0.122628f
C263 minus.n24 a_n2524_n1288# 0.198107f
C264 minus.n25 a_n2524_n1288# 0.070656f
C265 minus.t13 a_n2524_n1288# 0.210181f
C266 minus.n26 a_n2524_n1288# 0.152374f
C267 minus.t1 a_n2524_n1288# 0.210181f
C268 minus.n27 a_n2524_n1288# 0.155251f
C269 minus.t7 a_n2524_n1288# 0.210181f
C270 minus.n28 a_n2524_n1288# 0.152374f
C271 minus.n29 a_n2524_n1288# 0.070656f
C272 minus.n30 a_n2524_n1288# 0.056604f
C273 minus.n31 a_n2524_n1288# 0.04242f
C274 minus.t2 a_n2524_n1288# 0.210181f
C275 minus.n32 a_n2524_n1288# 0.142225f
C276 minus.n33 a_n2524_n1288# 0.009626f
C277 minus.t9 a_n2524_n1288# 0.210181f
C278 minus.n34 a_n2524_n1288# 0.143271f
C279 minus.n35 a_n2524_n1288# 0.29967f
C280 minus.n36 a_n2524_n1288# 1.46162f
.ends

