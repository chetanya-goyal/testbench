* NGSPICE file created from diffpair326.ext - technology: sky130A

.subckt diffpair326 minus drain_right drain_left source plus
X0 a_n1756_n2688# a_n1756_n2688# a_n1756_n2688# a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=34.2 ps=151.6 w=9 l=0.15
X1 drain_left.t13 plus.t0 source.t23 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X2 a_n1756_n2688# a_n1756_n2688# a_n1756_n2688# a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X3 drain_left.t12 plus.t1 source.t18 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X4 source.t15 plus.t2 drain_left.t11 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X5 a_n1756_n2688# a_n1756_n2688# a_n1756_n2688# a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X6 drain_right.t13 minus.t0 source.t6 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X7 drain_left.t10 plus.t3 source.t24 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X8 source.t8 minus.t1 drain_right.t12 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X9 drain_left.t9 plus.t4 source.t27 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X10 a_n1756_n2688# a_n1756_n2688# a_n1756_n2688# a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X11 source.t0 minus.t2 drain_right.t11 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X12 source.t11 minus.t3 drain_right.t10 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X13 source.t21 plus.t5 drain_left.t8 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X14 drain_right.t9 minus.t4 source.t2 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X15 drain_right.t8 minus.t5 source.t1 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X16 drain_right.t7 minus.t6 source.t13 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X17 source.t4 minus.t7 drain_right.t6 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X18 drain_right.t5 minus.t8 source.t12 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X19 drain_left.t7 plus.t6 source.t16 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X20 drain_right.t4 minus.t9 source.t5 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X21 drain_right.t3 minus.t10 source.t7 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X22 source.t26 plus.t7 drain_left.t6 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X23 source.t9 minus.t11 drain_right.t2 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X24 source.t3 minus.t12 drain_right.t1 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X25 drain_left.t5 plus.t8 source.t25 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X26 drain_left.t4 plus.t9 source.t19 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X27 source.t14 plus.t10 drain_left.t3 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X28 source.t20 plus.t11 drain_left.t2 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X29 drain_right.t0 minus.t13 source.t10 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X30 source.t22 plus.t12 drain_left.t1 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X31 drain_left.t0 plus.t13 source.t17 a_n1756_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
R0 plus.n3 plus.t6 1720.59
R1 plus.n15 plus.t8 1720.59
R2 plus.n20 plus.t3 1720.59
R3 plus.n32 plus.t1 1720.59
R4 plus.n1 plus.t7 1654.87
R5 plus.n4 plus.t11 1654.87
R6 plus.n6 plus.t9 1654.87
R7 plus.n12 plus.t13 1654.87
R8 plus.n14 plus.t10 1654.87
R9 plus.n18 plus.t2 1654.87
R10 plus.n21 plus.t5 1654.87
R11 plus.n23 plus.t0 1654.87
R12 plus.n29 plus.t4 1654.87
R13 plus.n31 plus.t12 1654.87
R14 plus.n3 plus.n2 161.489
R15 plus.n20 plus.n19 161.489
R16 plus.n5 plus.n2 161.3
R17 plus.n8 plus.n7 161.3
R18 plus.n9 plus.n1 161.3
R19 plus.n11 plus.n10 161.3
R20 plus.n13 plus.n0 161.3
R21 plus.n16 plus.n15 161.3
R22 plus.n22 plus.n19 161.3
R23 plus.n25 plus.n24 161.3
R24 plus.n26 plus.n18 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n17 161.3
R27 plus.n33 plus.n32 161.3
R28 plus.n7 plus.n1 73.0308
R29 plus.n11 plus.n1 73.0308
R30 plus.n28 plus.n18 73.0308
R31 plus.n24 plus.n18 73.0308
R32 plus.n6 plus.n5 51.1217
R33 plus.n13 plus.n12 51.1217
R34 plus.n30 plus.n29 51.1217
R35 plus.n23 plus.n22 51.1217
R36 plus.n5 plus.n4 43.8187
R37 plus.n14 plus.n13 43.8187
R38 plus.n31 plus.n30 43.8187
R39 plus.n22 plus.n21 43.8187
R40 plus.n4 plus.n3 29.2126
R41 plus.n15 plus.n14 29.2126
R42 plus.n32 plus.n31 29.2126
R43 plus.n21 plus.n20 29.2126
R44 plus plus.n33 28.588
R45 plus.n7 plus.n6 21.9096
R46 plus.n12 plus.n11 21.9096
R47 plus.n29 plus.n28 21.9096
R48 plus.n24 plus.n23 21.9096
R49 plus plus.n16 11.0782
R50 plus.n8 plus.n2 0.189894
R51 plus.n9 plus.n8 0.189894
R52 plus.n10 plus.n9 0.189894
R53 plus.n10 plus.n0 0.189894
R54 plus.n16 plus.n0 0.189894
R55 plus.n33 plus.n17 0.189894
R56 plus.n27 plus.n17 0.189894
R57 plus.n27 plus.n26 0.189894
R58 plus.n26 plus.n25 0.189894
R59 plus.n25 plus.n19 0.189894
R60 source.n7 source.t2 52.1921
R61 source.n27 source.t12 52.1919
R62 source.n20 source.t24 52.1919
R63 source.n0 source.t25 52.1919
R64 source.n2 source.n1 48.8588
R65 source.n4 source.n3 48.8588
R66 source.n6 source.n5 48.8588
R67 source.n9 source.n8 48.8588
R68 source.n11 source.n10 48.8588
R69 source.n13 source.n12 48.8588
R70 source.n26 source.n25 48.8586
R71 source.n24 source.n23 48.8586
R72 source.n22 source.n21 48.8586
R73 source.n19 source.n18 48.8586
R74 source.n17 source.n16 48.8586
R75 source.n15 source.n14 48.8586
R76 source.n15 source.n13 20.1357
R77 source.n28 source.n0 14.0322
R78 source.n28 source.n27 5.5436
R79 source.n25 source.t6 3.33383
R80 source.n25 source.t0 3.33383
R81 source.n23 source.t13 3.33383
R82 source.n23 source.t3 3.33383
R83 source.n21 source.t10 3.33383
R84 source.n21 source.t8 3.33383
R85 source.n18 source.t23 3.33383
R86 source.n18 source.t21 3.33383
R87 source.n16 source.t27 3.33383
R88 source.n16 source.t15 3.33383
R89 source.n14 source.t18 3.33383
R90 source.n14 source.t22 3.33383
R91 source.n1 source.t17 3.33383
R92 source.n1 source.t14 3.33383
R93 source.n3 source.t19 3.33383
R94 source.n3 source.t26 3.33383
R95 source.n5 source.t16 3.33383
R96 source.n5 source.t20 3.33383
R97 source.n8 source.t5 3.33383
R98 source.n8 source.t11 3.33383
R99 source.n10 source.t1 3.33383
R100 source.n10 source.t4 3.33383
R101 source.n12 source.t7 3.33383
R102 source.n12 source.t9 3.33383
R103 source.n7 source.n6 0.7505
R104 source.n22 source.n20 0.7505
R105 source.n13 source.n11 0.560845
R106 source.n11 source.n9 0.560845
R107 source.n9 source.n7 0.560845
R108 source.n6 source.n4 0.560845
R109 source.n4 source.n2 0.560845
R110 source.n2 source.n0 0.560845
R111 source.n17 source.n15 0.560845
R112 source.n19 source.n17 0.560845
R113 source.n20 source.n19 0.560845
R114 source.n24 source.n22 0.560845
R115 source.n26 source.n24 0.560845
R116 source.n27 source.n26 0.560845
R117 source source.n28 0.188
R118 drain_left.n7 drain_left.t7 69.4313
R119 drain_left.n1 drain_left.t12 69.431
R120 drain_left.n4 drain_left.n2 66.0977
R121 drain_left.n9 drain_left.n8 65.5376
R122 drain_left.n7 drain_left.n6 65.5376
R123 drain_left.n11 drain_left.n10 65.5374
R124 drain_left.n4 drain_left.n3 65.5373
R125 drain_left.n1 drain_left.n0 65.5373
R126 drain_left drain_left.n5 28.3163
R127 drain_left drain_left.n11 6.21356
R128 drain_left.n2 drain_left.t8 3.33383
R129 drain_left.n2 drain_left.t10 3.33383
R130 drain_left.n3 drain_left.t11 3.33383
R131 drain_left.n3 drain_left.t13 3.33383
R132 drain_left.n0 drain_left.t1 3.33383
R133 drain_left.n0 drain_left.t9 3.33383
R134 drain_left.n10 drain_left.t3 3.33383
R135 drain_left.n10 drain_left.t5 3.33383
R136 drain_left.n8 drain_left.t6 3.33383
R137 drain_left.n8 drain_left.t0 3.33383
R138 drain_left.n6 drain_left.t2 3.33383
R139 drain_left.n6 drain_left.t4 3.33383
R140 drain_left.n9 drain_left.n7 0.560845
R141 drain_left.n11 drain_left.n9 0.560845
R142 drain_left.n5 drain_left.n1 0.365413
R143 drain_left.n5 drain_left.n4 0.0852402
R144 minus.n15 minus.t10 1720.59
R145 minus.n3 minus.t4 1720.59
R146 minus.n32 minus.t8 1720.59
R147 minus.n20 minus.t13 1720.59
R148 minus.n1 minus.t7 1654.87
R149 minus.n14 minus.t11 1654.87
R150 minus.n12 minus.t5 1654.87
R151 minus.n6 minus.t9 1654.87
R152 minus.n4 minus.t3 1654.87
R153 minus.n18 minus.t12 1654.87
R154 minus.n31 minus.t2 1654.87
R155 minus.n29 minus.t0 1654.87
R156 minus.n23 minus.t6 1654.87
R157 minus.n21 minus.t1 1654.87
R158 minus.n3 minus.n2 161.489
R159 minus.n20 minus.n19 161.489
R160 minus.n16 minus.n15 161.3
R161 minus.n13 minus.n0 161.3
R162 minus.n11 minus.n10 161.3
R163 minus.n9 minus.n1 161.3
R164 minus.n8 minus.n7 161.3
R165 minus.n5 minus.n2 161.3
R166 minus.n33 minus.n32 161.3
R167 minus.n30 minus.n17 161.3
R168 minus.n28 minus.n27 161.3
R169 minus.n26 minus.n18 161.3
R170 minus.n25 minus.n24 161.3
R171 minus.n22 minus.n19 161.3
R172 minus.n11 minus.n1 73.0308
R173 minus.n7 minus.n1 73.0308
R174 minus.n24 minus.n18 73.0308
R175 minus.n28 minus.n18 73.0308
R176 minus.n13 minus.n12 51.1217
R177 minus.n6 minus.n5 51.1217
R178 minus.n23 minus.n22 51.1217
R179 minus.n30 minus.n29 51.1217
R180 minus.n14 minus.n13 43.8187
R181 minus.n5 minus.n4 43.8187
R182 minus.n22 minus.n21 43.8187
R183 minus.n31 minus.n30 43.8187
R184 minus.n34 minus.n16 33.5706
R185 minus.n15 minus.n14 29.2126
R186 minus.n4 minus.n3 29.2126
R187 minus.n21 minus.n20 29.2126
R188 minus.n32 minus.n31 29.2126
R189 minus.n12 minus.n11 21.9096
R190 minus.n7 minus.n6 21.9096
R191 minus.n24 minus.n23 21.9096
R192 minus.n29 minus.n28 21.9096
R193 minus.n34 minus.n33 6.57058
R194 minus.n16 minus.n0 0.189894
R195 minus.n10 minus.n0 0.189894
R196 minus.n10 minus.n9 0.189894
R197 minus.n9 minus.n8 0.189894
R198 minus.n8 minus.n2 0.189894
R199 minus.n25 minus.n19 0.189894
R200 minus.n26 minus.n25 0.189894
R201 minus.n27 minus.n26 0.189894
R202 minus.n27 minus.n17 0.189894
R203 minus.n33 minus.n17 0.189894
R204 minus minus.n34 0.188
R205 drain_right.n1 drain_right.t0 69.431
R206 drain_right.n11 drain_right.t3 68.8709
R207 drain_right.n8 drain_right.n6 66.0978
R208 drain_right.n4 drain_right.n2 66.0977
R209 drain_right.n8 drain_right.n7 65.5376
R210 drain_right.n10 drain_right.n9 65.5376
R211 drain_right.n4 drain_right.n3 65.5373
R212 drain_right.n1 drain_right.n0 65.5373
R213 drain_right drain_right.n5 27.7631
R214 drain_right drain_right.n11 5.93339
R215 drain_right.n2 drain_right.t11 3.33383
R216 drain_right.n2 drain_right.t5 3.33383
R217 drain_right.n3 drain_right.t1 3.33383
R218 drain_right.n3 drain_right.t13 3.33383
R219 drain_right.n0 drain_right.t12 3.33383
R220 drain_right.n0 drain_right.t7 3.33383
R221 drain_right.n6 drain_right.t10 3.33383
R222 drain_right.n6 drain_right.t9 3.33383
R223 drain_right.n7 drain_right.t6 3.33383
R224 drain_right.n7 drain_right.t4 3.33383
R225 drain_right.n9 drain_right.t2 3.33383
R226 drain_right.n9 drain_right.t8 3.33383
R227 drain_right.n11 drain_right.n10 0.560845
R228 drain_right.n10 drain_right.n8 0.560845
R229 drain_right.n5 drain_right.n1 0.365413
R230 drain_right.n5 drain_right.n4 0.0852402
C0 source drain_left 22.1185f
C1 drain_right minus 2.51387f
C2 drain_right plus 0.325592f
C3 plus minus 4.76842f
C4 drain_right drain_left 0.900167f
C5 drain_right source 22.1106f
C6 minus drain_left 0.171187f
C7 plus drain_left 2.68183f
C8 minus source 2.15959f
C9 plus source 2.17411f
C10 drain_right a_n1756_n2688# 6.12255f
C11 drain_left a_n1756_n2688# 6.39945f
C12 source a_n1756_n2688# 5.233246f
C13 minus a_n1756_n2688# 6.257572f
C14 plus a_n1756_n2688# 8.20316f
C15 drain_right.t0 a_n1756_n2688# 2.22136f
C16 drain_right.t12 a_n1756_n2688# 0.280749f
C17 drain_right.t7 a_n1756_n2688# 0.280749f
C18 drain_right.n0 a_n1756_n2688# 1.81162f
C19 drain_right.n1 a_n1756_n2688# 0.649859f
C20 drain_right.t11 a_n1756_n2688# 0.280749f
C21 drain_right.t5 a_n1756_n2688# 0.280749f
C22 drain_right.n2 a_n1756_n2688# 1.81427f
C23 drain_right.t1 a_n1756_n2688# 0.280749f
C24 drain_right.t13 a_n1756_n2688# 0.280749f
C25 drain_right.n3 a_n1756_n2688# 1.81162f
C26 drain_right.n4 a_n1756_n2688# 0.580587f
C27 drain_right.n5 a_n1756_n2688# 1.01997f
C28 drain_right.t10 a_n1756_n2688# 0.280749f
C29 drain_right.t9 a_n1756_n2688# 0.280749f
C30 drain_right.n6 a_n1756_n2688# 1.81427f
C31 drain_right.t6 a_n1756_n2688# 0.280749f
C32 drain_right.t4 a_n1756_n2688# 0.280749f
C33 drain_right.n7 a_n1756_n2688# 1.81162f
C34 drain_right.n8 a_n1756_n2688# 0.613386f
C35 drain_right.t2 a_n1756_n2688# 0.280749f
C36 drain_right.t8 a_n1756_n2688# 0.280749f
C37 drain_right.n9 a_n1756_n2688# 1.81162f
C38 drain_right.n10 a_n1756_n2688# 0.302771f
C39 drain_right.t3 a_n1756_n2688# 2.21842f
C40 drain_right.n11 a_n1756_n2688# 0.583243f
C41 minus.n0 a_n1756_n2688# 0.054626f
C42 minus.t10 a_n1756_n2688# 0.212747f
C43 minus.t11 a_n1756_n2688# 0.208964f
C44 minus.t5 a_n1756_n2688# 0.208964f
C45 minus.t7 a_n1756_n2688# 0.208964f
C46 minus.n1 a_n1756_n2688# 0.1138f
C47 minus.n2 a_n1756_n2688# 0.127689f
C48 minus.t9 a_n1756_n2688# 0.208964f
C49 minus.t3 a_n1756_n2688# 0.208964f
C50 minus.t4 a_n1756_n2688# 0.212747f
C51 minus.n3 a_n1756_n2688# 0.118522f
C52 minus.n4 a_n1756_n2688# 0.095679f
C53 minus.n5 a_n1756_n2688# 0.023173f
C54 minus.n6 a_n1756_n2688# 0.095679f
C55 minus.n7 a_n1756_n2688# 0.023173f
C56 minus.n8 a_n1756_n2688# 0.054626f
C57 minus.n9 a_n1756_n2688# 0.054626f
C58 minus.n10 a_n1756_n2688# 0.054626f
C59 minus.n11 a_n1756_n2688# 0.023173f
C60 minus.n12 a_n1756_n2688# 0.095679f
C61 minus.n13 a_n1756_n2688# 0.023173f
C62 minus.n14 a_n1756_n2688# 0.095679f
C63 minus.n15 a_n1756_n2688# 0.118437f
C64 minus.n16 a_n1756_n2688# 1.7161f
C65 minus.n17 a_n1756_n2688# 0.054626f
C66 minus.t2 a_n1756_n2688# 0.208964f
C67 minus.t0 a_n1756_n2688# 0.208964f
C68 minus.t12 a_n1756_n2688# 0.208964f
C69 minus.n18 a_n1756_n2688# 0.1138f
C70 minus.n19 a_n1756_n2688# 0.127689f
C71 minus.t6 a_n1756_n2688# 0.208964f
C72 minus.t1 a_n1756_n2688# 0.208964f
C73 minus.t13 a_n1756_n2688# 0.212747f
C74 minus.n20 a_n1756_n2688# 0.118522f
C75 minus.n21 a_n1756_n2688# 0.095679f
C76 minus.n22 a_n1756_n2688# 0.023173f
C77 minus.n23 a_n1756_n2688# 0.095679f
C78 minus.n24 a_n1756_n2688# 0.023173f
C79 minus.n25 a_n1756_n2688# 0.054626f
C80 minus.n26 a_n1756_n2688# 0.054626f
C81 minus.n27 a_n1756_n2688# 0.054626f
C82 minus.n28 a_n1756_n2688# 0.023173f
C83 minus.n29 a_n1756_n2688# 0.095679f
C84 minus.n30 a_n1756_n2688# 0.023173f
C85 minus.n31 a_n1756_n2688# 0.095679f
C86 minus.t8 a_n1756_n2688# 0.212747f
C87 minus.n32 a_n1756_n2688# 0.118437f
C88 minus.n33 a_n1756_n2688# 0.366181f
C89 minus.n34 a_n1756_n2688# 2.0965f
C90 drain_left.t12 a_n1756_n2688# 2.23018f
C91 drain_left.t1 a_n1756_n2688# 0.281864f
C92 drain_left.t9 a_n1756_n2688# 0.281864f
C93 drain_left.n0 a_n1756_n2688# 1.81881f
C94 drain_left.n1 a_n1756_n2688# 0.652439f
C95 drain_left.t8 a_n1756_n2688# 0.281864f
C96 drain_left.t10 a_n1756_n2688# 0.281864f
C97 drain_left.n2 a_n1756_n2688# 1.82148f
C98 drain_left.t11 a_n1756_n2688# 0.281864f
C99 drain_left.t13 a_n1756_n2688# 0.281864f
C100 drain_left.n3 a_n1756_n2688# 1.81881f
C101 drain_left.n4 a_n1756_n2688# 0.582892f
C102 drain_left.n5 a_n1756_n2688# 1.07795f
C103 drain_left.t7 a_n1756_n2688# 2.23018f
C104 drain_left.t2 a_n1756_n2688# 0.281864f
C105 drain_left.t4 a_n1756_n2688# 0.281864f
C106 drain_left.n6 a_n1756_n2688# 1.81881f
C107 drain_left.n7 a_n1756_n2688# 0.667242f
C108 drain_left.t6 a_n1756_n2688# 0.281864f
C109 drain_left.t0 a_n1756_n2688# 0.281864f
C110 drain_left.n8 a_n1756_n2688# 1.81881f
C111 drain_left.n9 a_n1756_n2688# 0.303973f
C112 drain_left.t3 a_n1756_n2688# 0.281864f
C113 drain_left.t5 a_n1756_n2688# 0.281864f
C114 drain_left.n10 a_n1756_n2688# 1.81881f
C115 drain_left.n11 a_n1756_n2688# 0.522418f
C116 source.t25 a_n1756_n2688# 2.21081f
C117 source.n0 a_n1756_n2688# 1.23323f
C118 source.t17 a_n1756_n2688# 0.292525f
C119 source.t14 a_n1756_n2688# 0.292525f
C120 source.n1 a_n1756_n2688# 1.81514f
C121 source.n2 a_n1756_n2688# 0.351036f
C122 source.t19 a_n1756_n2688# 0.292525f
C123 source.t26 a_n1756_n2688# 0.292525f
C124 source.n3 a_n1756_n2688# 1.81514f
C125 source.n4 a_n1756_n2688# 0.351036f
C126 source.t16 a_n1756_n2688# 0.292525f
C127 source.t20 a_n1756_n2688# 0.292525f
C128 source.n5 a_n1756_n2688# 1.81514f
C129 source.n6 a_n1756_n2688# 0.367626f
C130 source.t2 a_n1756_n2688# 2.21081f
C131 source.n7 a_n1756_n2688# 0.4985f
C132 source.t5 a_n1756_n2688# 0.292525f
C133 source.t11 a_n1756_n2688# 0.292525f
C134 source.n8 a_n1756_n2688# 1.81514f
C135 source.n9 a_n1756_n2688# 0.351036f
C136 source.t1 a_n1756_n2688# 0.292525f
C137 source.t4 a_n1756_n2688# 0.292525f
C138 source.n10 a_n1756_n2688# 1.81514f
C139 source.n11 a_n1756_n2688# 0.351036f
C140 source.t7 a_n1756_n2688# 0.292525f
C141 source.t9 a_n1756_n2688# 0.292525f
C142 source.n12 a_n1756_n2688# 1.81514f
C143 source.n13 a_n1756_n2688# 1.54629f
C144 source.t18 a_n1756_n2688# 0.292525f
C145 source.t22 a_n1756_n2688# 0.292525f
C146 source.n14 a_n1756_n2688# 1.81514f
C147 source.n15 a_n1756_n2688# 1.5463f
C148 source.t27 a_n1756_n2688# 0.292525f
C149 source.t15 a_n1756_n2688# 0.292525f
C150 source.n16 a_n1756_n2688# 1.81514f
C151 source.n17 a_n1756_n2688# 0.351041f
C152 source.t23 a_n1756_n2688# 0.292525f
C153 source.t21 a_n1756_n2688# 0.292525f
C154 source.n18 a_n1756_n2688# 1.81514f
C155 source.n19 a_n1756_n2688# 0.351041f
C156 source.t24 a_n1756_n2688# 2.21081f
C157 source.n20 a_n1756_n2688# 0.498505f
C158 source.t10 a_n1756_n2688# 0.292525f
C159 source.t8 a_n1756_n2688# 0.292525f
C160 source.n21 a_n1756_n2688# 1.81514f
C161 source.n22 a_n1756_n2688# 0.367631f
C162 source.t13 a_n1756_n2688# 0.292525f
C163 source.t3 a_n1756_n2688# 0.292525f
C164 source.n23 a_n1756_n2688# 1.81514f
C165 source.n24 a_n1756_n2688# 0.351041f
C166 source.t6 a_n1756_n2688# 0.292525f
C167 source.t0 a_n1756_n2688# 0.292525f
C168 source.n25 a_n1756_n2688# 1.81514f
C169 source.n26 a_n1756_n2688# 0.351041f
C170 source.t12 a_n1756_n2688# 2.21081f
C171 source.n27 a_n1756_n2688# 0.628443f
C172 source.n28 a_n1756_n2688# 1.41395f
C173 plus.n0 a_n1756_n2688# 0.056432f
C174 plus.t10 a_n1756_n2688# 0.215873f
C175 plus.t13 a_n1756_n2688# 0.215873f
C176 plus.t7 a_n1756_n2688# 0.215873f
C177 plus.n1 a_n1756_n2688# 0.117563f
C178 plus.n2 a_n1756_n2688# 0.131911f
C179 plus.t9 a_n1756_n2688# 0.215873f
C180 plus.t11 a_n1756_n2688# 0.215873f
C181 plus.t6 a_n1756_n2688# 0.219782f
C182 plus.n3 a_n1756_n2688# 0.122441f
C183 plus.n4 a_n1756_n2688# 0.098843f
C184 plus.n5 a_n1756_n2688# 0.023939f
C185 plus.n6 a_n1756_n2688# 0.098843f
C186 plus.n7 a_n1756_n2688# 0.023939f
C187 plus.n8 a_n1756_n2688# 0.056432f
C188 plus.n9 a_n1756_n2688# 0.056432f
C189 plus.n10 a_n1756_n2688# 0.056432f
C190 plus.n11 a_n1756_n2688# 0.023939f
C191 plus.n12 a_n1756_n2688# 0.098843f
C192 plus.n13 a_n1756_n2688# 0.023939f
C193 plus.n14 a_n1756_n2688# 0.098843f
C194 plus.t8 a_n1756_n2688# 0.219782f
C195 plus.n15 a_n1756_n2688# 0.122353f
C196 plus.n16 a_n1756_n2688# 0.563971f
C197 plus.n17 a_n1756_n2688# 0.056432f
C198 plus.t1 a_n1756_n2688# 0.219782f
C199 plus.t12 a_n1756_n2688# 0.215873f
C200 plus.t4 a_n1756_n2688# 0.215873f
C201 plus.t2 a_n1756_n2688# 0.215873f
C202 plus.n18 a_n1756_n2688# 0.117563f
C203 plus.n19 a_n1756_n2688# 0.131911f
C204 plus.t0 a_n1756_n2688# 0.215873f
C205 plus.t5 a_n1756_n2688# 0.215873f
C206 plus.t3 a_n1756_n2688# 0.219782f
C207 plus.n20 a_n1756_n2688# 0.122441f
C208 plus.n21 a_n1756_n2688# 0.098843f
C209 plus.n22 a_n1756_n2688# 0.023939f
C210 plus.n23 a_n1756_n2688# 0.098843f
C211 plus.n24 a_n1756_n2688# 0.023939f
C212 plus.n25 a_n1756_n2688# 0.056432f
C213 plus.n26 a_n1756_n2688# 0.056432f
C214 plus.n27 a_n1756_n2688# 0.056432f
C215 plus.n28 a_n1756_n2688# 0.023939f
C216 plus.n29 a_n1756_n2688# 0.098843f
C217 plus.n30 a_n1756_n2688# 0.023939f
C218 plus.n31 a_n1756_n2688# 0.098843f
C219 plus.n32 a_n1756_n2688# 0.122353f
C220 plus.n33 a_n1756_n2688# 1.54665f
.ends

