* NGSPICE file created from diffpair226.ext - technology: sky130A

.subckt diffpair226 minus drain_right drain_left source plus
X0 source.t24 minus.t0 drain_right.t4 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X1 drain_right.t11 minus.t1 source.t23 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X2 a_n2364_n1488# a_n2364_n1488# a_n2364_n1488# a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.7
X3 drain_left.t13 plus.t0 source.t6 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X4 drain_left.t12 plus.t1 source.t7 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X5 source.t22 minus.t2 drain_right.t1 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X6 a_n2364_n1488# a_n2364_n1488# a_n2364_n1488# a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X7 drain_left.t11 plus.t2 source.t0 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X8 drain_left.t10 plus.t3 source.t1 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X9 source.t21 minus.t3 drain_right.t8 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X10 drain_right.t0 minus.t4 source.t20 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X11 drain_right.t2 minus.t5 source.t19 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X12 drain_left.t9 plus.t4 source.t2 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X13 source.t9 plus.t5 drain_left.t8 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X14 a_n2364_n1488# a_n2364_n1488# a_n2364_n1488# a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X15 drain_right.t12 minus.t6 source.t18 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X16 drain_right.t9 minus.t7 source.t17 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X17 drain_right.t13 minus.t8 source.t16 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X18 source.t15 minus.t9 drain_right.t5 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X19 drain_left.t7 plus.t6 source.t25 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X20 drain_right.t6 minus.t10 source.t14 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X21 source.t26 plus.t7 drain_left.t6 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X22 source.t5 plus.t8 drain_left.t5 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X23 drain_right.t7 minus.t11 source.t13 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X24 a_n2364_n1488# a_n2364_n1488# a_n2364_n1488# a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X25 source.t4 plus.t9 drain_left.t4 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X26 drain_left.t3 plus.t10 source.t10 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X27 source.t3 plus.t11 drain_left.t2 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X28 drain_left.t1 plus.t12 source.t8 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X29 source.t12 minus.t12 drain_right.t3 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X30 source.t11 minus.t13 drain_right.t10 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X31 source.t27 plus.t13 drain_left.t0 a_n2364_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
R0 minus.n5 minus.t11 183.251
R1 minus.n27 minus.t1 183.251
R2 minus.n21 minus.n20 161.3
R3 minus.n19 minus.n0 161.3
R4 minus.n18 minus.n17 161.3
R5 minus.n16 minus.n1 161.3
R6 minus.n15 minus.n14 161.3
R7 minus.n13 minus.n2 161.3
R8 minus.n12 minus.n11 161.3
R9 minus.n10 minus.n3 161.3
R10 minus.n9 minus.n8 161.3
R11 minus.n7 minus.n4 161.3
R12 minus.n43 minus.n42 161.3
R13 minus.n41 minus.n22 161.3
R14 minus.n40 minus.n39 161.3
R15 minus.n38 minus.n23 161.3
R16 minus.n37 minus.n36 161.3
R17 minus.n35 minus.n24 161.3
R18 minus.n34 minus.n33 161.3
R19 minus.n32 minus.n25 161.3
R20 minus.n31 minus.n30 161.3
R21 minus.n29 minus.n26 161.3
R22 minus.n6 minus.t2 159.405
R23 minus.n8 minus.t10 159.405
R24 minus.n12 minus.t12 159.405
R25 minus.n14 minus.t7 159.405
R26 minus.n18 minus.t13 159.405
R27 minus.n20 minus.t6 159.405
R28 minus.n28 minus.t0 159.405
R29 minus.n30 minus.t4 159.405
R30 minus.n34 minus.t3 159.405
R31 minus.n36 minus.t5 159.405
R32 minus.n40 minus.t9 159.405
R33 minus.n42 minus.t8 159.405
R34 minus.n5 minus.n4 44.9119
R35 minus.n27 minus.n26 44.9119
R36 minus.n20 minus.n19 35.055
R37 minus.n42 minus.n41 35.055
R38 minus.n44 minus.n21 31.4077
R39 minus.n7 minus.n6 30.6732
R40 minus.n18 minus.n1 30.6732
R41 minus.n29 minus.n28 30.6732
R42 minus.n40 minus.n23 30.6732
R43 minus.n8 minus.n3 26.2914
R44 minus.n14 minus.n13 26.2914
R45 minus.n30 minus.n25 26.2914
R46 minus.n36 minus.n35 26.2914
R47 minus.n12 minus.n3 21.9096
R48 minus.n13 minus.n12 21.9096
R49 minus.n34 minus.n25 21.9096
R50 minus.n35 minus.n34 21.9096
R51 minus.n6 minus.n5 17.739
R52 minus.n28 minus.n27 17.739
R53 minus.n8 minus.n7 17.5278
R54 minus.n14 minus.n1 17.5278
R55 minus.n30 minus.n29 17.5278
R56 minus.n36 minus.n23 17.5278
R57 minus.n19 minus.n18 13.146
R58 minus.n41 minus.n40 13.146
R59 minus.n44 minus.n43 6.65012
R60 minus.n21 minus.n0 0.189894
R61 minus.n17 minus.n0 0.189894
R62 minus.n17 minus.n16 0.189894
R63 minus.n16 minus.n15 0.189894
R64 minus.n15 minus.n2 0.189894
R65 minus.n11 minus.n2 0.189894
R66 minus.n11 minus.n10 0.189894
R67 minus.n10 minus.n9 0.189894
R68 minus.n9 minus.n4 0.189894
R69 minus.n31 minus.n26 0.189894
R70 minus.n32 minus.n31 0.189894
R71 minus.n33 minus.n32 0.189894
R72 minus.n33 minus.n24 0.189894
R73 minus.n37 minus.n24 0.189894
R74 minus.n38 minus.n37 0.189894
R75 minus.n39 minus.n38 0.189894
R76 minus.n39 minus.n22 0.189894
R77 minus.n43 minus.n22 0.189894
R78 minus minus.n44 0.188
R79 drain_right.n1 drain_right.t11 87.2609
R80 drain_right.n11 drain_right.t12 86.3731
R81 drain_right.n8 drain_right.n6 80.661
R82 drain_right.n4 drain_right.n2 80.6609
R83 drain_right.n8 drain_right.n7 79.7731
R84 drain_right.n10 drain_right.n9 79.7731
R85 drain_right.n4 drain_right.n3 79.773
R86 drain_right.n1 drain_right.n0 79.773
R87 drain_right drain_right.n5 25.1013
R88 drain_right.n2 drain_right.t5 6.6005
R89 drain_right.n2 drain_right.t13 6.6005
R90 drain_right.n3 drain_right.t8 6.6005
R91 drain_right.n3 drain_right.t2 6.6005
R92 drain_right.n0 drain_right.t4 6.6005
R93 drain_right.n0 drain_right.t0 6.6005
R94 drain_right.n6 drain_right.t1 6.6005
R95 drain_right.n6 drain_right.t7 6.6005
R96 drain_right.n7 drain_right.t3 6.6005
R97 drain_right.n7 drain_right.t6 6.6005
R98 drain_right.n9 drain_right.t10 6.6005
R99 drain_right.n9 drain_right.t9 6.6005
R100 drain_right drain_right.n11 6.09718
R101 drain_right.n11 drain_right.n10 0.888431
R102 drain_right.n10 drain_right.n8 0.888431
R103 drain_right.n5 drain_right.n1 0.611102
R104 drain_right.n5 drain_right.n4 0.167137
R105 source.n0 source.t6 69.6943
R106 source.n7 source.t13 69.6943
R107 source.n27 source.t16 69.6942
R108 source.n20 source.t2 69.6942
R109 source.n2 source.n1 63.0943
R110 source.n4 source.n3 63.0943
R111 source.n6 source.n5 63.0943
R112 source.n9 source.n8 63.0943
R113 source.n11 source.n10 63.0943
R114 source.n13 source.n12 63.0943
R115 source.n26 source.n25 63.0942
R116 source.n24 source.n23 63.0942
R117 source.n22 source.n21 63.0942
R118 source.n19 source.n18 63.0942
R119 source.n17 source.n16 63.0942
R120 source.n15 source.n14 63.0942
R121 source.n15 source.n13 16.2454
R122 source.n28 source.n0 9.65058
R123 source.n25 source.t19 6.6005
R124 source.n25 source.t15 6.6005
R125 source.n23 source.t20 6.6005
R126 source.n23 source.t21 6.6005
R127 source.n21 source.t23 6.6005
R128 source.n21 source.t24 6.6005
R129 source.n18 source.t25 6.6005
R130 source.n18 source.t9 6.6005
R131 source.n16 source.t10 6.6005
R132 source.n16 source.t3 6.6005
R133 source.n14 source.t8 6.6005
R134 source.n14 source.t27 6.6005
R135 source.n1 source.t0 6.6005
R136 source.n1 source.t5 6.6005
R137 source.n3 source.t7 6.6005
R138 source.n3 source.t26 6.6005
R139 source.n5 source.t1 6.6005
R140 source.n5 source.t4 6.6005
R141 source.n8 source.t14 6.6005
R142 source.n8 source.t22 6.6005
R143 source.n10 source.t17 6.6005
R144 source.n10 source.t12 6.6005
R145 source.n12 source.t18 6.6005
R146 source.n12 source.t11 6.6005
R147 source.n28 source.n27 5.7074
R148 source.n7 source.n6 0.914293
R149 source.n22 source.n20 0.914293
R150 source.n13 source.n11 0.888431
R151 source.n11 source.n9 0.888431
R152 source.n9 source.n7 0.888431
R153 source.n6 source.n4 0.888431
R154 source.n4 source.n2 0.888431
R155 source.n2 source.n0 0.888431
R156 source.n17 source.n15 0.888431
R157 source.n19 source.n17 0.888431
R158 source.n20 source.n19 0.888431
R159 source.n24 source.n22 0.888431
R160 source.n26 source.n24 0.888431
R161 source.n27 source.n26 0.888431
R162 source source.n28 0.188
R163 plus.n5 plus.t3 183.251
R164 plus.n27 plus.t4 183.251
R165 plus.n8 plus.n7 161.3
R166 plus.n9 plus.n4 161.3
R167 plus.n11 plus.n10 161.3
R168 plus.n12 plus.n3 161.3
R169 plus.n14 plus.n13 161.3
R170 plus.n15 plus.n2 161.3
R171 plus.n17 plus.n16 161.3
R172 plus.n18 plus.n1 161.3
R173 plus.n19 plus.n0 161.3
R174 plus.n21 plus.n20 161.3
R175 plus.n30 plus.n29 161.3
R176 plus.n31 plus.n26 161.3
R177 plus.n33 plus.n32 161.3
R178 plus.n34 plus.n25 161.3
R179 plus.n36 plus.n35 161.3
R180 plus.n37 plus.n24 161.3
R181 plus.n39 plus.n38 161.3
R182 plus.n40 plus.n23 161.3
R183 plus.n41 plus.n22 161.3
R184 plus.n43 plus.n42 161.3
R185 plus.n20 plus.t0 159.405
R186 plus.n18 plus.t8 159.405
R187 plus.n2 plus.t2 159.405
R188 plus.n12 plus.t7 159.405
R189 plus.n4 plus.t1 159.405
R190 plus.n6 plus.t9 159.405
R191 plus.n42 plus.t12 159.405
R192 plus.n40 plus.t13 159.405
R193 plus.n24 plus.t10 159.405
R194 plus.n34 plus.t11 159.405
R195 plus.n26 plus.t6 159.405
R196 plus.n28 plus.t5 159.405
R197 plus.n30 plus.n27 44.9119
R198 plus.n8 plus.n5 44.9119
R199 plus.n20 plus.n19 35.055
R200 plus.n42 plus.n41 35.055
R201 plus.n18 plus.n17 30.6732
R202 plus.n7 plus.n6 30.6732
R203 plus.n40 plus.n39 30.6732
R204 plus.n29 plus.n28 30.6732
R205 plus plus.n43 28.6979
R206 plus.n13 plus.n2 26.2914
R207 plus.n11 plus.n4 26.2914
R208 plus.n35 plus.n24 26.2914
R209 plus.n33 plus.n26 26.2914
R210 plus.n13 plus.n12 21.9096
R211 plus.n12 plus.n11 21.9096
R212 plus.n35 plus.n34 21.9096
R213 plus.n34 plus.n33 21.9096
R214 plus.n28 plus.n27 17.739
R215 plus.n6 plus.n5 17.739
R216 plus.n17 plus.n2 17.5278
R217 plus.n7 plus.n4 17.5278
R218 plus.n39 plus.n24 17.5278
R219 plus.n29 plus.n26 17.5278
R220 plus.n19 plus.n18 13.146
R221 plus.n41 plus.n40 13.146
R222 plus plus.n21 8.88497
R223 plus.n9 plus.n8 0.189894
R224 plus.n10 plus.n9 0.189894
R225 plus.n10 plus.n3 0.189894
R226 plus.n14 plus.n3 0.189894
R227 plus.n15 plus.n14 0.189894
R228 plus.n16 plus.n15 0.189894
R229 plus.n16 plus.n1 0.189894
R230 plus.n1 plus.n0 0.189894
R231 plus.n21 plus.n0 0.189894
R232 plus.n43 plus.n22 0.189894
R233 plus.n23 plus.n22 0.189894
R234 plus.n38 plus.n23 0.189894
R235 plus.n38 plus.n37 0.189894
R236 plus.n37 plus.n36 0.189894
R237 plus.n36 plus.n25 0.189894
R238 plus.n32 plus.n25 0.189894
R239 plus.n32 plus.n31 0.189894
R240 plus.n31 plus.n30 0.189894
R241 drain_left.n7 drain_left.t10 87.261
R242 drain_left.n1 drain_left.t1 87.2609
R243 drain_left.n4 drain_left.n2 80.6609
R244 drain_left.n11 drain_left.n10 79.7731
R245 drain_left.n9 drain_left.n8 79.7731
R246 drain_left.n7 drain_left.n6 79.7731
R247 drain_left.n4 drain_left.n3 79.773
R248 drain_left.n1 drain_left.n0 79.773
R249 drain_left drain_left.n5 25.6545
R250 drain_left.n2 drain_left.t8 6.6005
R251 drain_left.n2 drain_left.t9 6.6005
R252 drain_left.n3 drain_left.t2 6.6005
R253 drain_left.n3 drain_left.t7 6.6005
R254 drain_left.n0 drain_left.t0 6.6005
R255 drain_left.n0 drain_left.t3 6.6005
R256 drain_left.n10 drain_left.t5 6.6005
R257 drain_left.n10 drain_left.t13 6.6005
R258 drain_left.n8 drain_left.t6 6.6005
R259 drain_left.n8 drain_left.t11 6.6005
R260 drain_left.n6 drain_left.t4 6.6005
R261 drain_left.n6 drain_left.t12 6.6005
R262 drain_left drain_left.n11 6.54115
R263 drain_left.n9 drain_left.n7 0.888431
R264 drain_left.n11 drain_left.n9 0.888431
R265 drain_left.n5 drain_left.n1 0.611102
R266 drain_left.n5 drain_left.n4 0.167137
C0 plus drain_right 0.395426f
C1 plus source 3.13274f
C2 minus drain_right 2.67553f
C3 minus source 3.11862f
C4 drain_left drain_right 1.23103f
C5 drain_left source 7.07413f
C6 plus minus 4.43246f
C7 drain_right source 7.07353f
C8 drain_left plus 2.90806f
C9 drain_left minus 0.17789f
C10 drain_right a_n2364_n1488# 5.00421f
C11 drain_left a_n2364_n1488# 5.36517f
C12 source a_n2364_n1488# 3.164833f
C13 minus a_n2364_n1488# 8.637661f
C14 plus a_n2364_n1488# 9.93221f
C15 drain_left.t1 a_n2364_n1488# 0.563271f
C16 drain_left.t0 a_n2364_n1488# 0.060493f
C17 drain_left.t3 a_n2364_n1488# 0.060493f
C18 drain_left.n0 a_n2364_n1488# 0.436266f
C19 drain_left.n1 a_n2364_n1488# 0.653955f
C20 drain_left.t8 a_n2364_n1488# 0.060493f
C21 drain_left.t9 a_n2364_n1488# 0.060493f
C22 drain_left.n2 a_n2364_n1488# 0.440235f
C23 drain_left.t2 a_n2364_n1488# 0.060493f
C24 drain_left.t7 a_n2364_n1488# 0.060493f
C25 drain_left.n3 a_n2364_n1488# 0.436266f
C26 drain_left.n4 a_n2364_n1488# 0.651096f
C27 drain_left.n5 a_n2364_n1488# 0.926473f
C28 drain_left.t10 a_n2364_n1488# 0.563273f
C29 drain_left.t4 a_n2364_n1488# 0.060493f
C30 drain_left.t12 a_n2364_n1488# 0.060493f
C31 drain_left.n6 a_n2364_n1488# 0.436268f
C32 drain_left.n7 a_n2364_n1488# 0.675784f
C33 drain_left.t6 a_n2364_n1488# 0.060493f
C34 drain_left.t11 a_n2364_n1488# 0.060493f
C35 drain_left.n8 a_n2364_n1488# 0.436268f
C36 drain_left.n9 a_n2364_n1488# 0.350269f
C37 drain_left.t5 a_n2364_n1488# 0.060493f
C38 drain_left.t13 a_n2364_n1488# 0.060493f
C39 drain_left.n10 a_n2364_n1488# 0.436268f
C40 drain_left.n11 a_n2364_n1488# 0.575967f
C41 plus.n0 a_n2364_n1488# 0.044274f
C42 plus.t0 a_n2364_n1488# 0.2788f
C43 plus.t8 a_n2364_n1488# 0.2788f
C44 plus.n1 a_n2364_n1488# 0.044274f
C45 plus.t2 a_n2364_n1488# 0.2788f
C46 plus.n2 a_n2364_n1488# 0.162379f
C47 plus.n3 a_n2364_n1488# 0.044274f
C48 plus.t7 a_n2364_n1488# 0.2788f
C49 plus.t1 a_n2364_n1488# 0.2788f
C50 plus.n4 a_n2364_n1488# 0.162379f
C51 plus.t3 a_n2364_n1488# 0.299936f
C52 plus.n5 a_n2364_n1488# 0.14509f
C53 plus.t9 a_n2364_n1488# 0.2788f
C54 plus.n6 a_n2364_n1488# 0.167864f
C55 plus.n7 a_n2364_n1488# 0.010047f
C56 plus.n8 a_n2364_n1488# 0.186545f
C57 plus.n9 a_n2364_n1488# 0.044274f
C58 plus.n10 a_n2364_n1488# 0.044274f
C59 plus.n11 a_n2364_n1488# 0.010047f
C60 plus.n12 a_n2364_n1488# 0.162379f
C61 plus.n13 a_n2364_n1488# 0.010047f
C62 plus.n14 a_n2364_n1488# 0.044274f
C63 plus.n15 a_n2364_n1488# 0.044274f
C64 plus.n16 a_n2364_n1488# 0.044274f
C65 plus.n17 a_n2364_n1488# 0.010047f
C66 plus.n18 a_n2364_n1488# 0.162379f
C67 plus.n19 a_n2364_n1488# 0.010047f
C68 plus.n20 a_n2364_n1488# 0.160742f
C69 plus.n21 a_n2364_n1488# 0.347105f
C70 plus.n22 a_n2364_n1488# 0.044274f
C71 plus.t12 a_n2364_n1488# 0.2788f
C72 plus.n23 a_n2364_n1488# 0.044274f
C73 plus.t13 a_n2364_n1488# 0.2788f
C74 plus.t10 a_n2364_n1488# 0.2788f
C75 plus.n24 a_n2364_n1488# 0.162379f
C76 plus.n25 a_n2364_n1488# 0.044274f
C77 plus.t11 a_n2364_n1488# 0.2788f
C78 plus.t6 a_n2364_n1488# 0.2788f
C79 plus.n26 a_n2364_n1488# 0.162379f
C80 plus.t4 a_n2364_n1488# 0.299936f
C81 plus.n27 a_n2364_n1488# 0.14509f
C82 plus.t5 a_n2364_n1488# 0.2788f
C83 plus.n28 a_n2364_n1488# 0.167864f
C84 plus.n29 a_n2364_n1488# 0.010047f
C85 plus.n30 a_n2364_n1488# 0.186545f
C86 plus.n31 a_n2364_n1488# 0.044274f
C87 plus.n32 a_n2364_n1488# 0.044274f
C88 plus.n33 a_n2364_n1488# 0.010047f
C89 plus.n34 a_n2364_n1488# 0.162379f
C90 plus.n35 a_n2364_n1488# 0.010047f
C91 plus.n36 a_n2364_n1488# 0.044274f
C92 plus.n37 a_n2364_n1488# 0.044274f
C93 plus.n38 a_n2364_n1488# 0.044274f
C94 plus.n39 a_n2364_n1488# 0.010047f
C95 plus.n40 a_n2364_n1488# 0.162379f
C96 plus.n41 a_n2364_n1488# 0.010047f
C97 plus.n42 a_n2364_n1488# 0.160742f
C98 plus.n43 a_n2364_n1488# 1.17446f
C99 source.t6 a_n2364_n1488# 0.612473f
C100 source.n0 a_n2364_n1488# 0.896341f
C101 source.t0 a_n2364_n1488# 0.073758f
C102 source.t5 a_n2364_n1488# 0.073758f
C103 source.n1 a_n2364_n1488# 0.467668f
C104 source.n2 a_n2364_n1488# 0.449062f
C105 source.t7 a_n2364_n1488# 0.073758f
C106 source.t26 a_n2364_n1488# 0.073758f
C107 source.n3 a_n2364_n1488# 0.467668f
C108 source.n4 a_n2364_n1488# 0.449062f
C109 source.t1 a_n2364_n1488# 0.073758f
C110 source.t4 a_n2364_n1488# 0.073758f
C111 source.n5 a_n2364_n1488# 0.467668f
C112 source.n6 a_n2364_n1488# 0.451655f
C113 source.t13 a_n2364_n1488# 0.612473f
C114 source.n7 a_n2364_n1488# 0.508007f
C115 source.t14 a_n2364_n1488# 0.073758f
C116 source.t22 a_n2364_n1488# 0.073758f
C117 source.n8 a_n2364_n1488# 0.467668f
C118 source.n9 a_n2364_n1488# 0.449062f
C119 source.t17 a_n2364_n1488# 0.073758f
C120 source.t12 a_n2364_n1488# 0.073758f
C121 source.n10 a_n2364_n1488# 0.467668f
C122 source.n11 a_n2364_n1488# 0.449062f
C123 source.t18 a_n2364_n1488# 0.073758f
C124 source.t11 a_n2364_n1488# 0.073758f
C125 source.n12 a_n2364_n1488# 0.467668f
C126 source.n13 a_n2364_n1488# 1.26173f
C127 source.t8 a_n2364_n1488# 0.073758f
C128 source.t27 a_n2364_n1488# 0.073758f
C129 source.n14 a_n2364_n1488# 0.467665f
C130 source.n15 a_n2364_n1488# 1.26173f
C131 source.t10 a_n2364_n1488# 0.073758f
C132 source.t3 a_n2364_n1488# 0.073758f
C133 source.n16 a_n2364_n1488# 0.467665f
C134 source.n17 a_n2364_n1488# 0.449065f
C135 source.t25 a_n2364_n1488# 0.073758f
C136 source.t9 a_n2364_n1488# 0.073758f
C137 source.n18 a_n2364_n1488# 0.467665f
C138 source.n19 a_n2364_n1488# 0.449065f
C139 source.t2 a_n2364_n1488# 0.61247f
C140 source.n20 a_n2364_n1488# 0.508011f
C141 source.t23 a_n2364_n1488# 0.073758f
C142 source.t24 a_n2364_n1488# 0.073758f
C143 source.n21 a_n2364_n1488# 0.467665f
C144 source.n22 a_n2364_n1488# 0.451658f
C145 source.t20 a_n2364_n1488# 0.073758f
C146 source.t21 a_n2364_n1488# 0.073758f
C147 source.n23 a_n2364_n1488# 0.467665f
C148 source.n24 a_n2364_n1488# 0.449065f
C149 source.t19 a_n2364_n1488# 0.073758f
C150 source.t15 a_n2364_n1488# 0.073758f
C151 source.n25 a_n2364_n1488# 0.467665f
C152 source.n26 a_n2364_n1488# 0.449065f
C153 source.t16 a_n2364_n1488# 0.61247f
C154 source.n27 a_n2364_n1488# 0.66645f
C155 source.n28 a_n2364_n1488# 0.917467f
C156 drain_right.t11 a_n2364_n1488# 0.557571f
C157 drain_right.t4 a_n2364_n1488# 0.05988f
C158 drain_right.t0 a_n2364_n1488# 0.05988f
C159 drain_right.n0 a_n2364_n1488# 0.431851f
C160 drain_right.n1 a_n2364_n1488# 0.647337f
C161 drain_right.t5 a_n2364_n1488# 0.05988f
C162 drain_right.t13 a_n2364_n1488# 0.05988f
C163 drain_right.n2 a_n2364_n1488# 0.43578f
C164 drain_right.t8 a_n2364_n1488# 0.05988f
C165 drain_right.t2 a_n2364_n1488# 0.05988f
C166 drain_right.n3 a_n2364_n1488# 0.431851f
C167 drain_right.n4 a_n2364_n1488# 0.644507f
C168 drain_right.n5 a_n2364_n1488# 0.867353f
C169 drain_right.t1 a_n2364_n1488# 0.05988f
C170 drain_right.t7 a_n2364_n1488# 0.05988f
C171 drain_right.n6 a_n2364_n1488# 0.435782f
C172 drain_right.t3 a_n2364_n1488# 0.05988f
C173 drain_right.t6 a_n2364_n1488# 0.05988f
C174 drain_right.n7 a_n2364_n1488# 0.431853f
C175 drain_right.n8 a_n2364_n1488# 0.699694f
C176 drain_right.t10 a_n2364_n1488# 0.05988f
C177 drain_right.t9 a_n2364_n1488# 0.05988f
C178 drain_right.n9 a_n2364_n1488# 0.431853f
C179 drain_right.n10 a_n2364_n1488# 0.346725f
C180 drain_right.t12 a_n2364_n1488# 0.554261f
C181 drain_right.n11 a_n2364_n1488# 0.557674f
C182 minus.n0 a_n2364_n1488# 0.043052f
C183 minus.n1 a_n2364_n1488# 0.009769f
C184 minus.t13 a_n2364_n1488# 0.271104f
C185 minus.n2 a_n2364_n1488# 0.043052f
C186 minus.n3 a_n2364_n1488# 0.009769f
C187 minus.t12 a_n2364_n1488# 0.271104f
C188 minus.n4 a_n2364_n1488# 0.181396f
C189 minus.t11 a_n2364_n1488# 0.291657f
C190 minus.n5 a_n2364_n1488# 0.141086f
C191 minus.t2 a_n2364_n1488# 0.271104f
C192 minus.n6 a_n2364_n1488# 0.16323f
C193 minus.n7 a_n2364_n1488# 0.009769f
C194 minus.t10 a_n2364_n1488# 0.271104f
C195 minus.n8 a_n2364_n1488# 0.157897f
C196 minus.n9 a_n2364_n1488# 0.043052f
C197 minus.n10 a_n2364_n1488# 0.043052f
C198 minus.n11 a_n2364_n1488# 0.043052f
C199 minus.n12 a_n2364_n1488# 0.157897f
C200 minus.n13 a_n2364_n1488# 0.009769f
C201 minus.t7 a_n2364_n1488# 0.271104f
C202 minus.n14 a_n2364_n1488# 0.157897f
C203 minus.n15 a_n2364_n1488# 0.043052f
C204 minus.n16 a_n2364_n1488# 0.043052f
C205 minus.n17 a_n2364_n1488# 0.043052f
C206 minus.n18 a_n2364_n1488# 0.157897f
C207 minus.n19 a_n2364_n1488# 0.009769f
C208 minus.t6 a_n2364_n1488# 0.271104f
C209 minus.n20 a_n2364_n1488# 0.156305f
C210 minus.n21 a_n2364_n1488# 1.21584f
C211 minus.n22 a_n2364_n1488# 0.043052f
C212 minus.n23 a_n2364_n1488# 0.009769f
C213 minus.n24 a_n2364_n1488# 0.043052f
C214 minus.n25 a_n2364_n1488# 0.009769f
C215 minus.n26 a_n2364_n1488# 0.181396f
C216 minus.t1 a_n2364_n1488# 0.291657f
C217 minus.n27 a_n2364_n1488# 0.141086f
C218 minus.t0 a_n2364_n1488# 0.271104f
C219 minus.n28 a_n2364_n1488# 0.16323f
C220 minus.n29 a_n2364_n1488# 0.009769f
C221 minus.t4 a_n2364_n1488# 0.271104f
C222 minus.n30 a_n2364_n1488# 0.157897f
C223 minus.n31 a_n2364_n1488# 0.043052f
C224 minus.n32 a_n2364_n1488# 0.043052f
C225 minus.n33 a_n2364_n1488# 0.043052f
C226 minus.t3 a_n2364_n1488# 0.271104f
C227 minus.n34 a_n2364_n1488# 0.157897f
C228 minus.n35 a_n2364_n1488# 0.009769f
C229 minus.t5 a_n2364_n1488# 0.271104f
C230 minus.n36 a_n2364_n1488# 0.157897f
C231 minus.n37 a_n2364_n1488# 0.043052f
C232 minus.n38 a_n2364_n1488# 0.043052f
C233 minus.n39 a_n2364_n1488# 0.043052f
C234 minus.t9 a_n2364_n1488# 0.271104f
C235 minus.n40 a_n2364_n1488# 0.157897f
C236 minus.n41 a_n2364_n1488# 0.009769f
C237 minus.t8 a_n2364_n1488# 0.271104f
C238 minus.n42 a_n2364_n1488# 0.156305f
C239 minus.n43 a_n2364_n1488# 0.296582f
C240 minus.n44 a_n2364_n1488# 1.489f
.ends

