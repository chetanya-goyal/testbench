* NGSPICE file created from diffpair95.ext - technology: sky130A

.subckt diffpair95 minus drain_right drain_left source plus
X0 source.t23 minus.t0 drain_right.t7 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X1 drain_right.t2 minus.t1 source.t22 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X2 source.t6 plus.t0 drain_left.t11 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X3 drain_right.t4 minus.t2 source.t21 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X4 source.t0 plus.t1 drain_left.t10 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X5 a_n1458_n1288# a_n1458_n1288# a_n1458_n1288# a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.2
X6 drain_left.t9 plus.t2 source.t9 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X7 drain_left.t8 plus.t3 source.t1 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X8 source.t20 minus.t3 drain_right.t10 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X9 source.t19 minus.t4 drain_right.t3 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X10 a_n1458_n1288# a_n1458_n1288# a_n1458_n1288# a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X11 drain_left.t7 plus.t4 source.t4 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X12 source.t2 plus.t5 drain_left.t6 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X13 drain_right.t9 minus.t5 source.t18 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X14 source.t17 minus.t6 drain_right.t5 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X15 drain_left.t5 plus.t6 source.t8 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X16 drain_right.t0 minus.t7 source.t16 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X17 drain_right.t11 minus.t8 source.t15 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X18 a_n1458_n1288# a_n1458_n1288# a_n1458_n1288# a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X19 a_n1458_n1288# a_n1458_n1288# a_n1458_n1288# a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X20 source.t11 plus.t7 drain_left.t4 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X21 drain_left.t3 plus.t8 source.t10 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X22 drain_right.t6 minus.t9 source.t14 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X23 source.t3 plus.t9 drain_left.t2 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X24 source.t13 minus.t10 drain_right.t1 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X25 source.t12 minus.t11 drain_right.t8 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X26 drain_left.t1 plus.t10 source.t5 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X27 source.t7 plus.t11 drain_left.t0 a_n1458_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
R0 minus.n11 minus.t3 445.12
R1 minus.n2 minus.t7 445.12
R2 minus.n24 minus.t5 445.12
R3 minus.n15 minus.t11 445.12
R4 minus.n10 minus.t8 397.651
R5 minus.n8 minus.t10 397.651
R6 minus.n1 minus.t2 397.651
R7 minus.n3 minus.t4 397.651
R8 minus.n23 minus.t0 397.651
R9 minus.n21 minus.t9 397.651
R10 minus.n14 minus.t6 397.651
R11 minus.n16 minus.t1 397.651
R12 minus.n5 minus.n2 161.489
R13 minus.n18 minus.n15 161.489
R14 minus.n12 minus.n11 161.3
R15 minus.n9 minus.n0 161.3
R16 minus.n7 minus.n6 161.3
R17 minus.n5 minus.n4 161.3
R18 minus.n25 minus.n24 161.3
R19 minus.n22 minus.n13 161.3
R20 minus.n20 minus.n19 161.3
R21 minus.n18 minus.n17 161.3
R22 minus.n10 minus.n9 43.0884
R23 minus.n4 minus.n3 43.0884
R24 minus.n17 minus.n16 43.0884
R25 minus.n23 minus.n22 43.0884
R26 minus.n8 minus.n7 38.7066
R27 minus.n7 minus.n1 38.7066
R28 minus.n20 minus.n14 38.7066
R29 minus.n21 minus.n20 38.7066
R30 minus.n9 minus.n8 34.3247
R31 minus.n4 minus.n1 34.3247
R32 minus.n17 minus.n14 34.3247
R33 minus.n22 minus.n21 34.3247
R34 minus.n11 minus.n10 29.9429
R35 minus.n3 minus.n2 29.9429
R36 minus.n16 minus.n15 29.9429
R37 minus.n24 minus.n23 29.9429
R38 minus.n26 minus.n12 27.0232
R39 minus.n26 minus.n25 6.45505
R40 minus.n12 minus.n0 0.189894
R41 minus.n6 minus.n0 0.189894
R42 minus.n6 minus.n5 0.189894
R43 minus.n19 minus.n18 0.189894
R44 minus.n19 minus.n13 0.189894
R45 minus.n25 minus.n13 0.189894
R46 minus minus.n26 0.188
R47 drain_right.n6 drain_right.n4 101.252
R48 drain_right.n3 drain_right.n2 101.198
R49 drain_right.n3 drain_right.n0 101.198
R50 drain_right.n6 drain_right.n5 100.796
R51 drain_right.n8 drain_right.n7 100.796
R52 drain_right.n3 drain_right.n1 100.796
R53 drain_right drain_right.n3 21.5226
R54 drain_right.n1 drain_right.t5 9.9005
R55 drain_right.n1 drain_right.t6 9.9005
R56 drain_right.n2 drain_right.t7 9.9005
R57 drain_right.n2 drain_right.t9 9.9005
R58 drain_right.n0 drain_right.t8 9.9005
R59 drain_right.n0 drain_right.t2 9.9005
R60 drain_right.n4 drain_right.t3 9.9005
R61 drain_right.n4 drain_right.t0 9.9005
R62 drain_right.n5 drain_right.t1 9.9005
R63 drain_right.n5 drain_right.t4 9.9005
R64 drain_right.n7 drain_right.t10 9.9005
R65 drain_right.n7 drain_right.t11 9.9005
R66 drain_right drain_right.n8 6.11011
R67 drain_right.n8 drain_right.n6 0.457397
R68 source.n74 source.n72 289.615
R69 source.n62 source.n60 289.615
R70 source.n54 source.n52 289.615
R71 source.n42 source.n40 289.615
R72 source.n2 source.n0 289.615
R73 source.n14 source.n12 289.615
R74 source.n22 source.n20 289.615
R75 source.n34 source.n32 289.615
R76 source.n75 source.n74 185
R77 source.n63 source.n62 185
R78 source.n55 source.n54 185
R79 source.n43 source.n42 185
R80 source.n3 source.n2 185
R81 source.n15 source.n14 185
R82 source.n23 source.n22 185
R83 source.n35 source.n34 185
R84 source.t18 source.n73 167.117
R85 source.t12 source.n61 167.117
R86 source.t5 source.n53 167.117
R87 source.t3 source.n41 167.117
R88 source.t4 source.n1 167.117
R89 source.t2 source.n13 167.117
R90 source.t16 source.n21 167.117
R91 source.t20 source.n33 167.117
R92 source.n9 source.n8 84.1169
R93 source.n11 source.n10 84.1169
R94 source.n29 source.n28 84.1169
R95 source.n31 source.n30 84.1169
R96 source.n71 source.n70 84.1168
R97 source.n69 source.n68 84.1168
R98 source.n51 source.n50 84.1168
R99 source.n49 source.n48 84.1168
R100 source.n74 source.t18 52.3082
R101 source.n62 source.t12 52.3082
R102 source.n54 source.t5 52.3082
R103 source.n42 source.t3 52.3082
R104 source.n2 source.t4 52.3082
R105 source.n14 source.t2 52.3082
R106 source.n22 source.t16 52.3082
R107 source.n34 source.t20 52.3082
R108 source.n79 source.n78 31.4096
R109 source.n67 source.n66 31.4096
R110 source.n59 source.n58 31.4096
R111 source.n47 source.n46 31.4096
R112 source.n7 source.n6 31.4096
R113 source.n19 source.n18 31.4096
R114 source.n27 source.n26 31.4096
R115 source.n39 source.n38 31.4096
R116 source.n47 source.n39 14.1689
R117 source.n70 source.t14 9.9005
R118 source.n70 source.t23 9.9005
R119 source.n68 source.t22 9.9005
R120 source.n68 source.t17 9.9005
R121 source.n50 source.t8 9.9005
R122 source.n50 source.t0 9.9005
R123 source.n48 source.t1 9.9005
R124 source.n48 source.t6 9.9005
R125 source.n8 source.t10 9.9005
R126 source.n8 source.t11 9.9005
R127 source.n10 source.t9 9.9005
R128 source.n10 source.t7 9.9005
R129 source.n28 source.t21 9.9005
R130 source.n28 source.t19 9.9005
R131 source.n30 source.t15 9.9005
R132 source.n30 source.t13 9.9005
R133 source.n75 source.n73 9.71174
R134 source.n63 source.n61 9.71174
R135 source.n55 source.n53 9.71174
R136 source.n43 source.n41 9.71174
R137 source.n3 source.n1 9.71174
R138 source.n15 source.n13 9.71174
R139 source.n23 source.n21 9.71174
R140 source.n35 source.n33 9.71174
R141 source.n78 source.n77 9.45567
R142 source.n66 source.n65 9.45567
R143 source.n58 source.n57 9.45567
R144 source.n46 source.n45 9.45567
R145 source.n6 source.n5 9.45567
R146 source.n18 source.n17 9.45567
R147 source.n26 source.n25 9.45567
R148 source.n38 source.n37 9.45567
R149 source.n77 source.n76 9.3005
R150 source.n65 source.n64 9.3005
R151 source.n57 source.n56 9.3005
R152 source.n45 source.n44 9.3005
R153 source.n5 source.n4 9.3005
R154 source.n17 source.n16 9.3005
R155 source.n25 source.n24 9.3005
R156 source.n37 source.n36 9.3005
R157 source.n80 source.n7 8.67749
R158 source.n78 source.n72 8.14595
R159 source.n66 source.n60 8.14595
R160 source.n58 source.n52 8.14595
R161 source.n46 source.n40 8.14595
R162 source.n6 source.n0 8.14595
R163 source.n18 source.n12 8.14595
R164 source.n26 source.n20 8.14595
R165 source.n38 source.n32 8.14595
R166 source.n76 source.n75 7.3702
R167 source.n64 source.n63 7.3702
R168 source.n56 source.n55 7.3702
R169 source.n44 source.n43 7.3702
R170 source.n4 source.n3 7.3702
R171 source.n16 source.n15 7.3702
R172 source.n24 source.n23 7.3702
R173 source.n36 source.n35 7.3702
R174 source.n76 source.n72 5.81868
R175 source.n64 source.n60 5.81868
R176 source.n56 source.n52 5.81868
R177 source.n44 source.n40 5.81868
R178 source.n4 source.n0 5.81868
R179 source.n16 source.n12 5.81868
R180 source.n24 source.n20 5.81868
R181 source.n36 source.n32 5.81868
R182 source.n80 source.n79 5.49188
R183 source.n77 source.n73 3.44771
R184 source.n65 source.n61 3.44771
R185 source.n57 source.n53 3.44771
R186 source.n45 source.n41 3.44771
R187 source.n5 source.n1 3.44771
R188 source.n17 source.n13 3.44771
R189 source.n25 source.n21 3.44771
R190 source.n37 source.n33 3.44771
R191 source.n27 source.n19 0.470328
R192 source.n67 source.n59 0.470328
R193 source.n39 source.n31 0.457397
R194 source.n31 source.n29 0.457397
R195 source.n29 source.n27 0.457397
R196 source.n19 source.n11 0.457397
R197 source.n11 source.n9 0.457397
R198 source.n9 source.n7 0.457397
R199 source.n49 source.n47 0.457397
R200 source.n51 source.n49 0.457397
R201 source.n59 source.n51 0.457397
R202 source.n69 source.n67 0.457397
R203 source.n71 source.n69 0.457397
R204 source.n79 source.n71 0.457397
R205 source source.n80 0.188
R206 plus.n2 plus.t5 445.12
R207 plus.n11 plus.t4 445.12
R208 plus.n15 plus.t10 445.12
R209 plus.n24 plus.t9 445.12
R210 plus.n3 plus.t2 397.651
R211 plus.n1 plus.t11 397.651
R212 plus.n8 plus.t8 397.651
R213 plus.n10 plus.t7 397.651
R214 plus.n16 plus.t1 397.651
R215 plus.n14 plus.t6 397.651
R216 plus.n21 plus.t0 397.651
R217 plus.n23 plus.t3 397.651
R218 plus.n5 plus.n2 161.489
R219 plus.n18 plus.n15 161.489
R220 plus.n5 plus.n4 161.3
R221 plus.n7 plus.n6 161.3
R222 plus.n9 plus.n0 161.3
R223 plus.n12 plus.n11 161.3
R224 plus.n18 plus.n17 161.3
R225 plus.n20 plus.n19 161.3
R226 plus.n22 plus.n13 161.3
R227 plus.n25 plus.n24 161.3
R228 plus.n4 plus.n3 43.0884
R229 plus.n10 plus.n9 43.0884
R230 plus.n23 plus.n22 43.0884
R231 plus.n17 plus.n16 43.0884
R232 plus.n7 plus.n1 38.7066
R233 plus.n8 plus.n7 38.7066
R234 plus.n21 plus.n20 38.7066
R235 plus.n20 plus.n14 38.7066
R236 plus.n4 plus.n1 34.3247
R237 plus.n9 plus.n8 34.3247
R238 plus.n22 plus.n21 34.3247
R239 plus.n17 plus.n14 34.3247
R240 plus.n3 plus.n2 29.9429
R241 plus.n11 plus.n10 29.9429
R242 plus.n24 plus.n23 29.9429
R243 plus.n16 plus.n15 29.9429
R244 plus plus.n25 24.6922
R245 plus plus.n12 8.31111
R246 plus.n6 plus.n5 0.189894
R247 plus.n6 plus.n0 0.189894
R248 plus.n12 plus.n0 0.189894
R249 plus.n25 plus.n13 0.189894
R250 plus.n19 plus.n13 0.189894
R251 plus.n19 plus.n18 0.189894
R252 drain_left.n6 drain_left.n4 101.252
R253 drain_left.n3 drain_left.n2 101.198
R254 drain_left.n3 drain_left.n0 101.198
R255 drain_left.n8 drain_left.n7 100.796
R256 drain_left.n6 drain_left.n5 100.796
R257 drain_left.n3 drain_left.n1 100.796
R258 drain_left drain_left.n3 22.0758
R259 drain_left.n1 drain_left.t11 9.9005
R260 drain_left.n1 drain_left.t5 9.9005
R261 drain_left.n2 drain_left.t10 9.9005
R262 drain_left.n2 drain_left.t1 9.9005
R263 drain_left.n0 drain_left.t2 9.9005
R264 drain_left.n0 drain_left.t8 9.9005
R265 drain_left.n7 drain_left.t4 9.9005
R266 drain_left.n7 drain_left.t7 9.9005
R267 drain_left.n5 drain_left.t0 9.9005
R268 drain_left.n5 drain_left.t3 9.9005
R269 drain_left.n4 drain_left.t6 9.9005
R270 drain_left.n4 drain_left.t9 9.9005
R271 drain_left drain_left.n8 6.11011
R272 drain_left.n8 drain_left.n6 0.457397
C0 drain_left minus 0.176308f
C1 drain_right plus 0.298665f
C2 source plus 1.02787f
C3 source drain_right 6.5528f
C4 drain_left plus 1.08189f
C5 minus plus 3.12867f
C6 drain_left drain_right 0.71208f
C7 drain_right minus 0.942983f
C8 drain_left source 6.55367f
C9 source minus 1.01391f
C10 drain_right a_n1458_n1288# 3.54992f
C11 drain_left a_n1458_n1288# 3.75544f
C12 source a_n1458_n1288# 2.933112f
C13 minus a_n1458_n1288# 4.837504f
C14 plus a_n1458_n1288# 5.531555f
C15 drain_left.t2 a_n1458_n1288# 0.046179f
C16 drain_left.t8 a_n1458_n1288# 0.046179f
C17 drain_left.n0 a_n1458_n1288# 0.291369f
C18 drain_left.t11 a_n1458_n1288# 0.046179f
C19 drain_left.t5 a_n1458_n1288# 0.046179f
C20 drain_left.n1 a_n1458_n1288# 0.290108f
C21 drain_left.t10 a_n1458_n1288# 0.046179f
C22 drain_left.t1 a_n1458_n1288# 0.046179f
C23 drain_left.n2 a_n1458_n1288# 0.291369f
C24 drain_left.n3 a_n1458_n1288# 1.61922f
C25 drain_left.t6 a_n1458_n1288# 0.046179f
C26 drain_left.t9 a_n1458_n1288# 0.046179f
C27 drain_left.n4 a_n1458_n1288# 0.291559f
C28 drain_left.t0 a_n1458_n1288# 0.046179f
C29 drain_left.t3 a_n1458_n1288# 0.046179f
C30 drain_left.n5 a_n1458_n1288# 0.290109f
C31 drain_left.n6 a_n1458_n1288# 0.62965f
C32 drain_left.t4 a_n1458_n1288# 0.046179f
C33 drain_left.t7 a_n1458_n1288# 0.046179f
C34 drain_left.n7 a_n1458_n1288# 0.290109f
C35 drain_left.n8 a_n1458_n1288# 0.548791f
C36 plus.n0 a_n1458_n1288# 0.034194f
C37 plus.t7 a_n1458_n1288# 0.040247f
C38 plus.t8 a_n1458_n1288# 0.040247f
C39 plus.t11 a_n1458_n1288# 0.040247f
C40 plus.n1 a_n1458_n1288# 0.031623f
C41 plus.t5 a_n1458_n1288# 0.043676f
C42 plus.n2 a_n1458_n1288# 0.040745f
C43 plus.t2 a_n1458_n1288# 0.040247f
C44 plus.n3 a_n1458_n1288# 0.031623f
C45 plus.n4 a_n1458_n1288# 0.011976f
C46 plus.n5 a_n1458_n1288# 0.075717f
C47 plus.n6 a_n1458_n1288# 0.034194f
C48 plus.n7 a_n1458_n1288# 0.011976f
C49 plus.n8 a_n1458_n1288# 0.031623f
C50 plus.n9 a_n1458_n1288# 0.011976f
C51 plus.n10 a_n1458_n1288# 0.031623f
C52 plus.t4 a_n1458_n1288# 0.043676f
C53 plus.n11 a_n1458_n1288# 0.040697f
C54 plus.n12 a_n1458_n1288# 0.240623f
C55 plus.n13 a_n1458_n1288# 0.034194f
C56 plus.t9 a_n1458_n1288# 0.043676f
C57 plus.t3 a_n1458_n1288# 0.040247f
C58 plus.t0 a_n1458_n1288# 0.040247f
C59 plus.t6 a_n1458_n1288# 0.040247f
C60 plus.n14 a_n1458_n1288# 0.031623f
C61 plus.t10 a_n1458_n1288# 0.043676f
C62 plus.n15 a_n1458_n1288# 0.040745f
C63 plus.t1 a_n1458_n1288# 0.040247f
C64 plus.n16 a_n1458_n1288# 0.031623f
C65 plus.n17 a_n1458_n1288# 0.011976f
C66 plus.n18 a_n1458_n1288# 0.075717f
C67 plus.n19 a_n1458_n1288# 0.034194f
C68 plus.n20 a_n1458_n1288# 0.011976f
C69 plus.n21 a_n1458_n1288# 0.031623f
C70 plus.n22 a_n1458_n1288# 0.011976f
C71 plus.n23 a_n1458_n1288# 0.031623f
C72 plus.n24 a_n1458_n1288# 0.040697f
C73 plus.n25 a_n1458_n1288# 0.708309f
C74 source.n0 a_n1458_n1288# 0.04287f
C75 source.n1 a_n1458_n1288# 0.094855f
C76 source.t4 a_n1458_n1288# 0.071183f
C77 source.n2 a_n1458_n1288# 0.074237f
C78 source.n3 a_n1458_n1288# 0.023931f
C79 source.n4 a_n1458_n1288# 0.015783f
C80 source.n5 a_n1458_n1288# 0.209082f
C81 source.n6 a_n1458_n1288# 0.046995f
C82 source.n7 a_n1458_n1288# 0.428954f
C83 source.t10 a_n1458_n1288# 0.046421f
C84 source.t11 a_n1458_n1288# 0.046421f
C85 source.n8 a_n1458_n1288# 0.248164f
C86 source.n9 a_n1458_n1288# 0.314834f
C87 source.t9 a_n1458_n1288# 0.046421f
C88 source.t7 a_n1458_n1288# 0.046421f
C89 source.n10 a_n1458_n1288# 0.248164f
C90 source.n11 a_n1458_n1288# 0.314834f
C91 source.n12 a_n1458_n1288# 0.04287f
C92 source.n13 a_n1458_n1288# 0.094854f
C93 source.t2 a_n1458_n1288# 0.071183f
C94 source.n14 a_n1458_n1288# 0.074237f
C95 source.n15 a_n1458_n1288# 0.023931f
C96 source.n16 a_n1458_n1288# 0.015783f
C97 source.n17 a_n1458_n1288# 0.209082f
C98 source.n18 a_n1458_n1288# 0.046995f
C99 source.n19 a_n1458_n1288# 0.111887f
C100 source.n20 a_n1458_n1288# 0.04287f
C101 source.n21 a_n1458_n1288# 0.094854f
C102 source.t16 a_n1458_n1288# 0.071183f
C103 source.n22 a_n1458_n1288# 0.074237f
C104 source.n23 a_n1458_n1288# 0.023931f
C105 source.n24 a_n1458_n1288# 0.015783f
C106 source.n25 a_n1458_n1288# 0.209082f
C107 source.n26 a_n1458_n1288# 0.046995f
C108 source.n27 a_n1458_n1288# 0.111887f
C109 source.t21 a_n1458_n1288# 0.046421f
C110 source.t19 a_n1458_n1288# 0.046421f
C111 source.n28 a_n1458_n1288# 0.248164f
C112 source.n29 a_n1458_n1288# 0.314834f
C113 source.t15 a_n1458_n1288# 0.046421f
C114 source.t13 a_n1458_n1288# 0.046421f
C115 source.n30 a_n1458_n1288# 0.248164f
C116 source.n31 a_n1458_n1288# 0.314834f
C117 source.n32 a_n1458_n1288# 0.04287f
C118 source.n33 a_n1458_n1288# 0.094854f
C119 source.t20 a_n1458_n1288# 0.071183f
C120 source.n34 a_n1458_n1288# 0.074237f
C121 source.n35 a_n1458_n1288# 0.023931f
C122 source.n36 a_n1458_n1288# 0.015783f
C123 source.n37 a_n1458_n1288# 0.209082f
C124 source.n38 a_n1458_n1288# 0.046995f
C125 source.n39 a_n1458_n1288# 0.700979f
C126 source.n40 a_n1458_n1288# 0.04287f
C127 source.n41 a_n1458_n1288# 0.094854f
C128 source.t3 a_n1458_n1288# 0.071184f
C129 source.n42 a_n1458_n1288# 0.074237f
C130 source.n43 a_n1458_n1288# 0.023931f
C131 source.n44 a_n1458_n1288# 0.015783f
C132 source.n45 a_n1458_n1288# 0.209082f
C133 source.n46 a_n1458_n1288# 0.046995f
C134 source.n47 a_n1458_n1288# 0.700979f
C135 source.t1 a_n1458_n1288# 0.046421f
C136 source.t6 a_n1458_n1288# 0.046421f
C137 source.n48 a_n1458_n1288# 0.248162f
C138 source.n49 a_n1458_n1288# 0.314836f
C139 source.t8 a_n1458_n1288# 0.046421f
C140 source.t0 a_n1458_n1288# 0.046421f
C141 source.n50 a_n1458_n1288# 0.248162f
C142 source.n51 a_n1458_n1288# 0.314836f
C143 source.n52 a_n1458_n1288# 0.04287f
C144 source.n53 a_n1458_n1288# 0.094854f
C145 source.t5 a_n1458_n1288# 0.071184f
C146 source.n54 a_n1458_n1288# 0.074237f
C147 source.n55 a_n1458_n1288# 0.023931f
C148 source.n56 a_n1458_n1288# 0.015783f
C149 source.n57 a_n1458_n1288# 0.209082f
C150 source.n58 a_n1458_n1288# 0.046995f
C151 source.n59 a_n1458_n1288# 0.111887f
C152 source.n60 a_n1458_n1288# 0.04287f
C153 source.n61 a_n1458_n1288# 0.094854f
C154 source.t12 a_n1458_n1288# 0.071184f
C155 source.n62 a_n1458_n1288# 0.074237f
C156 source.n63 a_n1458_n1288# 0.023931f
C157 source.n64 a_n1458_n1288# 0.015783f
C158 source.n65 a_n1458_n1288# 0.209082f
C159 source.n66 a_n1458_n1288# 0.046995f
C160 source.n67 a_n1458_n1288# 0.111887f
C161 source.t22 a_n1458_n1288# 0.046421f
C162 source.t17 a_n1458_n1288# 0.046421f
C163 source.n68 a_n1458_n1288# 0.248162f
C164 source.n69 a_n1458_n1288# 0.314836f
C165 source.t14 a_n1458_n1288# 0.046421f
C166 source.t23 a_n1458_n1288# 0.046421f
C167 source.n70 a_n1458_n1288# 0.248162f
C168 source.n71 a_n1458_n1288# 0.314836f
C169 source.n72 a_n1458_n1288# 0.04287f
C170 source.n73 a_n1458_n1288# 0.094854f
C171 source.t18 a_n1458_n1288# 0.071184f
C172 source.n74 a_n1458_n1288# 0.074237f
C173 source.n75 a_n1458_n1288# 0.023931f
C174 source.n76 a_n1458_n1288# 0.015783f
C175 source.n77 a_n1458_n1288# 0.209082f
C176 source.n78 a_n1458_n1288# 0.046995f
C177 source.n79 a_n1458_n1288# 0.271149f
C178 source.n80 a_n1458_n1288# 0.722747f
C179 drain_right.t8 a_n1458_n1288# 0.046992f
C180 drain_right.t2 a_n1458_n1288# 0.046992f
C181 drain_right.n0 a_n1458_n1288# 0.296504f
C182 drain_right.t5 a_n1458_n1288# 0.046992f
C183 drain_right.t6 a_n1458_n1288# 0.046992f
C184 drain_right.n1 a_n1458_n1288# 0.29522f
C185 drain_right.t7 a_n1458_n1288# 0.046992f
C186 drain_right.t9 a_n1458_n1288# 0.046992f
C187 drain_right.n2 a_n1458_n1288# 0.296504f
C188 drain_right.n3 a_n1458_n1288# 1.58928f
C189 drain_right.t3 a_n1458_n1288# 0.046992f
C190 drain_right.t0 a_n1458_n1288# 0.046992f
C191 drain_right.n4 a_n1458_n1288# 0.296698f
C192 drain_right.t1 a_n1458_n1288# 0.046992f
C193 drain_right.t4 a_n1458_n1288# 0.046992f
C194 drain_right.n5 a_n1458_n1288# 0.295222f
C195 drain_right.n6 a_n1458_n1288# 0.640746f
C196 drain_right.t10 a_n1458_n1288# 0.046992f
C197 drain_right.t11 a_n1458_n1288# 0.046992f
C198 drain_right.n7 a_n1458_n1288# 0.295222f
C199 drain_right.n8 a_n1458_n1288# 0.558462f
C200 minus.n0 a_n1458_n1288# 0.033447f
C201 minus.t3 a_n1458_n1288# 0.042723f
C202 minus.t8 a_n1458_n1288# 0.039369f
C203 minus.t10 a_n1458_n1288# 0.039369f
C204 minus.t2 a_n1458_n1288# 0.039369f
C205 minus.n1 a_n1458_n1288# 0.030933f
C206 minus.t7 a_n1458_n1288# 0.042723f
C207 minus.n2 a_n1458_n1288# 0.039856f
C208 minus.t4 a_n1458_n1288# 0.039369f
C209 minus.n3 a_n1458_n1288# 0.030933f
C210 minus.n4 a_n1458_n1288# 0.011714f
C211 minus.n5 a_n1458_n1288# 0.074065f
C212 minus.n6 a_n1458_n1288# 0.033447f
C213 minus.n7 a_n1458_n1288# 0.011714f
C214 minus.n8 a_n1458_n1288# 0.030933f
C215 minus.n9 a_n1458_n1288# 0.011714f
C216 minus.n10 a_n1458_n1288# 0.030933f
C217 minus.n11 a_n1458_n1288# 0.039809f
C218 minus.n12 a_n1458_n1288# 0.722741f
C219 minus.n13 a_n1458_n1288# 0.033447f
C220 minus.t0 a_n1458_n1288# 0.039369f
C221 minus.t9 a_n1458_n1288# 0.039369f
C222 minus.t6 a_n1458_n1288# 0.039369f
C223 minus.n14 a_n1458_n1288# 0.030933f
C224 minus.t11 a_n1458_n1288# 0.042723f
C225 minus.n15 a_n1458_n1288# 0.039856f
C226 minus.t1 a_n1458_n1288# 0.039369f
C227 minus.n16 a_n1458_n1288# 0.030933f
C228 minus.n17 a_n1458_n1288# 0.011714f
C229 minus.n18 a_n1458_n1288# 0.074065f
C230 minus.n19 a_n1458_n1288# 0.033447f
C231 minus.n20 a_n1458_n1288# 0.011714f
C232 minus.n21 a_n1458_n1288# 0.030933f
C233 minus.n22 a_n1458_n1288# 0.011714f
C234 minus.n23 a_n1458_n1288# 0.030933f
C235 minus.t5 a_n1458_n1288# 0.042723f
C236 minus.n24 a_n1458_n1288# 0.039809f
C237 minus.n25 a_n1458_n1288# 0.21512f
C238 minus.n26 a_n1458_n1288# 0.895338f
.ends

