* NGSPICE file created from diffpair498.ext - technology: sky130A

.subckt diffpair498 minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t28 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X1 drain_left.t18 plus.t1 source.t37 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X2 drain_left.t17 plus.t2 source.t36 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X3 drain_right.t19 minus.t0 source.t12 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X4 drain_right.t18 minus.t1 source.t15 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X5 source.t25 plus.t3 drain_left.t16 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X6 source.t24 plus.t4 drain_left.t15 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X7 drain_left.t14 plus.t5 source.t31 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X8 source.t9 minus.t2 drain_right.t17 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X9 source.t11 minus.t3 drain_right.t16 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X10 source.t7 minus.t4 drain_right.t15 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X11 source.t1 minus.t5 drain_right.t14 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X12 drain_left.t13 plus.t6 source.t20 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X13 source.t3 minus.t6 drain_right.t13 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X14 drain_left.t12 plus.t7 source.t22 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X15 source.t33 plus.t8 drain_left.t11 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X16 drain_right.t12 minus.t7 source.t8 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X17 drain_right.t11 minus.t8 source.t2 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X18 drain_right.t10 minus.t9 source.t6 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X19 a_n1882_n3888# a_n1882_n3888# a_n1882_n3888# a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.2
X20 drain_right.t9 minus.t10 source.t10 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X21 drain_right.t8 minus.t11 source.t13 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X22 drain_right.t7 minus.t12 source.t16 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X23 source.t17 minus.t13 drain_right.t6 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X24 drain_right.t5 minus.t14 source.t38 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X25 drain_right.t4 minus.t15 source.t39 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X26 source.t5 minus.t16 drain_right.t3 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X27 source.t32 plus.t9 drain_left.t10 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X28 source.t0 minus.t17 drain_right.t2 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X29 source.t34 plus.t10 drain_left.t9 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X30 a_n1882_n3888# a_n1882_n3888# a_n1882_n3888# a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X31 drain_left.t8 plus.t11 source.t18 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X32 source.t29 plus.t12 drain_left.t7 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X33 drain_left.t6 plus.t13 source.t30 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X34 a_n1882_n3888# a_n1882_n3888# a_n1882_n3888# a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X35 source.t4 minus.t18 drain_right.t1 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X36 source.t14 minus.t19 drain_right.t0 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X37 source.t23 plus.t14 drain_left.t5 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X38 source.t21 plus.t15 drain_left.t4 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X39 source.t19 plus.t16 drain_left.t3 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X40 drain_left.t2 plus.t17 source.t35 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X41 source.t27 plus.t18 drain_left.t1 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X42 a_n1882_n3888# a_n1882_n3888# a_n1882_n3888# a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X43 drain_left.t0 plus.t19 source.t26 a_n1882_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
R0 plus.n5 plus.t8 2020.38
R1 plus.n23 plus.t6 2020.38
R2 plus.n30 plus.t2 2020.38
R3 plus.n48 plus.t9 2020.38
R4 plus.n6 plus.t5 1964.15
R5 plus.n8 plus.t18 1964.15
R6 plus.n3 plus.t13 1964.15
R7 plus.n13 plus.t12 1964.15
R8 plus.n15 plus.t7 1964.15
R9 plus.n1 plus.t4 1964.15
R10 plus.n20 plus.t17 1964.15
R11 plus.n22 plus.t10 1964.15
R12 plus.n31 plus.t3 1964.15
R13 plus.n33 plus.t1 1964.15
R14 plus.n28 plus.t15 1964.15
R15 plus.n38 plus.t0 1964.15
R16 plus.n40 plus.t16 1964.15
R17 plus.n26 plus.t19 1964.15
R18 plus.n45 plus.t14 1964.15
R19 plus.n47 plus.t11 1964.15
R20 plus.n5 plus.n4 161.489
R21 plus.n30 plus.n29 161.489
R22 plus.n7 plus.n4 161.3
R23 plus.n10 plus.n9 161.3
R24 plus.n12 plus.n11 161.3
R25 plus.n14 plus.n2 161.3
R26 plus.n17 plus.n16 161.3
R27 plus.n19 plus.n18 161.3
R28 plus.n21 plus.n0 161.3
R29 plus.n24 plus.n23 161.3
R30 plus.n32 plus.n29 161.3
R31 plus.n35 plus.n34 161.3
R32 plus.n37 plus.n36 161.3
R33 plus.n39 plus.n27 161.3
R34 plus.n42 plus.n41 161.3
R35 plus.n44 plus.n43 161.3
R36 plus.n46 plus.n25 161.3
R37 plus.n49 plus.n48 161.3
R38 plus.n7 plus.n6 51.852
R39 plus.n22 plus.n21 51.852
R40 plus.n47 plus.n46 51.852
R41 plus.n32 plus.n31 51.852
R42 plus.n9 plus.n8 47.4702
R43 plus.n20 plus.n19 47.4702
R44 plus.n45 plus.n44 47.4702
R45 plus.n34 plus.n33 47.4702
R46 plus.n12 plus.n3 43.0884
R47 plus.n16 plus.n1 43.0884
R48 plus.n41 plus.n26 43.0884
R49 plus.n37 plus.n28 43.0884
R50 plus.n14 plus.n13 38.7066
R51 plus.n15 plus.n14 38.7066
R52 plus.n40 plus.n39 38.7066
R53 plus.n39 plus.n38 38.7066
R54 plus.n13 plus.n12 34.3247
R55 plus.n16 plus.n15 34.3247
R56 plus.n41 plus.n40 34.3247
R57 plus.n38 plus.n37 34.3247
R58 plus plus.n49 31.2452
R59 plus.n9 plus.n3 29.9429
R60 plus.n19 plus.n1 29.9429
R61 plus.n44 plus.n26 29.9429
R62 plus.n34 plus.n28 29.9429
R63 plus.n8 plus.n7 25.5611
R64 plus.n21 plus.n20 25.5611
R65 plus.n46 plus.n45 25.5611
R66 plus.n33 plus.n32 25.5611
R67 plus.n6 plus.n5 21.1793
R68 plus.n23 plus.n22 21.1793
R69 plus.n48 plus.n47 21.1793
R70 plus.n31 plus.n30 21.1793
R71 plus plus.n24 13.2581
R72 plus.n10 plus.n4 0.189894
R73 plus.n11 plus.n10 0.189894
R74 plus.n11 plus.n2 0.189894
R75 plus.n17 plus.n2 0.189894
R76 plus.n18 plus.n17 0.189894
R77 plus.n18 plus.n0 0.189894
R78 plus.n24 plus.n0 0.189894
R79 plus.n49 plus.n25 0.189894
R80 plus.n43 plus.n25 0.189894
R81 plus.n43 plus.n42 0.189894
R82 plus.n42 plus.n27 0.189894
R83 plus.n36 plus.n27 0.189894
R84 plus.n36 plus.n35 0.189894
R85 plus.n35 plus.n29 0.189894
R86 source.n9 source.t33 45.521
R87 source.n10 source.t38 45.521
R88 source.n19 source.t3 45.521
R89 source.n39 source.t8 45.5208
R90 source.n30 source.t1 45.5208
R91 source.n29 source.t36 45.5208
R92 source.n20 source.t32 45.5208
R93 source.n0 source.t20 45.5208
R94 source.n2 source.n1 44.201
R95 source.n4 source.n3 44.201
R96 source.n6 source.n5 44.201
R97 source.n8 source.n7 44.201
R98 source.n12 source.n11 44.201
R99 source.n14 source.n13 44.201
R100 source.n16 source.n15 44.201
R101 source.n18 source.n17 44.201
R102 source.n38 source.n37 44.2008
R103 source.n36 source.n35 44.2008
R104 source.n34 source.n33 44.2008
R105 source.n32 source.n31 44.2008
R106 source.n28 source.n27 44.2008
R107 source.n26 source.n25 44.2008
R108 source.n24 source.n23 44.2008
R109 source.n22 source.n21 44.2008
R110 source.n20 source.n19 24.0173
R111 source.n40 source.n0 18.526
R112 source.n40 source.n39 5.49188
R113 source.n37 source.t10 1.3205
R114 source.n37 source.t17 1.3205
R115 source.n35 source.t13 1.3205
R116 source.n35 source.t5 1.3205
R117 source.n33 source.t2 1.3205
R118 source.n33 source.t0 1.3205
R119 source.n31 source.t6 1.3205
R120 source.n31 source.t11 1.3205
R121 source.n27 source.t37 1.3205
R122 source.n27 source.t25 1.3205
R123 source.n25 source.t28 1.3205
R124 source.n25 source.t21 1.3205
R125 source.n23 source.t26 1.3205
R126 source.n23 source.t19 1.3205
R127 source.n21 source.t18 1.3205
R128 source.n21 source.t23 1.3205
R129 source.n1 source.t35 1.3205
R130 source.n1 source.t34 1.3205
R131 source.n3 source.t22 1.3205
R132 source.n3 source.t24 1.3205
R133 source.n5 source.t30 1.3205
R134 source.n5 source.t29 1.3205
R135 source.n7 source.t31 1.3205
R136 source.n7 source.t27 1.3205
R137 source.n11 source.t12 1.3205
R138 source.n11 source.t7 1.3205
R139 source.n13 source.t39 1.3205
R140 source.n13 source.t4 1.3205
R141 source.n15 source.t15 1.3205
R142 source.n15 source.t9 1.3205
R143 source.n17 source.t16 1.3205
R144 source.n17 source.t14 1.3205
R145 source.n10 source.n9 0.470328
R146 source.n30 source.n29 0.470328
R147 source.n19 source.n18 0.457397
R148 source.n18 source.n16 0.457397
R149 source.n16 source.n14 0.457397
R150 source.n14 source.n12 0.457397
R151 source.n12 source.n10 0.457397
R152 source.n9 source.n8 0.457397
R153 source.n8 source.n6 0.457397
R154 source.n6 source.n4 0.457397
R155 source.n4 source.n2 0.457397
R156 source.n2 source.n0 0.457397
R157 source.n22 source.n20 0.457397
R158 source.n24 source.n22 0.457397
R159 source.n26 source.n24 0.457397
R160 source.n28 source.n26 0.457397
R161 source.n29 source.n28 0.457397
R162 source.n32 source.n30 0.457397
R163 source.n34 source.n32 0.457397
R164 source.n36 source.n34 0.457397
R165 source.n38 source.n36 0.457397
R166 source.n39 source.n38 0.457397
R167 source source.n40 0.188
R168 drain_left.n10 drain_left.n8 61.3367
R169 drain_left.n6 drain_left.n4 61.3365
R170 drain_left.n2 drain_left.n0 61.3365
R171 drain_left.n14 drain_left.n13 60.8798
R172 drain_left.n12 drain_left.n11 60.8798
R173 drain_left.n10 drain_left.n9 60.8798
R174 drain_left.n16 drain_left.n15 60.8796
R175 drain_left.n7 drain_left.n3 60.8796
R176 drain_left.n6 drain_left.n5 60.8796
R177 drain_left.n2 drain_left.n1 60.8796
R178 drain_left drain_left.n7 33.295
R179 drain_left drain_left.n16 6.11011
R180 drain_left.n3 drain_left.t3 1.3205
R181 drain_left.n3 drain_left.t19 1.3205
R182 drain_left.n4 drain_left.t16 1.3205
R183 drain_left.n4 drain_left.t17 1.3205
R184 drain_left.n5 drain_left.t4 1.3205
R185 drain_left.n5 drain_left.t18 1.3205
R186 drain_left.n1 drain_left.t5 1.3205
R187 drain_left.n1 drain_left.t0 1.3205
R188 drain_left.n0 drain_left.t10 1.3205
R189 drain_left.n0 drain_left.t8 1.3205
R190 drain_left.n15 drain_left.t9 1.3205
R191 drain_left.n15 drain_left.t13 1.3205
R192 drain_left.n13 drain_left.t15 1.3205
R193 drain_left.n13 drain_left.t2 1.3205
R194 drain_left.n11 drain_left.t7 1.3205
R195 drain_left.n11 drain_left.t12 1.3205
R196 drain_left.n9 drain_left.t1 1.3205
R197 drain_left.n9 drain_left.t6 1.3205
R198 drain_left.n8 drain_left.t11 1.3205
R199 drain_left.n8 drain_left.t14 1.3205
R200 drain_left.n12 drain_left.n10 0.457397
R201 drain_left.n14 drain_left.n12 0.457397
R202 drain_left.n16 drain_left.n14 0.457397
R203 drain_left.n7 drain_left.n6 0.402051
R204 drain_left.n7 drain_left.n2 0.402051
R205 minus.n23 minus.t6 2020.38
R206 minus.n5 minus.t14 2020.38
R207 minus.n48 minus.t7 2020.38
R208 minus.n30 minus.t5 2020.38
R209 minus.n22 minus.t12 1964.15
R210 minus.n20 minus.t19 1964.15
R211 minus.n1 minus.t1 1964.15
R212 minus.n15 minus.t2 1964.15
R213 minus.n13 minus.t15 1964.15
R214 minus.n3 minus.t18 1964.15
R215 minus.n8 minus.t0 1964.15
R216 minus.n6 minus.t4 1964.15
R217 minus.n47 minus.t13 1964.15
R218 minus.n45 minus.t10 1964.15
R219 minus.n26 minus.t16 1964.15
R220 minus.n40 minus.t11 1964.15
R221 minus.n38 minus.t17 1964.15
R222 minus.n28 minus.t8 1964.15
R223 minus.n33 minus.t3 1964.15
R224 minus.n31 minus.t9 1964.15
R225 minus.n5 minus.n4 161.489
R226 minus.n30 minus.n29 161.489
R227 minus.n24 minus.n23 161.3
R228 minus.n21 minus.n0 161.3
R229 minus.n19 minus.n18 161.3
R230 minus.n17 minus.n16 161.3
R231 minus.n14 minus.n2 161.3
R232 minus.n12 minus.n11 161.3
R233 minus.n10 minus.n9 161.3
R234 minus.n7 minus.n4 161.3
R235 minus.n49 minus.n48 161.3
R236 minus.n46 minus.n25 161.3
R237 minus.n44 minus.n43 161.3
R238 minus.n42 minus.n41 161.3
R239 minus.n39 minus.n27 161.3
R240 minus.n37 minus.n36 161.3
R241 minus.n35 minus.n34 161.3
R242 minus.n32 minus.n29 161.3
R243 minus.n22 minus.n21 51.852
R244 minus.n7 minus.n6 51.852
R245 minus.n32 minus.n31 51.852
R246 minus.n47 minus.n46 51.852
R247 minus.n20 minus.n19 47.4702
R248 minus.n9 minus.n8 47.4702
R249 minus.n34 minus.n33 47.4702
R250 minus.n45 minus.n44 47.4702
R251 minus.n16 minus.n1 43.0884
R252 minus.n12 minus.n3 43.0884
R253 minus.n37 minus.n28 43.0884
R254 minus.n41 minus.n26 43.0884
R255 minus.n15 minus.n14 38.7066
R256 minus.n14 minus.n13 38.7066
R257 minus.n39 minus.n38 38.7066
R258 minus.n40 minus.n39 38.7066
R259 minus.n50 minus.n24 38.5005
R260 minus.n16 minus.n15 34.3247
R261 minus.n13 minus.n12 34.3247
R262 minus.n38 minus.n37 34.3247
R263 minus.n41 minus.n40 34.3247
R264 minus.n19 minus.n1 29.9429
R265 minus.n9 minus.n3 29.9429
R266 minus.n34 minus.n28 29.9429
R267 minus.n44 minus.n26 29.9429
R268 minus.n21 minus.n20 25.5611
R269 minus.n8 minus.n7 25.5611
R270 minus.n33 minus.n32 25.5611
R271 minus.n46 minus.n45 25.5611
R272 minus.n23 minus.n22 21.1793
R273 minus.n6 minus.n5 21.1793
R274 minus.n31 minus.n30 21.1793
R275 minus.n48 minus.n47 21.1793
R276 minus.n50 minus.n49 6.47777
R277 minus.n24 minus.n0 0.189894
R278 minus.n18 minus.n0 0.189894
R279 minus.n18 minus.n17 0.189894
R280 minus.n17 minus.n2 0.189894
R281 minus.n11 minus.n2 0.189894
R282 minus.n11 minus.n10 0.189894
R283 minus.n10 minus.n4 0.189894
R284 minus.n35 minus.n29 0.189894
R285 minus.n36 minus.n35 0.189894
R286 minus.n36 minus.n27 0.189894
R287 minus.n42 minus.n27 0.189894
R288 minus.n43 minus.n42 0.189894
R289 minus.n43 minus.n25 0.189894
R290 minus.n49 minus.n25 0.189894
R291 minus minus.n50 0.188
R292 drain_right.n10 drain_right.n8 61.3365
R293 drain_right.n6 drain_right.n4 61.3365
R294 drain_right.n2 drain_right.n0 61.3365
R295 drain_right.n10 drain_right.n9 60.8798
R296 drain_right.n12 drain_right.n11 60.8798
R297 drain_right.n14 drain_right.n13 60.8798
R298 drain_right.n16 drain_right.n15 60.8798
R299 drain_right.n7 drain_right.n3 60.8796
R300 drain_right.n6 drain_right.n5 60.8796
R301 drain_right.n2 drain_right.n1 60.8796
R302 drain_right drain_right.n7 32.7417
R303 drain_right drain_right.n16 6.11011
R304 drain_right.n3 drain_right.t2 1.3205
R305 drain_right.n3 drain_right.t8 1.3205
R306 drain_right.n4 drain_right.t6 1.3205
R307 drain_right.n4 drain_right.t12 1.3205
R308 drain_right.n5 drain_right.t3 1.3205
R309 drain_right.n5 drain_right.t9 1.3205
R310 drain_right.n1 drain_right.t16 1.3205
R311 drain_right.n1 drain_right.t11 1.3205
R312 drain_right.n0 drain_right.t14 1.3205
R313 drain_right.n0 drain_right.t10 1.3205
R314 drain_right.n8 drain_right.t15 1.3205
R315 drain_right.n8 drain_right.t5 1.3205
R316 drain_right.n9 drain_right.t1 1.3205
R317 drain_right.n9 drain_right.t19 1.3205
R318 drain_right.n11 drain_right.t17 1.3205
R319 drain_right.n11 drain_right.t4 1.3205
R320 drain_right.n13 drain_right.t0 1.3205
R321 drain_right.n13 drain_right.t18 1.3205
R322 drain_right.n15 drain_right.t13 1.3205
R323 drain_right.n15 drain_right.t7 1.3205
R324 drain_right.n16 drain_right.n14 0.457397
R325 drain_right.n14 drain_right.n12 0.457397
R326 drain_right.n12 drain_right.n10 0.457397
R327 drain_right.n7 drain_right.n6 0.402051
R328 drain_right.n7 drain_right.n2 0.402051
C0 plus drain_right 0.337271f
C1 plus minus 6.05723f
C2 drain_left plus 6.69466f
C3 source drain_right 55.7054f
C4 source minus 6.01706f
C5 source drain_left 55.7055f
C6 minus drain_right 6.5116f
C7 drain_left drain_right 0.982035f
C8 drain_left minus 0.171252f
C9 source plus 6.0311f
C10 drain_right a_n1882_n3888# 7.83197f
C11 drain_left a_n1882_n3888# 8.133161f
C12 source a_n1882_n3888# 10.200675f
C13 minus a_n1882_n3888# 7.513767f
C14 plus a_n1882_n3888# 9.81307f
C15 drain_right.t14 a_n1882_n3888# 0.463499f
C16 drain_right.t10 a_n1882_n3888# 0.463499f
C17 drain_right.n0 a_n1882_n3888# 4.19285f
C18 drain_right.t16 a_n1882_n3888# 0.463499f
C19 drain_right.t11 a_n1882_n3888# 0.463499f
C20 drain_right.n1 a_n1882_n3888# 4.18949f
C21 drain_right.n2 a_n1882_n3888# 0.878488f
C22 drain_right.t2 a_n1882_n3888# 0.463499f
C23 drain_right.t8 a_n1882_n3888# 0.463499f
C24 drain_right.n3 a_n1882_n3888# 4.18949f
C25 drain_right.t6 a_n1882_n3888# 0.463499f
C26 drain_right.t12 a_n1882_n3888# 0.463499f
C27 drain_right.n4 a_n1882_n3888# 4.19285f
C28 drain_right.t3 a_n1882_n3888# 0.463499f
C29 drain_right.t9 a_n1882_n3888# 0.463499f
C30 drain_right.n5 a_n1882_n3888# 4.18949f
C31 drain_right.n6 a_n1882_n3888# 0.878488f
C32 drain_right.n7 a_n1882_n3888# 2.50063f
C33 drain_right.t15 a_n1882_n3888# 0.463499f
C34 drain_right.t5 a_n1882_n3888# 0.463499f
C35 drain_right.n8 a_n1882_n3888# 4.19284f
C36 drain_right.t1 a_n1882_n3888# 0.463499f
C37 drain_right.t19 a_n1882_n3888# 0.463499f
C38 drain_right.n9 a_n1882_n3888# 4.18949f
C39 drain_right.n10 a_n1882_n3888# 0.883212f
C40 drain_right.t17 a_n1882_n3888# 0.463499f
C41 drain_right.t4 a_n1882_n3888# 0.463499f
C42 drain_right.n11 a_n1882_n3888# 4.18949f
C43 drain_right.n12 a_n1882_n3888# 0.435404f
C44 drain_right.t0 a_n1882_n3888# 0.463499f
C45 drain_right.t18 a_n1882_n3888# 0.463499f
C46 drain_right.n13 a_n1882_n3888# 4.18949f
C47 drain_right.n14 a_n1882_n3888# 0.435404f
C48 drain_right.t13 a_n1882_n3888# 0.463499f
C49 drain_right.t7 a_n1882_n3888# 0.463499f
C50 drain_right.n15 a_n1882_n3888# 4.18949f
C51 drain_right.n16 a_n1882_n3888# 0.75542f
C52 minus.n0 a_n1882_n3888# 0.052791f
C53 minus.t6 a_n1882_n3888# 0.451794f
C54 minus.t12 a_n1882_n3888# 0.44679f
C55 minus.t19 a_n1882_n3888# 0.44679f
C56 minus.t1 a_n1882_n3888# 0.44679f
C57 minus.n1 a_n1882_n3888# 0.177039f
C58 minus.n2 a_n1882_n3888# 0.052791f
C59 minus.t2 a_n1882_n3888# 0.44679f
C60 minus.t15 a_n1882_n3888# 0.44679f
C61 minus.t18 a_n1882_n3888# 0.44679f
C62 minus.n3 a_n1882_n3888# 0.177039f
C63 minus.n4 a_n1882_n3888# 0.120798f
C64 minus.t0 a_n1882_n3888# 0.44679f
C65 minus.t4 a_n1882_n3888# 0.44679f
C66 minus.t14 a_n1882_n3888# 0.451794f
C67 minus.n5 a_n1882_n3888# 0.19337f
C68 minus.n6 a_n1882_n3888# 0.177039f
C69 minus.n7 a_n1882_n3888# 0.018489f
C70 minus.n8 a_n1882_n3888# 0.177039f
C71 minus.n9 a_n1882_n3888# 0.018489f
C72 minus.n10 a_n1882_n3888# 0.052791f
C73 minus.n11 a_n1882_n3888# 0.052791f
C74 minus.n12 a_n1882_n3888# 0.018489f
C75 minus.n13 a_n1882_n3888# 0.177039f
C76 minus.n14 a_n1882_n3888# 0.018489f
C77 minus.n15 a_n1882_n3888# 0.177039f
C78 minus.n16 a_n1882_n3888# 0.018489f
C79 minus.n17 a_n1882_n3888# 0.052791f
C80 minus.n18 a_n1882_n3888# 0.052791f
C81 minus.n19 a_n1882_n3888# 0.018489f
C82 minus.n20 a_n1882_n3888# 0.177039f
C83 minus.n21 a_n1882_n3888# 0.018489f
C84 minus.n22 a_n1882_n3888# 0.177039f
C85 minus.n23 a_n1882_n3888# 0.19329f
C86 minus.n24 a_n1882_n3888# 2.05147f
C87 minus.n25 a_n1882_n3888# 0.052791f
C88 minus.t13 a_n1882_n3888# 0.44679f
C89 minus.t10 a_n1882_n3888# 0.44679f
C90 minus.t16 a_n1882_n3888# 0.44679f
C91 minus.n26 a_n1882_n3888# 0.177039f
C92 minus.n27 a_n1882_n3888# 0.052791f
C93 minus.t11 a_n1882_n3888# 0.44679f
C94 minus.t17 a_n1882_n3888# 0.44679f
C95 minus.t8 a_n1882_n3888# 0.44679f
C96 minus.n28 a_n1882_n3888# 0.177039f
C97 minus.n29 a_n1882_n3888# 0.120798f
C98 minus.t3 a_n1882_n3888# 0.44679f
C99 minus.t9 a_n1882_n3888# 0.44679f
C100 minus.t5 a_n1882_n3888# 0.451794f
C101 minus.n30 a_n1882_n3888# 0.19337f
C102 minus.n31 a_n1882_n3888# 0.177039f
C103 minus.n32 a_n1882_n3888# 0.018489f
C104 minus.n33 a_n1882_n3888# 0.177039f
C105 minus.n34 a_n1882_n3888# 0.018489f
C106 minus.n35 a_n1882_n3888# 0.052791f
C107 minus.n36 a_n1882_n3888# 0.052791f
C108 minus.n37 a_n1882_n3888# 0.018489f
C109 minus.n38 a_n1882_n3888# 0.177039f
C110 minus.n39 a_n1882_n3888# 0.018489f
C111 minus.n40 a_n1882_n3888# 0.177039f
C112 minus.n41 a_n1882_n3888# 0.018489f
C113 minus.n42 a_n1882_n3888# 0.052791f
C114 minus.n43 a_n1882_n3888# 0.052791f
C115 minus.n44 a_n1882_n3888# 0.018489f
C116 minus.n45 a_n1882_n3888# 0.177039f
C117 minus.n46 a_n1882_n3888# 0.018489f
C118 minus.n47 a_n1882_n3888# 0.177039f
C119 minus.t7 a_n1882_n3888# 0.451794f
C120 minus.n48 a_n1882_n3888# 0.19329f
C121 minus.n49 a_n1882_n3888# 0.342363f
C122 minus.n50 a_n1882_n3888# 2.47582f
C123 drain_left.t10 a_n1882_n3888# 0.463848f
C124 drain_left.t8 a_n1882_n3888# 0.463848f
C125 drain_left.n0 a_n1882_n3888# 4.19601f
C126 drain_left.t5 a_n1882_n3888# 0.463848f
C127 drain_left.t0 a_n1882_n3888# 0.463848f
C128 drain_left.n1 a_n1882_n3888# 4.19265f
C129 drain_left.n2 a_n1882_n3888# 0.879151f
C130 drain_left.t3 a_n1882_n3888# 0.463848f
C131 drain_left.t19 a_n1882_n3888# 0.463848f
C132 drain_left.n3 a_n1882_n3888# 4.19265f
C133 drain_left.t16 a_n1882_n3888# 0.463848f
C134 drain_left.t17 a_n1882_n3888# 0.463848f
C135 drain_left.n4 a_n1882_n3888# 4.19601f
C136 drain_left.t4 a_n1882_n3888# 0.463848f
C137 drain_left.t18 a_n1882_n3888# 0.463848f
C138 drain_left.n5 a_n1882_n3888# 4.19265f
C139 drain_left.n6 a_n1882_n3888# 0.879151f
C140 drain_left.n7 a_n1882_n3888# 2.58389f
C141 drain_left.t11 a_n1882_n3888# 0.463848f
C142 drain_left.t14 a_n1882_n3888# 0.463848f
C143 drain_left.n8 a_n1882_n3888# 4.19601f
C144 drain_left.t1 a_n1882_n3888# 0.463848f
C145 drain_left.t6 a_n1882_n3888# 0.463848f
C146 drain_left.n9 a_n1882_n3888# 4.19265f
C147 drain_left.n10 a_n1882_n3888# 0.883863f
C148 drain_left.t7 a_n1882_n3888# 0.463848f
C149 drain_left.t12 a_n1882_n3888# 0.463848f
C150 drain_left.n11 a_n1882_n3888# 4.19265f
C151 drain_left.n12 a_n1882_n3888# 0.435732f
C152 drain_left.t15 a_n1882_n3888# 0.463848f
C153 drain_left.t2 a_n1882_n3888# 0.463848f
C154 drain_left.n13 a_n1882_n3888# 4.19265f
C155 drain_left.n14 a_n1882_n3888# 0.435732f
C156 drain_left.t9 a_n1882_n3888# 0.463848f
C157 drain_left.t13 a_n1882_n3888# 0.463848f
C158 drain_left.n15 a_n1882_n3888# 4.19264f
C159 drain_left.n16 a_n1882_n3888# 0.756005f
C160 source.t20 a_n1882_n3888# 4.44078f
C161 source.n0 a_n1882_n3888# 2.0419f
C162 source.t35 a_n1882_n3888# 0.396264f
C163 source.t34 a_n1882_n3888# 0.396264f
C164 source.n1 a_n1882_n3888# 3.48085f
C165 source.n2 a_n1882_n3888# 0.427726f
C166 source.t22 a_n1882_n3888# 0.396264f
C167 source.t24 a_n1882_n3888# 0.396264f
C168 source.n3 a_n1882_n3888# 3.48085f
C169 source.n4 a_n1882_n3888# 0.427726f
C170 source.t30 a_n1882_n3888# 0.396264f
C171 source.t29 a_n1882_n3888# 0.396264f
C172 source.n5 a_n1882_n3888# 3.48085f
C173 source.n6 a_n1882_n3888# 0.427726f
C174 source.t31 a_n1882_n3888# 0.396264f
C175 source.t27 a_n1882_n3888# 0.396264f
C176 source.n7 a_n1882_n3888# 3.48085f
C177 source.n8 a_n1882_n3888# 0.427726f
C178 source.t33 a_n1882_n3888# 4.44078f
C179 source.n9 a_n1882_n3888# 0.549904f
C180 source.t38 a_n1882_n3888# 4.44078f
C181 source.n10 a_n1882_n3888# 0.549904f
C182 source.t12 a_n1882_n3888# 0.396264f
C183 source.t7 a_n1882_n3888# 0.396264f
C184 source.n11 a_n1882_n3888# 3.48085f
C185 source.n12 a_n1882_n3888# 0.427726f
C186 source.t39 a_n1882_n3888# 0.396264f
C187 source.t4 a_n1882_n3888# 0.396264f
C188 source.n13 a_n1882_n3888# 3.48085f
C189 source.n14 a_n1882_n3888# 0.427726f
C190 source.t15 a_n1882_n3888# 0.396264f
C191 source.t9 a_n1882_n3888# 0.396264f
C192 source.n15 a_n1882_n3888# 3.48085f
C193 source.n16 a_n1882_n3888# 0.427726f
C194 source.t16 a_n1882_n3888# 0.396264f
C195 source.t14 a_n1882_n3888# 0.396264f
C196 source.n17 a_n1882_n3888# 3.48085f
C197 source.n18 a_n1882_n3888# 0.427726f
C198 source.t3 a_n1882_n3888# 4.44078f
C199 source.n19 a_n1882_n3888# 2.59411f
C200 source.t32 a_n1882_n3888# 4.44078f
C201 source.n20 a_n1882_n3888# 2.59412f
C202 source.t18 a_n1882_n3888# 0.396264f
C203 source.t23 a_n1882_n3888# 0.396264f
C204 source.n21 a_n1882_n3888# 3.48084f
C205 source.n22 a_n1882_n3888# 0.42773f
C206 source.t26 a_n1882_n3888# 0.396264f
C207 source.t19 a_n1882_n3888# 0.396264f
C208 source.n23 a_n1882_n3888# 3.48084f
C209 source.n24 a_n1882_n3888# 0.42773f
C210 source.t28 a_n1882_n3888# 0.396264f
C211 source.t21 a_n1882_n3888# 0.396264f
C212 source.n25 a_n1882_n3888# 3.48084f
C213 source.n26 a_n1882_n3888# 0.42773f
C214 source.t37 a_n1882_n3888# 0.396264f
C215 source.t25 a_n1882_n3888# 0.396264f
C216 source.n27 a_n1882_n3888# 3.48084f
C217 source.n28 a_n1882_n3888# 0.42773f
C218 source.t36 a_n1882_n3888# 4.44078f
C219 source.n29 a_n1882_n3888# 0.549909f
C220 source.t1 a_n1882_n3888# 4.44078f
C221 source.n30 a_n1882_n3888# 0.549909f
C222 source.t6 a_n1882_n3888# 0.396264f
C223 source.t11 a_n1882_n3888# 0.396264f
C224 source.n31 a_n1882_n3888# 3.48084f
C225 source.n32 a_n1882_n3888# 0.42773f
C226 source.t2 a_n1882_n3888# 0.396264f
C227 source.t0 a_n1882_n3888# 0.396264f
C228 source.n33 a_n1882_n3888# 3.48084f
C229 source.n34 a_n1882_n3888# 0.42773f
C230 source.t13 a_n1882_n3888# 0.396264f
C231 source.t5 a_n1882_n3888# 0.396264f
C232 source.n35 a_n1882_n3888# 3.48084f
C233 source.n36 a_n1882_n3888# 0.42773f
C234 source.t10 a_n1882_n3888# 0.396264f
C235 source.t17 a_n1882_n3888# 0.396264f
C236 source.n37 a_n1882_n3888# 3.48084f
C237 source.n38 a_n1882_n3888# 0.42773f
C238 source.t8 a_n1882_n3888# 4.44078f
C239 source.n39 a_n1882_n3888# 0.731178f
C240 source.n40 a_n1882_n3888# 2.43894f
C241 plus.n0 a_n1882_n3888# 0.053666f
C242 plus.t10 a_n1882_n3888# 0.454201f
C243 plus.t17 a_n1882_n3888# 0.454201f
C244 plus.t4 a_n1882_n3888# 0.454201f
C245 plus.n1 a_n1882_n3888# 0.179976f
C246 plus.n2 a_n1882_n3888# 0.053666f
C247 plus.t7 a_n1882_n3888# 0.454201f
C248 plus.t12 a_n1882_n3888# 0.454201f
C249 plus.t13 a_n1882_n3888# 0.454201f
C250 plus.n3 a_n1882_n3888# 0.179976f
C251 plus.n4 a_n1882_n3888# 0.122802f
C252 plus.t18 a_n1882_n3888# 0.454201f
C253 plus.t5 a_n1882_n3888# 0.454201f
C254 plus.t8 a_n1882_n3888# 0.459288f
C255 plus.n5 a_n1882_n3888# 0.196577f
C256 plus.n6 a_n1882_n3888# 0.179976f
C257 plus.n7 a_n1882_n3888# 0.018795f
C258 plus.n8 a_n1882_n3888# 0.179976f
C259 plus.n9 a_n1882_n3888# 0.018795f
C260 plus.n10 a_n1882_n3888# 0.053666f
C261 plus.n11 a_n1882_n3888# 0.053666f
C262 plus.n12 a_n1882_n3888# 0.018795f
C263 plus.n13 a_n1882_n3888# 0.179976f
C264 plus.n14 a_n1882_n3888# 0.018795f
C265 plus.n15 a_n1882_n3888# 0.179976f
C266 plus.n16 a_n1882_n3888# 0.018795f
C267 plus.n17 a_n1882_n3888# 0.053666f
C268 plus.n18 a_n1882_n3888# 0.053666f
C269 plus.n19 a_n1882_n3888# 0.018795f
C270 plus.n20 a_n1882_n3888# 0.179976f
C271 plus.n21 a_n1882_n3888# 0.018795f
C272 plus.n22 a_n1882_n3888# 0.179976f
C273 plus.t6 a_n1882_n3888# 0.459288f
C274 plus.n23 a_n1882_n3888# 0.196496f
C275 plus.n24 a_n1882_n3888# 0.675358f
C276 plus.n25 a_n1882_n3888# 0.053666f
C277 plus.t9 a_n1882_n3888# 0.459288f
C278 plus.t11 a_n1882_n3888# 0.454201f
C279 plus.t14 a_n1882_n3888# 0.454201f
C280 plus.t19 a_n1882_n3888# 0.454201f
C281 plus.n26 a_n1882_n3888# 0.179976f
C282 plus.n27 a_n1882_n3888# 0.053666f
C283 plus.t16 a_n1882_n3888# 0.454201f
C284 plus.t0 a_n1882_n3888# 0.454201f
C285 plus.t15 a_n1882_n3888# 0.454201f
C286 plus.n28 a_n1882_n3888# 0.179976f
C287 plus.n29 a_n1882_n3888# 0.122802f
C288 plus.t1 a_n1882_n3888# 0.454201f
C289 plus.t3 a_n1882_n3888# 0.454201f
C290 plus.t2 a_n1882_n3888# 0.459288f
C291 plus.n30 a_n1882_n3888# 0.196577f
C292 plus.n31 a_n1882_n3888# 0.179976f
C293 plus.n32 a_n1882_n3888# 0.018795f
C294 plus.n33 a_n1882_n3888# 0.179976f
C295 plus.n34 a_n1882_n3888# 0.018795f
C296 plus.n35 a_n1882_n3888# 0.053666f
C297 plus.n36 a_n1882_n3888# 0.053666f
C298 plus.n37 a_n1882_n3888# 0.018795f
C299 plus.n38 a_n1882_n3888# 0.179976f
C300 plus.n39 a_n1882_n3888# 0.018795f
C301 plus.n40 a_n1882_n3888# 0.179976f
C302 plus.n41 a_n1882_n3888# 0.018795f
C303 plus.n42 a_n1882_n3888# 0.053666f
C304 plus.n43 a_n1882_n3888# 0.053666f
C305 plus.n44 a_n1882_n3888# 0.018795f
C306 plus.n45 a_n1882_n3888# 0.179976f
C307 plus.n46 a_n1882_n3888# 0.018795f
C308 plus.n47 a_n1882_n3888# 0.179976f
C309 plus.n48 a_n1882_n3888# 0.196496f
C310 plus.n49 a_n1882_n3888# 1.71602f
.ends

