* NGSPICE file created from diffpair359.ext - technology: sky130A

.subckt diffpair359 minus drain_right drain_left source plus
X0 source.t47 plus.t0 drain_left.t15 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X1 drain_left.t7 plus.t1 source.t46 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X2 source.t0 minus.t0 drain_right.t23 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X3 drain_left.t23 plus.t2 source.t45 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X4 drain_left.t10 plus.t3 source.t44 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X5 drain_right.t22 minus.t1 source.t15 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X6 drain_right.t21 minus.t2 source.t19 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X7 source.t23 minus.t3 drain_right.t20 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X8 source.t43 plus.t4 drain_left.t9 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X9 source.t16 minus.t4 drain_right.t19 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X10 source.t1 minus.t5 drain_right.t18 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X11 a_n2354_n2688# a_n2354_n2688# a_n2354_n2688# a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.3
X12 drain_left.t17 plus.t5 source.t42 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X13 a_n2354_n2688# a_n2354_n2688# a_n2354_n2688# a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X14 drain_right.t17 minus.t6 source.t5 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X15 source.t6 minus.t7 drain_right.t16 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X16 drain_left.t18 plus.t6 source.t41 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X17 source.t11 minus.t8 drain_right.t15 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X18 source.t40 plus.t7 drain_left.t22 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X19 source.t39 plus.t8 drain_left.t8 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X20 source.t38 plus.t9 drain_left.t16 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X21 source.t37 plus.t10 drain_left.t14 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X22 drain_left.t6 plus.t11 source.t36 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X23 drain_right.t14 minus.t9 source.t8 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X24 drain_right.t13 minus.t10 source.t2 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X25 source.t10 minus.t11 drain_right.t12 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X26 a_n2354_n2688# a_n2354_n2688# a_n2354_n2688# a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X27 source.t13 minus.t12 drain_right.t11 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X28 source.t35 plus.t12 drain_left.t21 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X29 drain_right.t10 minus.t13 source.t18 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X30 drain_right.t9 minus.t14 source.t20 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X31 source.t34 plus.t13 drain_left.t20 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X32 source.t33 plus.t14 drain_left.t19 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X33 drain_right.t8 minus.t15 source.t12 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X34 drain_left.t13 plus.t15 source.t32 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X35 drain_left.t5 plus.t16 source.t31 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X36 source.t30 plus.t17 drain_left.t0 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X37 drain_left.t3 plus.t18 source.t29 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X38 drain_left.t2 plus.t19 source.t28 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X39 drain_right.t7 minus.t16 source.t17 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X40 drain_right.t6 minus.t17 source.t21 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X41 a_n2354_n2688# a_n2354_n2688# a_n2354_n2688# a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X42 source.t22 minus.t18 drain_right.t5 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X43 source.t4 minus.t19 drain_right.t4 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X44 source.t9 minus.t20 drain_right.t3 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X45 source.t3 minus.t21 drain_right.t2 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X46 source.t27 plus.t20 drain_left.t12 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X47 drain_right.t1 minus.t22 source.t7 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X48 drain_right.t0 minus.t23 source.t14 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X49 source.t26 plus.t21 drain_left.t1 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X50 drain_left.t11 plus.t22 source.t25 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X51 drain_left.t4 plus.t23 source.t24 a_n2354_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
R0 plus.n9 plus.t4 858.837
R1 plus.n35 plus.t5 858.837
R2 plus.n46 plus.t16 858.837
R3 plus.n72 plus.t21 858.837
R4 plus.n8 plus.t11 827.433
R5 plus.n13 plus.t17 827.433
R6 plus.n15 plus.t22 827.433
R7 plus.n5 plus.t8 827.433
R8 plus.n20 plus.t15 827.433
R9 plus.n3 plus.t20 827.433
R10 plus.n26 plus.t1 827.433
R11 plus.n28 plus.t12 827.433
R12 plus.n1 plus.t19 827.433
R13 plus.n34 plus.t0 827.433
R14 plus.n45 plus.t7 827.433
R15 plus.n50 plus.t18 827.433
R16 plus.n52 plus.t9 827.433
R17 plus.n42 plus.t2 827.433
R18 plus.n57 plus.t10 827.433
R19 plus.n40 plus.t3 827.433
R20 plus.n63 plus.t13 827.433
R21 plus.n65 plus.t23 827.433
R22 plus.n38 plus.t14 827.433
R23 plus.n71 plus.t6 827.433
R24 plus.n10 plus.n9 161.489
R25 plus.n47 plus.n46 161.489
R26 plus.n10 plus.n7 161.3
R27 plus.n12 plus.n11 161.3
R28 plus.n14 plus.n6 161.3
R29 plus.n17 plus.n16 161.3
R30 plus.n19 plus.n18 161.3
R31 plus.n21 plus.n4 161.3
R32 plus.n23 plus.n22 161.3
R33 plus.n25 plus.n24 161.3
R34 plus.n27 plus.n2 161.3
R35 plus.n30 plus.n29 161.3
R36 plus.n32 plus.n31 161.3
R37 plus.n33 plus.n0 161.3
R38 plus.n36 plus.n35 161.3
R39 plus.n47 plus.n44 161.3
R40 plus.n49 plus.n48 161.3
R41 plus.n51 plus.n43 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n56 plus.n55 161.3
R44 plus.n58 plus.n41 161.3
R45 plus.n60 plus.n59 161.3
R46 plus.n62 plus.n61 161.3
R47 plus.n64 plus.n39 161.3
R48 plus.n67 plus.n66 161.3
R49 plus.n69 plus.n68 161.3
R50 plus.n70 plus.n37 161.3
R51 plus.n73 plus.n72 161.3
R52 plus.n12 plus.n7 73.0308
R53 plus.n22 plus.n21 73.0308
R54 plus.n33 plus.n32 73.0308
R55 plus.n70 plus.n69 73.0308
R56 plus.n59 plus.n58 73.0308
R57 plus.n49 plus.n44 73.0308
R58 plus.n14 plus.n13 66.4581
R59 plus.n29 plus.n1 66.4581
R60 plus.n66 plus.n38 66.4581
R61 plus.n51 plus.n50 66.4581
R62 plus.n20 plus.n19 63.5369
R63 plus.n25 plus.n3 63.5369
R64 plus.n62 plus.n40 63.5369
R65 plus.n57 plus.n56 63.5369
R66 plus.n9 plus.n8 60.6157
R67 plus.n35 plus.n34 60.6157
R68 plus.n72 plus.n71 60.6157
R69 plus.n46 plus.n45 60.6157
R70 plus.n16 plus.n15 47.4702
R71 plus.n28 plus.n27 47.4702
R72 plus.n65 plus.n64 47.4702
R73 plus.n53 plus.n52 47.4702
R74 plus.n16 plus.n5 44.549
R75 plus.n27 plus.n26 44.549
R76 plus.n64 plus.n63 44.549
R77 plus.n53 plus.n42 44.549
R78 plus plus.n73 30.7528
R79 plus.n19 plus.n5 28.4823
R80 plus.n26 plus.n25 28.4823
R81 plus.n63 plus.n62 28.4823
R82 plus.n56 plus.n42 28.4823
R83 plus.n15 plus.n14 25.5611
R84 plus.n29 plus.n28 25.5611
R85 plus.n66 plus.n65 25.5611
R86 plus.n52 plus.n51 25.5611
R87 plus.n8 plus.n7 12.4157
R88 plus.n34 plus.n33 12.4157
R89 plus.n71 plus.n70 12.4157
R90 plus.n45 plus.n44 12.4157
R91 plus plus.n36 10.9778
R92 plus.n21 plus.n20 9.49444
R93 plus.n22 plus.n3 9.49444
R94 plus.n59 plus.n40 9.49444
R95 plus.n58 plus.n57 9.49444
R96 plus.n13 plus.n12 6.57323
R97 plus.n32 plus.n1 6.57323
R98 plus.n69 plus.n38 6.57323
R99 plus.n50 plus.n49 6.57323
R100 plus.n11 plus.n10 0.189894
R101 plus.n11 plus.n6 0.189894
R102 plus.n17 plus.n6 0.189894
R103 plus.n18 plus.n17 0.189894
R104 plus.n18 plus.n4 0.189894
R105 plus.n23 plus.n4 0.189894
R106 plus.n24 plus.n23 0.189894
R107 plus.n24 plus.n2 0.189894
R108 plus.n30 plus.n2 0.189894
R109 plus.n31 plus.n30 0.189894
R110 plus.n31 plus.n0 0.189894
R111 plus.n36 plus.n0 0.189894
R112 plus.n73 plus.n37 0.189894
R113 plus.n68 plus.n37 0.189894
R114 plus.n68 plus.n67 0.189894
R115 plus.n67 plus.n39 0.189894
R116 plus.n61 plus.n39 0.189894
R117 plus.n61 plus.n60 0.189894
R118 plus.n60 plus.n41 0.189894
R119 plus.n55 plus.n41 0.189894
R120 plus.n55 plus.n54 0.189894
R121 plus.n54 plus.n43 0.189894
R122 plus.n48 plus.n43 0.189894
R123 plus.n48 plus.n47 0.189894
R124 drain_left.n13 drain_left.n11 66.0807
R125 drain_left.n7 drain_left.n5 66.0804
R126 drain_left.n2 drain_left.n0 66.0804
R127 drain_left.n19 drain_left.n18 65.5376
R128 drain_left.n17 drain_left.n16 65.5376
R129 drain_left.n15 drain_left.n14 65.5376
R130 drain_left.n13 drain_left.n12 65.5376
R131 drain_left.n21 drain_left.n20 65.5374
R132 drain_left.n7 drain_left.n6 65.5373
R133 drain_left.n9 drain_left.n8 65.5373
R134 drain_left.n4 drain_left.n3 65.5373
R135 drain_left.n2 drain_left.n1 65.5373
R136 drain_left drain_left.n10 30.2538
R137 drain_left drain_left.n21 6.19632
R138 drain_left.n5 drain_left.t22 2.2005
R139 drain_left.n5 drain_left.t5 2.2005
R140 drain_left.n6 drain_left.t16 2.2005
R141 drain_left.n6 drain_left.t3 2.2005
R142 drain_left.n8 drain_left.t14 2.2005
R143 drain_left.n8 drain_left.t23 2.2005
R144 drain_left.n3 drain_left.t20 2.2005
R145 drain_left.n3 drain_left.t10 2.2005
R146 drain_left.n1 drain_left.t19 2.2005
R147 drain_left.n1 drain_left.t4 2.2005
R148 drain_left.n0 drain_left.t1 2.2005
R149 drain_left.n0 drain_left.t18 2.2005
R150 drain_left.n20 drain_left.t15 2.2005
R151 drain_left.n20 drain_left.t17 2.2005
R152 drain_left.n18 drain_left.t21 2.2005
R153 drain_left.n18 drain_left.t2 2.2005
R154 drain_left.n16 drain_left.t12 2.2005
R155 drain_left.n16 drain_left.t7 2.2005
R156 drain_left.n14 drain_left.t8 2.2005
R157 drain_left.n14 drain_left.t13 2.2005
R158 drain_left.n12 drain_left.t0 2.2005
R159 drain_left.n12 drain_left.t11 2.2005
R160 drain_left.n11 drain_left.t9 2.2005
R161 drain_left.n11 drain_left.t6 2.2005
R162 drain_left.n9 drain_left.n7 0.543603
R163 drain_left.n4 drain_left.n2 0.543603
R164 drain_left.n15 drain_left.n13 0.543603
R165 drain_left.n17 drain_left.n15 0.543603
R166 drain_left.n19 drain_left.n17 0.543603
R167 drain_left.n21 drain_left.n19 0.543603
R168 drain_left.n10 drain_left.n9 0.216706
R169 drain_left.n10 drain_left.n4 0.216706
R170 source.n11 source.t43 51.0588
R171 source.n12 source.t12 51.0588
R172 source.n23 source.t23 51.0588
R173 source.n47 source.t7 51.0586
R174 source.n36 source.t3 51.0586
R175 source.n35 source.t31 51.0586
R176 source.n24 source.t26 51.0586
R177 source.n0 source.t42 51.0586
R178 source.n2 source.n1 48.8588
R179 source.n4 source.n3 48.8588
R180 source.n6 source.n5 48.8588
R181 source.n8 source.n7 48.8588
R182 source.n10 source.n9 48.8588
R183 source.n14 source.n13 48.8588
R184 source.n16 source.n15 48.8588
R185 source.n18 source.n17 48.8588
R186 source.n20 source.n19 48.8588
R187 source.n22 source.n21 48.8588
R188 source.n46 source.n45 48.8586
R189 source.n44 source.n43 48.8586
R190 source.n42 source.n41 48.8586
R191 source.n40 source.n39 48.8586
R192 source.n38 source.n37 48.8586
R193 source.n34 source.n33 48.8586
R194 source.n32 source.n31 48.8586
R195 source.n30 source.n29 48.8586
R196 source.n28 source.n27 48.8586
R197 source.n26 source.n25 48.8586
R198 source.n24 source.n23 19.5581
R199 source.n48 source.n0 14.0236
R200 source.n48 source.n47 5.53498
R201 source.n45 source.t14 2.2005
R202 source.n45 source.t6 2.2005
R203 source.n43 source.t18 2.2005
R204 source.n43 source.t13 2.2005
R205 source.n41 source.t20 2.2005
R206 source.n41 source.t16 2.2005
R207 source.n39 source.t8 2.2005
R208 source.n39 source.t1 2.2005
R209 source.n37 source.t2 2.2005
R210 source.n37 source.t9 2.2005
R211 source.n33 source.t29 2.2005
R212 source.n33 source.t40 2.2005
R213 source.n31 source.t45 2.2005
R214 source.n31 source.t38 2.2005
R215 source.n29 source.t44 2.2005
R216 source.n29 source.t37 2.2005
R217 source.n27 source.t24 2.2005
R218 source.n27 source.t34 2.2005
R219 source.n25 source.t41 2.2005
R220 source.n25 source.t33 2.2005
R221 source.n1 source.t28 2.2005
R222 source.n1 source.t47 2.2005
R223 source.n3 source.t46 2.2005
R224 source.n3 source.t35 2.2005
R225 source.n5 source.t32 2.2005
R226 source.n5 source.t27 2.2005
R227 source.n7 source.t25 2.2005
R228 source.n7 source.t39 2.2005
R229 source.n9 source.t36 2.2005
R230 source.n9 source.t30 2.2005
R231 source.n13 source.t15 2.2005
R232 source.n13 source.t22 2.2005
R233 source.n15 source.t17 2.2005
R234 source.n15 source.t10 2.2005
R235 source.n17 source.t5 2.2005
R236 source.n17 source.t0 2.2005
R237 source.n19 source.t19 2.2005
R238 source.n19 source.t4 2.2005
R239 source.n21 source.t21 2.2005
R240 source.n21 source.t11 2.2005
R241 source.n23 source.n22 0.543603
R242 source.n22 source.n20 0.543603
R243 source.n20 source.n18 0.543603
R244 source.n18 source.n16 0.543603
R245 source.n16 source.n14 0.543603
R246 source.n14 source.n12 0.543603
R247 source.n11 source.n10 0.543603
R248 source.n10 source.n8 0.543603
R249 source.n8 source.n6 0.543603
R250 source.n6 source.n4 0.543603
R251 source.n4 source.n2 0.543603
R252 source.n2 source.n0 0.543603
R253 source.n26 source.n24 0.543603
R254 source.n28 source.n26 0.543603
R255 source.n30 source.n28 0.543603
R256 source.n32 source.n30 0.543603
R257 source.n34 source.n32 0.543603
R258 source.n35 source.n34 0.543603
R259 source.n38 source.n36 0.543603
R260 source.n40 source.n38 0.543603
R261 source.n42 source.n40 0.543603
R262 source.n44 source.n42 0.543603
R263 source.n46 source.n44 0.543603
R264 source.n47 source.n46 0.543603
R265 source.n12 source.n11 0.470328
R266 source.n36 source.n35 0.470328
R267 source source.n48 0.188
R268 minus.n35 minus.t3 858.837
R269 minus.n9 minus.t15 858.837
R270 minus.n72 minus.t22 858.837
R271 minus.n46 minus.t21 858.837
R272 minus.n34 minus.t17 827.433
R273 minus.n1 minus.t8 827.433
R274 minus.n28 minus.t2 827.433
R275 minus.n26 minus.t19 827.433
R276 minus.n3 minus.t6 827.433
R277 minus.n20 minus.t0 827.433
R278 minus.n5 minus.t16 827.433
R279 minus.n15 minus.t11 827.433
R280 minus.n13 minus.t1 827.433
R281 minus.n8 minus.t18 827.433
R282 minus.n71 minus.t7 827.433
R283 minus.n38 minus.t23 827.433
R284 minus.n65 minus.t12 827.433
R285 minus.n63 minus.t13 827.433
R286 minus.n40 minus.t4 827.433
R287 minus.n57 minus.t14 827.433
R288 minus.n42 minus.t5 827.433
R289 minus.n52 minus.t9 827.433
R290 minus.n50 minus.t20 827.433
R291 minus.n45 minus.t10 827.433
R292 minus.n10 minus.n9 161.489
R293 minus.n47 minus.n46 161.489
R294 minus.n36 minus.n35 161.3
R295 minus.n33 minus.n0 161.3
R296 minus.n32 minus.n31 161.3
R297 minus.n30 minus.n29 161.3
R298 minus.n27 minus.n2 161.3
R299 minus.n25 minus.n24 161.3
R300 minus.n23 minus.n22 161.3
R301 minus.n21 minus.n4 161.3
R302 minus.n19 minus.n18 161.3
R303 minus.n17 minus.n16 161.3
R304 minus.n14 minus.n6 161.3
R305 minus.n12 minus.n11 161.3
R306 minus.n10 minus.n7 161.3
R307 minus.n73 minus.n72 161.3
R308 minus.n70 minus.n37 161.3
R309 minus.n69 minus.n68 161.3
R310 minus.n67 minus.n66 161.3
R311 minus.n64 minus.n39 161.3
R312 minus.n62 minus.n61 161.3
R313 minus.n60 minus.n59 161.3
R314 minus.n58 minus.n41 161.3
R315 minus.n56 minus.n55 161.3
R316 minus.n54 minus.n53 161.3
R317 minus.n51 minus.n43 161.3
R318 minus.n49 minus.n48 161.3
R319 minus.n47 minus.n44 161.3
R320 minus.n33 minus.n32 73.0308
R321 minus.n22 minus.n21 73.0308
R322 minus.n12 minus.n7 73.0308
R323 minus.n49 minus.n44 73.0308
R324 minus.n59 minus.n58 73.0308
R325 minus.n70 minus.n69 73.0308
R326 minus.n29 minus.n1 66.4581
R327 minus.n14 minus.n13 66.4581
R328 minus.n51 minus.n50 66.4581
R329 minus.n66 minus.n38 66.4581
R330 minus.n25 minus.n3 63.5369
R331 minus.n20 minus.n19 63.5369
R332 minus.n57 minus.n56 63.5369
R333 minus.n62 minus.n40 63.5369
R334 minus.n35 minus.n34 60.6157
R335 minus.n9 minus.n8 60.6157
R336 minus.n46 minus.n45 60.6157
R337 minus.n72 minus.n71 60.6157
R338 minus.n28 minus.n27 47.4702
R339 minus.n16 minus.n15 47.4702
R340 minus.n53 minus.n52 47.4702
R341 minus.n65 minus.n64 47.4702
R342 minus.n27 minus.n26 44.549
R343 minus.n16 minus.n5 44.549
R344 minus.n53 minus.n42 44.549
R345 minus.n64 minus.n63 44.549
R346 minus.n74 minus.n36 35.7354
R347 minus.n26 minus.n25 28.4823
R348 minus.n19 minus.n5 28.4823
R349 minus.n56 minus.n42 28.4823
R350 minus.n63 minus.n62 28.4823
R351 minus.n29 minus.n28 25.5611
R352 minus.n15 minus.n14 25.5611
R353 minus.n52 minus.n51 25.5611
R354 minus.n66 minus.n65 25.5611
R355 minus.n34 minus.n33 12.4157
R356 minus.n8 minus.n7 12.4157
R357 minus.n45 minus.n44 12.4157
R358 minus.n71 minus.n70 12.4157
R359 minus.n22 minus.n3 9.49444
R360 minus.n21 minus.n20 9.49444
R361 minus.n58 minus.n57 9.49444
R362 minus.n59 minus.n40 9.49444
R363 minus.n32 minus.n1 6.57323
R364 minus.n13 minus.n12 6.57323
R365 minus.n50 minus.n49 6.57323
R366 minus.n69 minus.n38 6.57323
R367 minus.n74 minus.n73 6.4702
R368 minus.n36 minus.n0 0.189894
R369 minus.n31 minus.n0 0.189894
R370 minus.n31 minus.n30 0.189894
R371 minus.n30 minus.n2 0.189894
R372 minus.n24 minus.n2 0.189894
R373 minus.n24 minus.n23 0.189894
R374 minus.n23 minus.n4 0.189894
R375 minus.n18 minus.n4 0.189894
R376 minus.n18 minus.n17 0.189894
R377 minus.n17 minus.n6 0.189894
R378 minus.n11 minus.n6 0.189894
R379 minus.n11 minus.n10 0.189894
R380 minus.n48 minus.n47 0.189894
R381 minus.n48 minus.n43 0.189894
R382 minus.n54 minus.n43 0.189894
R383 minus.n55 minus.n54 0.189894
R384 minus.n55 minus.n41 0.189894
R385 minus.n60 minus.n41 0.189894
R386 minus.n61 minus.n60 0.189894
R387 minus.n61 minus.n39 0.189894
R388 minus.n67 minus.n39 0.189894
R389 minus.n68 minus.n67 0.189894
R390 minus.n68 minus.n37 0.189894
R391 minus.n73 minus.n37 0.189894
R392 minus minus.n74 0.188
R393 drain_right.n13 drain_right.n11 66.0805
R394 drain_right.n7 drain_right.n5 66.0804
R395 drain_right.n2 drain_right.n0 66.0804
R396 drain_right.n13 drain_right.n12 65.5376
R397 drain_right.n15 drain_right.n14 65.5376
R398 drain_right.n17 drain_right.n16 65.5376
R399 drain_right.n19 drain_right.n18 65.5376
R400 drain_right.n21 drain_right.n20 65.5376
R401 drain_right.n7 drain_right.n6 65.5373
R402 drain_right.n9 drain_right.n8 65.5373
R403 drain_right.n4 drain_right.n3 65.5373
R404 drain_right.n2 drain_right.n1 65.5373
R405 drain_right drain_right.n10 29.7006
R406 drain_right drain_right.n21 6.19632
R407 drain_right.n5 drain_right.t16 2.2005
R408 drain_right.n5 drain_right.t1 2.2005
R409 drain_right.n6 drain_right.t11 2.2005
R410 drain_right.n6 drain_right.t0 2.2005
R411 drain_right.n8 drain_right.t19 2.2005
R412 drain_right.n8 drain_right.t10 2.2005
R413 drain_right.n3 drain_right.t18 2.2005
R414 drain_right.n3 drain_right.t9 2.2005
R415 drain_right.n1 drain_right.t3 2.2005
R416 drain_right.n1 drain_right.t14 2.2005
R417 drain_right.n0 drain_right.t2 2.2005
R418 drain_right.n0 drain_right.t13 2.2005
R419 drain_right.n11 drain_right.t5 2.2005
R420 drain_right.n11 drain_right.t8 2.2005
R421 drain_right.n12 drain_right.t12 2.2005
R422 drain_right.n12 drain_right.t22 2.2005
R423 drain_right.n14 drain_right.t23 2.2005
R424 drain_right.n14 drain_right.t7 2.2005
R425 drain_right.n16 drain_right.t4 2.2005
R426 drain_right.n16 drain_right.t17 2.2005
R427 drain_right.n18 drain_right.t15 2.2005
R428 drain_right.n18 drain_right.t21 2.2005
R429 drain_right.n20 drain_right.t20 2.2005
R430 drain_right.n20 drain_right.t6 2.2005
R431 drain_right.n9 drain_right.n7 0.543603
R432 drain_right.n4 drain_right.n2 0.543603
R433 drain_right.n21 drain_right.n19 0.543603
R434 drain_right.n19 drain_right.n17 0.543603
R435 drain_right.n17 drain_right.n15 0.543603
R436 drain_right.n15 drain_right.n13 0.543603
R437 drain_right.n10 drain_right.n9 0.216706
R438 drain_right.n10 drain_right.n4 0.216706
C0 drain_left plus 6.72734f
C1 plus drain_right 0.387992f
C2 drain_left drain_right 1.26597f
C3 plus minus 5.53846f
C4 drain_left minus 0.172624f
C5 drain_right minus 6.49513f
C6 plus source 6.44954f
C7 drain_left source 34.2775f
C8 drain_right source 34.278103f
C9 minus source 6.4355f
C10 drain_right a_n2354_n2688# 6.70327f
C11 drain_left a_n2354_n2688# 7.05467f
C12 source a_n2354_n2688# 7.313262f
C13 minus a_n2354_n2688# 9.075839f
C14 plus a_n2354_n2688# 10.927509f
C15 drain_right.t2 a_n2354_n2688# 0.242175f
C16 drain_right.t13 a_n2354_n2688# 0.242175f
C17 drain_right.n0 a_n2354_n2688# 2.12155f
C18 drain_right.t3 a_n2354_n2688# 0.242175f
C19 drain_right.t14 a_n2354_n2688# 0.242175f
C20 drain_right.n1 a_n2354_n2688# 2.11822f
C21 drain_right.n2 a_n2354_n2688# 0.794247f
C22 drain_right.t18 a_n2354_n2688# 0.242175f
C23 drain_right.t9 a_n2354_n2688# 0.242175f
C24 drain_right.n3 a_n2354_n2688# 2.11822f
C25 drain_right.n4 a_n2354_n2688# 0.359717f
C26 drain_right.t16 a_n2354_n2688# 0.242175f
C27 drain_right.t1 a_n2354_n2688# 0.242175f
C28 drain_right.n5 a_n2354_n2688# 2.12155f
C29 drain_right.t11 a_n2354_n2688# 0.242175f
C30 drain_right.t0 a_n2354_n2688# 0.242175f
C31 drain_right.n6 a_n2354_n2688# 2.11822f
C32 drain_right.n7 a_n2354_n2688# 0.794247f
C33 drain_right.t19 a_n2354_n2688# 0.242175f
C34 drain_right.t10 a_n2354_n2688# 0.242175f
C35 drain_right.n8 a_n2354_n2688# 2.11822f
C36 drain_right.n9 a_n2354_n2688# 0.359717f
C37 drain_right.n10 a_n2354_n2688# 1.54684f
C38 drain_right.t5 a_n2354_n2688# 0.242175f
C39 drain_right.t8 a_n2354_n2688# 0.242175f
C40 drain_right.n11 a_n2354_n2688# 2.12155f
C41 drain_right.t12 a_n2354_n2688# 0.242175f
C42 drain_right.t22 a_n2354_n2688# 0.242175f
C43 drain_right.n12 a_n2354_n2688# 2.11822f
C44 drain_right.n13 a_n2354_n2688# 0.794248f
C45 drain_right.t23 a_n2354_n2688# 0.242175f
C46 drain_right.t7 a_n2354_n2688# 0.242175f
C47 drain_right.n14 a_n2354_n2688# 2.11822f
C48 drain_right.n15 a_n2354_n2688# 0.391929f
C49 drain_right.t4 a_n2354_n2688# 0.242175f
C50 drain_right.t17 a_n2354_n2688# 0.242175f
C51 drain_right.n16 a_n2354_n2688# 2.11822f
C52 drain_right.n17 a_n2354_n2688# 0.391929f
C53 drain_right.t15 a_n2354_n2688# 0.242175f
C54 drain_right.t21 a_n2354_n2688# 0.242175f
C55 drain_right.n18 a_n2354_n2688# 2.11822f
C56 drain_right.n19 a_n2354_n2688# 0.391929f
C57 drain_right.t20 a_n2354_n2688# 0.242175f
C58 drain_right.t6 a_n2354_n2688# 0.242175f
C59 drain_right.n20 a_n2354_n2688# 2.11822f
C60 drain_right.n21 a_n2354_n2688# 0.675358f
C61 minus.n0 a_n2354_n2688# 0.048225f
C62 minus.t3 a_n2354_n2688# 0.37461f
C63 minus.t17 a_n2354_n2688# 0.36896f
C64 minus.t8 a_n2354_n2688# 0.36896f
C65 minus.n1 a_n2354_n2688# 0.154071f
C66 minus.n2 a_n2354_n2688# 0.048225f
C67 minus.t2 a_n2354_n2688# 0.36896f
C68 minus.t19 a_n2354_n2688# 0.36896f
C69 minus.t6 a_n2354_n2688# 0.36896f
C70 minus.n3 a_n2354_n2688# 0.154071f
C71 minus.n4 a_n2354_n2688# 0.048225f
C72 minus.t0 a_n2354_n2688# 0.36896f
C73 minus.t16 a_n2354_n2688# 0.36896f
C74 minus.n5 a_n2354_n2688# 0.154071f
C75 minus.n6 a_n2354_n2688# 0.048225f
C76 minus.t11 a_n2354_n2688# 0.36896f
C77 minus.t1 a_n2354_n2688# 0.36896f
C78 minus.n7 a_n2354_n2688# 0.018525f
C79 minus.t18 a_n2354_n2688# 0.36896f
C80 minus.n8 a_n2354_n2688# 0.154071f
C81 minus.t15 a_n2354_n2688# 0.37461f
C82 minus.n9 a_n2354_n2688# 0.168795f
C83 minus.n10 a_n2354_n2688# 0.103225f
C84 minus.n11 a_n2354_n2688# 0.048225f
C85 minus.n12 a_n2354_n2688# 0.017336f
C86 minus.n13 a_n2354_n2688# 0.154071f
C87 minus.n14 a_n2354_n2688# 0.019863f
C88 minus.n15 a_n2354_n2688# 0.154071f
C89 minus.n16 a_n2354_n2688# 0.019863f
C90 minus.n17 a_n2354_n2688# 0.048225f
C91 minus.n18 a_n2354_n2688# 0.048225f
C92 minus.n19 a_n2354_n2688# 0.019863f
C93 minus.n20 a_n2354_n2688# 0.154071f
C94 minus.n21 a_n2354_n2688# 0.017931f
C95 minus.n22 a_n2354_n2688# 0.017931f
C96 minus.n23 a_n2354_n2688# 0.048225f
C97 minus.n24 a_n2354_n2688# 0.048225f
C98 minus.n25 a_n2354_n2688# 0.019863f
C99 minus.n26 a_n2354_n2688# 0.154071f
C100 minus.n27 a_n2354_n2688# 0.019863f
C101 minus.n28 a_n2354_n2688# 0.154071f
C102 minus.n29 a_n2354_n2688# 0.019863f
C103 minus.n30 a_n2354_n2688# 0.048225f
C104 minus.n31 a_n2354_n2688# 0.048225f
C105 minus.n32 a_n2354_n2688# 0.017336f
C106 minus.n33 a_n2354_n2688# 0.018525f
C107 minus.n34 a_n2354_n2688# 0.154071f
C108 minus.n35 a_n2354_n2688# 0.168731f
C109 minus.n36 a_n2354_n2688# 1.66949f
C110 minus.n37 a_n2354_n2688# 0.048225f
C111 minus.t7 a_n2354_n2688# 0.36896f
C112 minus.t23 a_n2354_n2688# 0.36896f
C113 minus.n38 a_n2354_n2688# 0.154071f
C114 minus.n39 a_n2354_n2688# 0.048225f
C115 minus.t12 a_n2354_n2688# 0.36896f
C116 minus.t13 a_n2354_n2688# 0.36896f
C117 minus.t4 a_n2354_n2688# 0.36896f
C118 minus.n40 a_n2354_n2688# 0.154071f
C119 minus.n41 a_n2354_n2688# 0.048225f
C120 minus.t14 a_n2354_n2688# 0.36896f
C121 minus.t5 a_n2354_n2688# 0.36896f
C122 minus.n42 a_n2354_n2688# 0.154071f
C123 minus.n43 a_n2354_n2688# 0.048225f
C124 minus.t9 a_n2354_n2688# 0.36896f
C125 minus.t20 a_n2354_n2688# 0.36896f
C126 minus.n44 a_n2354_n2688# 0.018525f
C127 minus.t21 a_n2354_n2688# 0.37461f
C128 minus.t10 a_n2354_n2688# 0.36896f
C129 minus.n45 a_n2354_n2688# 0.154071f
C130 minus.n46 a_n2354_n2688# 0.168795f
C131 minus.n47 a_n2354_n2688# 0.103225f
C132 minus.n48 a_n2354_n2688# 0.048225f
C133 minus.n49 a_n2354_n2688# 0.017336f
C134 minus.n50 a_n2354_n2688# 0.154071f
C135 minus.n51 a_n2354_n2688# 0.019863f
C136 minus.n52 a_n2354_n2688# 0.154071f
C137 minus.n53 a_n2354_n2688# 0.019863f
C138 minus.n54 a_n2354_n2688# 0.048225f
C139 minus.n55 a_n2354_n2688# 0.048225f
C140 minus.n56 a_n2354_n2688# 0.019863f
C141 minus.n57 a_n2354_n2688# 0.154071f
C142 minus.n58 a_n2354_n2688# 0.017931f
C143 minus.n59 a_n2354_n2688# 0.017931f
C144 minus.n60 a_n2354_n2688# 0.048225f
C145 minus.n61 a_n2354_n2688# 0.048225f
C146 minus.n62 a_n2354_n2688# 0.019863f
C147 minus.n63 a_n2354_n2688# 0.154071f
C148 minus.n64 a_n2354_n2688# 0.019863f
C149 minus.n65 a_n2354_n2688# 0.154071f
C150 minus.n66 a_n2354_n2688# 0.019863f
C151 minus.n67 a_n2354_n2688# 0.048225f
C152 minus.n68 a_n2354_n2688# 0.048225f
C153 minus.n69 a_n2354_n2688# 0.017336f
C154 minus.n70 a_n2354_n2688# 0.018525f
C155 minus.n71 a_n2354_n2688# 0.154071f
C156 minus.t22 a_n2354_n2688# 0.37461f
C157 minus.n72 a_n2354_n2688# 0.168731f
C158 minus.n73 a_n2354_n2688# 0.311895f
C159 minus.n74 a_n2354_n2688# 2.03187f
C160 source.t42 a_n2354_n2688# 2.34191f
C161 source.n0 a_n2354_n2688# 1.34666f
C162 source.t28 a_n2354_n2688# 0.21962f
C163 source.t47 a_n2354_n2688# 0.21962f
C164 source.n1 a_n2354_n2688# 1.83851f
C165 source.n2 a_n2354_n2688# 0.395885f
C166 source.t46 a_n2354_n2688# 0.21962f
C167 source.t35 a_n2354_n2688# 0.21962f
C168 source.n3 a_n2354_n2688# 1.83851f
C169 source.n4 a_n2354_n2688# 0.395885f
C170 source.t32 a_n2354_n2688# 0.21962f
C171 source.t27 a_n2354_n2688# 0.21962f
C172 source.n5 a_n2354_n2688# 1.83851f
C173 source.n6 a_n2354_n2688# 0.395885f
C174 source.t25 a_n2354_n2688# 0.21962f
C175 source.t39 a_n2354_n2688# 0.21962f
C176 source.n7 a_n2354_n2688# 1.83851f
C177 source.n8 a_n2354_n2688# 0.395885f
C178 source.t36 a_n2354_n2688# 0.21962f
C179 source.t30 a_n2354_n2688# 0.21962f
C180 source.n9 a_n2354_n2688# 1.83851f
C181 source.n10 a_n2354_n2688# 0.395885f
C182 source.t43 a_n2354_n2688# 2.34191f
C183 source.n11 a_n2354_n2688# 0.484157f
C184 source.t12 a_n2354_n2688# 2.34191f
C185 source.n12 a_n2354_n2688# 0.484157f
C186 source.t15 a_n2354_n2688# 0.21962f
C187 source.t22 a_n2354_n2688# 0.21962f
C188 source.n13 a_n2354_n2688# 1.83851f
C189 source.n14 a_n2354_n2688# 0.395885f
C190 source.t17 a_n2354_n2688# 0.21962f
C191 source.t10 a_n2354_n2688# 0.21962f
C192 source.n15 a_n2354_n2688# 1.83851f
C193 source.n16 a_n2354_n2688# 0.395885f
C194 source.t5 a_n2354_n2688# 0.21962f
C195 source.t0 a_n2354_n2688# 0.21962f
C196 source.n17 a_n2354_n2688# 1.83851f
C197 source.n18 a_n2354_n2688# 0.395885f
C198 source.t19 a_n2354_n2688# 0.21962f
C199 source.t4 a_n2354_n2688# 0.21962f
C200 source.n19 a_n2354_n2688# 1.83851f
C201 source.n20 a_n2354_n2688# 0.395885f
C202 source.t21 a_n2354_n2688# 0.21962f
C203 source.t11 a_n2354_n2688# 0.21962f
C204 source.n21 a_n2354_n2688# 1.83851f
C205 source.n22 a_n2354_n2688# 0.395885f
C206 source.t23 a_n2354_n2688# 2.34191f
C207 source.n23 a_n2354_n2688# 1.79534f
C208 source.t26 a_n2354_n2688# 2.34191f
C209 source.n24 a_n2354_n2688# 1.79534f
C210 source.t41 a_n2354_n2688# 0.21962f
C211 source.t33 a_n2354_n2688# 0.21962f
C212 source.n25 a_n2354_n2688# 1.83851f
C213 source.n26 a_n2354_n2688# 0.395891f
C214 source.t24 a_n2354_n2688# 0.21962f
C215 source.t34 a_n2354_n2688# 0.21962f
C216 source.n27 a_n2354_n2688# 1.83851f
C217 source.n28 a_n2354_n2688# 0.395891f
C218 source.t44 a_n2354_n2688# 0.21962f
C219 source.t37 a_n2354_n2688# 0.21962f
C220 source.n29 a_n2354_n2688# 1.83851f
C221 source.n30 a_n2354_n2688# 0.395891f
C222 source.t45 a_n2354_n2688# 0.21962f
C223 source.t38 a_n2354_n2688# 0.21962f
C224 source.n31 a_n2354_n2688# 1.83851f
C225 source.n32 a_n2354_n2688# 0.395891f
C226 source.t29 a_n2354_n2688# 0.21962f
C227 source.t40 a_n2354_n2688# 0.21962f
C228 source.n33 a_n2354_n2688# 1.83851f
C229 source.n34 a_n2354_n2688# 0.395891f
C230 source.t31 a_n2354_n2688# 2.34191f
C231 source.n35 a_n2354_n2688# 0.484163f
C232 source.t3 a_n2354_n2688# 2.34191f
C233 source.n36 a_n2354_n2688# 0.484163f
C234 source.t2 a_n2354_n2688# 0.21962f
C235 source.t9 a_n2354_n2688# 0.21962f
C236 source.n37 a_n2354_n2688# 1.83851f
C237 source.n38 a_n2354_n2688# 0.395891f
C238 source.t8 a_n2354_n2688# 0.21962f
C239 source.t1 a_n2354_n2688# 0.21962f
C240 source.n39 a_n2354_n2688# 1.83851f
C241 source.n40 a_n2354_n2688# 0.395891f
C242 source.t20 a_n2354_n2688# 0.21962f
C243 source.t16 a_n2354_n2688# 0.21962f
C244 source.n41 a_n2354_n2688# 1.83851f
C245 source.n42 a_n2354_n2688# 0.395891f
C246 source.t18 a_n2354_n2688# 0.21962f
C247 source.t13 a_n2354_n2688# 0.21962f
C248 source.n43 a_n2354_n2688# 1.83851f
C249 source.n44 a_n2354_n2688# 0.395891f
C250 source.t14 a_n2354_n2688# 0.21962f
C251 source.t6 a_n2354_n2688# 0.21962f
C252 source.n45 a_n2354_n2688# 1.83851f
C253 source.n46 a_n2354_n2688# 0.395891f
C254 source.t7 a_n2354_n2688# 2.34191f
C255 source.n47 a_n2354_n2688# 0.658479f
C256 source.n48 a_n2354_n2688# 1.60751f
C257 drain_left.t1 a_n2354_n2688# 0.24257f
C258 drain_left.t18 a_n2354_n2688# 0.24257f
C259 drain_left.n0 a_n2354_n2688# 2.12501f
C260 drain_left.t19 a_n2354_n2688# 0.24257f
C261 drain_left.t4 a_n2354_n2688# 0.24257f
C262 drain_left.n1 a_n2354_n2688# 2.12168f
C263 drain_left.n2 a_n2354_n2688# 0.795543f
C264 drain_left.t20 a_n2354_n2688# 0.24257f
C265 drain_left.t10 a_n2354_n2688# 0.24257f
C266 drain_left.n3 a_n2354_n2688# 2.12168f
C267 drain_left.n4 a_n2354_n2688# 0.360304f
C268 drain_left.t22 a_n2354_n2688# 0.24257f
C269 drain_left.t5 a_n2354_n2688# 0.24257f
C270 drain_left.n5 a_n2354_n2688# 2.12501f
C271 drain_left.t16 a_n2354_n2688# 0.24257f
C272 drain_left.t3 a_n2354_n2688# 0.24257f
C273 drain_left.n6 a_n2354_n2688# 2.12168f
C274 drain_left.n7 a_n2354_n2688# 0.795543f
C275 drain_left.t14 a_n2354_n2688# 0.24257f
C276 drain_left.t23 a_n2354_n2688# 0.24257f
C277 drain_left.n8 a_n2354_n2688# 2.12168f
C278 drain_left.n9 a_n2354_n2688# 0.360304f
C279 drain_left.n10 a_n2354_n2688# 1.61895f
C280 drain_left.t9 a_n2354_n2688# 0.24257f
C281 drain_left.t6 a_n2354_n2688# 0.24257f
C282 drain_left.n11 a_n2354_n2688# 2.12502f
C283 drain_left.t0 a_n2354_n2688# 0.24257f
C284 drain_left.t11 a_n2354_n2688# 0.24257f
C285 drain_left.n12 a_n2354_n2688# 2.12168f
C286 drain_left.n13 a_n2354_n2688# 0.795535f
C287 drain_left.t8 a_n2354_n2688# 0.24257f
C288 drain_left.t13 a_n2354_n2688# 0.24257f
C289 drain_left.n14 a_n2354_n2688# 2.12168f
C290 drain_left.n15 a_n2354_n2688# 0.392568f
C291 drain_left.t12 a_n2354_n2688# 0.24257f
C292 drain_left.t7 a_n2354_n2688# 0.24257f
C293 drain_left.n16 a_n2354_n2688# 2.12168f
C294 drain_left.n17 a_n2354_n2688# 0.392568f
C295 drain_left.t21 a_n2354_n2688# 0.24257f
C296 drain_left.t2 a_n2354_n2688# 0.24257f
C297 drain_left.n18 a_n2354_n2688# 2.12168f
C298 drain_left.n19 a_n2354_n2688# 0.392568f
C299 drain_left.t15 a_n2354_n2688# 0.24257f
C300 drain_left.t17 a_n2354_n2688# 0.24257f
C301 drain_left.n20 a_n2354_n2688# 2.12167f
C302 drain_left.n21 a_n2354_n2688# 0.676469f
C303 plus.n0 a_n2354_n2688# 0.049009f
C304 plus.t0 a_n2354_n2688# 0.374958f
C305 plus.t19 a_n2354_n2688# 0.374958f
C306 plus.n1 a_n2354_n2688# 0.156576f
C307 plus.n2 a_n2354_n2688# 0.049009f
C308 plus.t12 a_n2354_n2688# 0.374958f
C309 plus.t1 a_n2354_n2688# 0.374958f
C310 plus.t20 a_n2354_n2688# 0.374958f
C311 plus.n3 a_n2354_n2688# 0.156576f
C312 plus.n4 a_n2354_n2688# 0.049009f
C313 plus.t15 a_n2354_n2688# 0.374958f
C314 plus.t8 a_n2354_n2688# 0.374958f
C315 plus.n5 a_n2354_n2688# 0.156576f
C316 plus.n6 a_n2354_n2688# 0.049009f
C317 plus.t22 a_n2354_n2688# 0.374958f
C318 plus.t17 a_n2354_n2688# 0.374958f
C319 plus.n7 a_n2354_n2688# 0.018826f
C320 plus.t4 a_n2354_n2688# 0.3807f
C321 plus.t11 a_n2354_n2688# 0.374958f
C322 plus.n8 a_n2354_n2688# 0.156576f
C323 plus.n9 a_n2354_n2688# 0.171539f
C324 plus.n10 a_n2354_n2688# 0.104903f
C325 plus.n11 a_n2354_n2688# 0.049009f
C326 plus.n12 a_n2354_n2688# 0.017618f
C327 plus.n13 a_n2354_n2688# 0.156576f
C328 plus.n14 a_n2354_n2688# 0.020186f
C329 plus.n15 a_n2354_n2688# 0.156576f
C330 plus.n16 a_n2354_n2688# 0.020186f
C331 plus.n17 a_n2354_n2688# 0.049009f
C332 plus.n18 a_n2354_n2688# 0.049009f
C333 plus.n19 a_n2354_n2688# 0.020186f
C334 plus.n20 a_n2354_n2688# 0.156576f
C335 plus.n21 a_n2354_n2688# 0.018222f
C336 plus.n22 a_n2354_n2688# 0.018222f
C337 plus.n23 a_n2354_n2688# 0.049009f
C338 plus.n24 a_n2354_n2688# 0.049009f
C339 plus.n25 a_n2354_n2688# 0.020186f
C340 plus.n26 a_n2354_n2688# 0.156576f
C341 plus.n27 a_n2354_n2688# 0.020186f
C342 plus.n28 a_n2354_n2688# 0.156576f
C343 plus.n29 a_n2354_n2688# 0.020186f
C344 plus.n30 a_n2354_n2688# 0.049009f
C345 plus.n31 a_n2354_n2688# 0.049009f
C346 plus.n32 a_n2354_n2688# 0.017618f
C347 plus.n33 a_n2354_n2688# 0.018826f
C348 plus.n34 a_n2354_n2688# 0.156576f
C349 plus.t5 a_n2354_n2688# 0.3807f
C350 plus.n35 a_n2354_n2688# 0.171474f
C351 plus.n36 a_n2354_n2688# 0.477872f
C352 plus.n37 a_n2354_n2688# 0.049009f
C353 plus.t21 a_n2354_n2688# 0.3807f
C354 plus.t6 a_n2354_n2688# 0.374958f
C355 plus.t14 a_n2354_n2688# 0.374958f
C356 plus.n38 a_n2354_n2688# 0.156576f
C357 plus.n39 a_n2354_n2688# 0.049009f
C358 plus.t23 a_n2354_n2688# 0.374958f
C359 plus.t13 a_n2354_n2688# 0.374958f
C360 plus.t3 a_n2354_n2688# 0.374958f
C361 plus.n40 a_n2354_n2688# 0.156576f
C362 plus.n41 a_n2354_n2688# 0.049009f
C363 plus.t10 a_n2354_n2688# 0.374958f
C364 plus.t2 a_n2354_n2688# 0.374958f
C365 plus.n42 a_n2354_n2688# 0.156576f
C366 plus.n43 a_n2354_n2688# 0.049009f
C367 plus.t9 a_n2354_n2688# 0.374958f
C368 plus.t18 a_n2354_n2688# 0.374958f
C369 plus.n44 a_n2354_n2688# 0.018826f
C370 plus.t7 a_n2354_n2688# 0.374958f
C371 plus.n45 a_n2354_n2688# 0.156576f
C372 plus.t16 a_n2354_n2688# 0.3807f
C373 plus.n46 a_n2354_n2688# 0.171539f
C374 plus.n47 a_n2354_n2688# 0.104903f
C375 plus.n48 a_n2354_n2688# 0.049009f
C376 plus.n49 a_n2354_n2688# 0.017618f
C377 plus.n50 a_n2354_n2688# 0.156576f
C378 plus.n51 a_n2354_n2688# 0.020186f
C379 plus.n52 a_n2354_n2688# 0.156576f
C380 plus.n53 a_n2354_n2688# 0.020186f
C381 plus.n54 a_n2354_n2688# 0.049009f
C382 plus.n55 a_n2354_n2688# 0.049009f
C383 plus.n56 a_n2354_n2688# 0.020186f
C384 plus.n57 a_n2354_n2688# 0.156576f
C385 plus.n58 a_n2354_n2688# 0.018222f
C386 plus.n59 a_n2354_n2688# 0.018222f
C387 plus.n60 a_n2354_n2688# 0.049009f
C388 plus.n61 a_n2354_n2688# 0.049009f
C389 plus.n62 a_n2354_n2688# 0.020186f
C390 plus.n63 a_n2354_n2688# 0.156576f
C391 plus.n64 a_n2354_n2688# 0.020186f
C392 plus.n65 a_n2354_n2688# 0.156576f
C393 plus.n66 a_n2354_n2688# 0.020186f
C394 plus.n67 a_n2354_n2688# 0.049009f
C395 plus.n68 a_n2354_n2688# 0.049009f
C396 plus.n69 a_n2354_n2688# 0.017618f
C397 plus.n70 a_n2354_n2688# 0.018826f
C398 plus.n71 a_n2354_n2688# 0.156576f
C399 plus.n72 a_n2354_n2688# 0.171474f
C400 plus.n73 a_n2354_n2688# 1.48349f
.ends

