* NGSPICE file created from diffpair228.ext - technology: sky130A

.subckt diffpair228 minus drain_right drain_left source plus
X0 drain_right.t19 minus.t0 source.t17 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X1 source.t13 minus.t1 drain_right.t18 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X2 source.t28 plus.t0 drain_left.t19 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X3 source.t31 plus.t1 drain_left.t18 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X4 source.t16 minus.t2 drain_right.t17 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X5 a_n2982_n1488# a_n2982_n1488# a_n2982_n1488# a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.7
X6 a_n2982_n1488# a_n2982_n1488# a_n2982_n1488# a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X7 drain_left.t17 plus.t2 source.t2 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X8 source.t0 plus.t3 drain_left.t16 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X9 source.t1 plus.t4 drain_left.t15 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X10 source.t3 plus.t5 drain_left.t14 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X11 drain_right.t16 minus.t3 source.t14 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X12 source.t15 minus.t4 drain_right.t15 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X13 drain_right.t14 minus.t5 source.t20 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X14 source.t19 minus.t6 drain_right.t13 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X15 drain_right.t12 minus.t7 source.t8 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X16 drain_left.t13 plus.t6 source.t29 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X17 source.t6 plus.t7 drain_left.t12 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X18 drain_left.t11 plus.t8 source.t36 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X19 source.t37 plus.t9 drain_left.t10 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X20 drain_right.t11 minus.t8 source.t9 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X21 drain_right.t10 minus.t9 source.t26 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X22 source.t7 minus.t10 drain_right.t9 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X23 drain_left.t9 plus.t10 source.t5 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X24 drain_right.t8 minus.t11 source.t21 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X25 drain_left.t8 plus.t11 source.t32 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X26 drain_right.t7 minus.t12 source.t10 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X27 drain_left.t7 plus.t12 source.t34 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X28 drain_left.t6 plus.t13 source.t27 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X29 drain_right.t6 minus.t13 source.t24 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X30 drain_left.t5 plus.t14 source.t30 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X31 a_n2982_n1488# a_n2982_n1488# a_n2982_n1488# a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X32 source.t22 minus.t14 drain_right.t5 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X33 a_n2982_n1488# a_n2982_n1488# a_n2982_n1488# a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X34 drain_right.t4 minus.t15 source.t11 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X35 drain_left.t4 plus.t15 source.t4 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X36 source.t23 minus.t16 drain_right.t3 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X37 source.t35 plus.t16 drain_left.t3 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X38 source.t18 minus.t17 drain_right.t2 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X39 drain_left.t2 plus.t17 source.t38 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X40 source.t12 minus.t18 drain_right.t1 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X41 source.t25 minus.t19 drain_right.t0 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X42 source.t33 plus.t18 drain_left.t1 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X43 source.t39 plus.t19 drain_left.t0 a_n2982_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
R0 minus.n9 minus.t13 184.798
R1 minus.n43 minus.t1 184.798
R2 minus.n33 minus.n32 161.3
R3 minus.n31 minus.n0 161.3
R4 minus.n30 minus.n29 161.3
R5 minus.n28 minus.n1 161.3
R6 minus.n27 minus.n26 161.3
R7 minus.n25 minus.n2 161.3
R8 minus.n24 minus.n23 161.3
R9 minus.n22 minus.n3 161.3
R10 minus.n21 minus.n20 161.3
R11 minus.n19 minus.n4 161.3
R12 minus.n18 minus.n17 161.3
R13 minus.n16 minus.n5 161.3
R14 minus.n15 minus.n14 161.3
R15 minus.n13 minus.n6 161.3
R16 minus.n12 minus.n11 161.3
R17 minus.n10 minus.n7 161.3
R18 minus.n67 minus.n66 161.3
R19 minus.n65 minus.n34 161.3
R20 minus.n64 minus.n63 161.3
R21 minus.n62 minus.n35 161.3
R22 minus.n61 minus.n60 161.3
R23 minus.n59 minus.n36 161.3
R24 minus.n58 minus.n57 161.3
R25 minus.n56 minus.n37 161.3
R26 minus.n55 minus.n54 161.3
R27 minus.n53 minus.n38 161.3
R28 minus.n52 minus.n51 161.3
R29 minus.n50 minus.n39 161.3
R30 minus.n49 minus.n48 161.3
R31 minus.n47 minus.n40 161.3
R32 minus.n46 minus.n45 161.3
R33 minus.n44 minus.n41 161.3
R34 minus.n8 minus.t2 159.405
R35 minus.n12 minus.t12 159.405
R36 minus.n14 minus.t18 159.405
R37 minus.n18 minus.t9 159.405
R38 minus.n20 minus.t19 159.405
R39 minus.n24 minus.t8 159.405
R40 minus.n26 minus.t17 159.405
R41 minus.n30 minus.t7 159.405
R42 minus.n32 minus.t16 159.405
R43 minus.n42 minus.t0 159.405
R44 minus.n46 minus.t4 159.405
R45 minus.n48 minus.t3 159.405
R46 minus.n52 minus.t6 159.405
R47 minus.n54 minus.t11 159.405
R48 minus.n58 minus.t10 159.405
R49 minus.n60 minus.t15 159.405
R50 minus.n64 minus.t14 159.405
R51 minus.n66 minus.t5 159.405
R52 minus.n10 minus.n9 45.0031
R53 minus.n44 minus.n43 45.0031
R54 minus.n32 minus.n31 41.6278
R55 minus.n66 minus.n65 41.6278
R56 minus.n8 minus.n7 37.246
R57 minus.n30 minus.n1 37.246
R58 minus.n42 minus.n41 37.246
R59 minus.n64 minus.n35 37.246
R60 minus.n68 minus.n33 33.7656
R61 minus.n13 minus.n12 32.8641
R62 minus.n26 minus.n25 32.8641
R63 minus.n47 minus.n46 32.8641
R64 minus.n60 minus.n59 32.8641
R65 minus.n14 minus.n5 28.4823
R66 minus.n24 minus.n3 28.4823
R67 minus.n48 minus.n39 28.4823
R68 minus.n58 minus.n37 28.4823
R69 minus.n20 minus.n19 24.1005
R70 minus.n19 minus.n18 24.1005
R71 minus.n53 minus.n52 24.1005
R72 minus.n54 minus.n53 24.1005
R73 minus.n18 minus.n5 19.7187
R74 minus.n20 minus.n3 19.7187
R75 minus.n52 minus.n39 19.7187
R76 minus.n54 minus.n37 19.7187
R77 minus.n9 minus.n8 15.6319
R78 minus.n43 minus.n42 15.6319
R79 minus.n14 minus.n13 15.3369
R80 minus.n25 minus.n24 15.3369
R81 minus.n48 minus.n47 15.3369
R82 minus.n59 minus.n58 15.3369
R83 minus.n12 minus.n7 10.955
R84 minus.n26 minus.n1 10.955
R85 minus.n46 minus.n41 10.955
R86 minus.n60 minus.n35 10.955
R87 minus.n68 minus.n67 6.66717
R88 minus.n31 minus.n30 6.57323
R89 minus.n65 minus.n64 6.57323
R90 minus.n33 minus.n0 0.189894
R91 minus.n29 minus.n0 0.189894
R92 minus.n29 minus.n28 0.189894
R93 minus.n28 minus.n27 0.189894
R94 minus.n27 minus.n2 0.189894
R95 minus.n23 minus.n2 0.189894
R96 minus.n23 minus.n22 0.189894
R97 minus.n22 minus.n21 0.189894
R98 minus.n21 minus.n4 0.189894
R99 minus.n17 minus.n4 0.189894
R100 minus.n17 minus.n16 0.189894
R101 minus.n16 minus.n15 0.189894
R102 minus.n15 minus.n6 0.189894
R103 minus.n11 minus.n6 0.189894
R104 minus.n11 minus.n10 0.189894
R105 minus.n45 minus.n44 0.189894
R106 minus.n45 minus.n40 0.189894
R107 minus.n49 minus.n40 0.189894
R108 minus.n50 minus.n49 0.189894
R109 minus.n51 minus.n50 0.189894
R110 minus.n51 minus.n38 0.189894
R111 minus.n55 minus.n38 0.189894
R112 minus.n56 minus.n55 0.189894
R113 minus.n57 minus.n56 0.189894
R114 minus.n57 minus.n36 0.189894
R115 minus.n61 minus.n36 0.189894
R116 minus.n62 minus.n61 0.189894
R117 minus.n63 minus.n62 0.189894
R118 minus.n63 minus.n34 0.189894
R119 minus.n67 minus.n34 0.189894
R120 minus minus.n68 0.188
R121 source.n0 source.t2 69.6943
R122 source.n9 source.t3 69.6943
R123 source.n10 source.t24 69.6943
R124 source.n19 source.t23 69.6943
R125 source.n39 source.t20 69.6942
R126 source.n30 source.t13 69.6942
R127 source.n29 source.t29 69.6942
R128 source.n20 source.t37 69.6942
R129 source.n2 source.n1 63.0943
R130 source.n4 source.n3 63.0943
R131 source.n6 source.n5 63.0943
R132 source.n8 source.n7 63.0943
R133 source.n12 source.n11 63.0943
R134 source.n14 source.n13 63.0943
R135 source.n16 source.n15 63.0943
R136 source.n18 source.n17 63.0943
R137 source.n38 source.n37 63.0942
R138 source.n36 source.n35 63.0942
R139 source.n34 source.n33 63.0942
R140 source.n32 source.n31 63.0942
R141 source.n28 source.n27 63.0942
R142 source.n26 source.n25 63.0942
R143 source.n24 source.n23 63.0942
R144 source.n22 source.n21 63.0942
R145 source.n20 source.n19 15.3575
R146 source.n40 source.n0 9.65058
R147 source.n37 source.t11 6.6005
R148 source.n37 source.t22 6.6005
R149 source.n35 source.t21 6.6005
R150 source.n35 source.t7 6.6005
R151 source.n33 source.t14 6.6005
R152 source.n33 source.t19 6.6005
R153 source.n31 source.t17 6.6005
R154 source.n31 source.t15 6.6005
R155 source.n27 source.t32 6.6005
R156 source.n27 source.t6 6.6005
R157 source.n25 source.t4 6.6005
R158 source.n25 source.t35 6.6005
R159 source.n23 source.t38 6.6005
R160 source.n23 source.t33 6.6005
R161 source.n21 source.t36 6.6005
R162 source.n21 source.t0 6.6005
R163 source.n1 source.t5 6.6005
R164 source.n1 source.t39 6.6005
R165 source.n3 source.t27 6.6005
R166 source.n3 source.t28 6.6005
R167 source.n5 source.t34 6.6005
R168 source.n5 source.t1 6.6005
R169 source.n7 source.t30 6.6005
R170 source.n7 source.t31 6.6005
R171 source.n11 source.t10 6.6005
R172 source.n11 source.t16 6.6005
R173 source.n13 source.t26 6.6005
R174 source.n13 source.t12 6.6005
R175 source.n15 source.t9 6.6005
R176 source.n15 source.t25 6.6005
R177 source.n17 source.t8 6.6005
R178 source.n17 source.t18 6.6005
R179 source.n40 source.n39 5.7074
R180 source.n19 source.n18 0.888431
R181 source.n18 source.n16 0.888431
R182 source.n16 source.n14 0.888431
R183 source.n14 source.n12 0.888431
R184 source.n12 source.n10 0.888431
R185 source.n9 source.n8 0.888431
R186 source.n8 source.n6 0.888431
R187 source.n6 source.n4 0.888431
R188 source.n4 source.n2 0.888431
R189 source.n2 source.n0 0.888431
R190 source.n22 source.n20 0.888431
R191 source.n24 source.n22 0.888431
R192 source.n26 source.n24 0.888431
R193 source.n28 source.n26 0.888431
R194 source.n29 source.n28 0.888431
R195 source.n32 source.n30 0.888431
R196 source.n34 source.n32 0.888431
R197 source.n36 source.n34 0.888431
R198 source.n38 source.n36 0.888431
R199 source.n39 source.n38 0.888431
R200 source.n10 source.n9 0.470328
R201 source.n30 source.n29 0.470328
R202 source source.n40 0.188
R203 drain_right.n10 drain_right.n8 80.661
R204 drain_right.n6 drain_right.n4 80.6609
R205 drain_right.n2 drain_right.n0 80.6609
R206 drain_right.n10 drain_right.n9 79.7731
R207 drain_right.n12 drain_right.n11 79.7731
R208 drain_right.n14 drain_right.n13 79.7731
R209 drain_right.n16 drain_right.n15 79.7731
R210 drain_right.n7 drain_right.n3 79.773
R211 drain_right.n6 drain_right.n5 79.773
R212 drain_right.n2 drain_right.n1 79.773
R213 drain_right drain_right.n7 27.0991
R214 drain_right.n3 drain_right.t13 6.6005
R215 drain_right.n3 drain_right.t8 6.6005
R216 drain_right.n4 drain_right.t5 6.6005
R217 drain_right.n4 drain_right.t14 6.6005
R218 drain_right.n5 drain_right.t9 6.6005
R219 drain_right.n5 drain_right.t4 6.6005
R220 drain_right.n1 drain_right.t15 6.6005
R221 drain_right.n1 drain_right.t16 6.6005
R222 drain_right.n0 drain_right.t18 6.6005
R223 drain_right.n0 drain_right.t19 6.6005
R224 drain_right.n8 drain_right.t17 6.6005
R225 drain_right.n8 drain_right.t6 6.6005
R226 drain_right.n9 drain_right.t1 6.6005
R227 drain_right.n9 drain_right.t7 6.6005
R228 drain_right.n11 drain_right.t0 6.6005
R229 drain_right.n11 drain_right.t10 6.6005
R230 drain_right.n13 drain_right.t2 6.6005
R231 drain_right.n13 drain_right.t11 6.6005
R232 drain_right.n15 drain_right.t3 6.6005
R233 drain_right.n15 drain_right.t12 6.6005
R234 drain_right drain_right.n16 6.54115
R235 drain_right.n16 drain_right.n14 0.888431
R236 drain_right.n14 drain_right.n12 0.888431
R237 drain_right.n12 drain_right.n10 0.888431
R238 drain_right.n7 drain_right.n6 0.833085
R239 drain_right.n7 drain_right.n2 0.833085
R240 plus.n9 plus.t5 184.798
R241 plus.n43 plus.t6 184.798
R242 plus.n11 plus.n10 161.3
R243 plus.n12 plus.n7 161.3
R244 plus.n14 plus.n13 161.3
R245 plus.n15 plus.n6 161.3
R246 plus.n17 plus.n16 161.3
R247 plus.n18 plus.n5 161.3
R248 plus.n20 plus.n19 161.3
R249 plus.n21 plus.n4 161.3
R250 plus.n23 plus.n22 161.3
R251 plus.n24 plus.n3 161.3
R252 plus.n26 plus.n25 161.3
R253 plus.n27 plus.n2 161.3
R254 plus.n29 plus.n28 161.3
R255 plus.n30 plus.n1 161.3
R256 plus.n31 plus.n0 161.3
R257 plus.n33 plus.n32 161.3
R258 plus.n45 plus.n44 161.3
R259 plus.n46 plus.n41 161.3
R260 plus.n48 plus.n47 161.3
R261 plus.n49 plus.n40 161.3
R262 plus.n51 plus.n50 161.3
R263 plus.n52 plus.n39 161.3
R264 plus.n54 plus.n53 161.3
R265 plus.n55 plus.n38 161.3
R266 plus.n57 plus.n56 161.3
R267 plus.n58 plus.n37 161.3
R268 plus.n60 plus.n59 161.3
R269 plus.n61 plus.n36 161.3
R270 plus.n63 plus.n62 161.3
R271 plus.n64 plus.n35 161.3
R272 plus.n65 plus.n34 161.3
R273 plus.n67 plus.n66 161.3
R274 plus.n32 plus.t2 159.405
R275 plus.n30 plus.t19 159.405
R276 plus.n2 plus.t10 159.405
R277 plus.n24 plus.t0 159.405
R278 plus.n4 plus.t13 159.405
R279 plus.n18 plus.t4 159.405
R280 plus.n6 plus.t12 159.405
R281 plus.n12 plus.t1 159.405
R282 plus.n8 plus.t14 159.405
R283 plus.n66 plus.t9 159.405
R284 plus.n64 plus.t8 159.405
R285 plus.n36 plus.t3 159.405
R286 plus.n58 plus.t17 159.405
R287 plus.n38 plus.t18 159.405
R288 plus.n52 plus.t15 159.405
R289 plus.n40 plus.t16 159.405
R290 plus.n46 plus.t11 159.405
R291 plus.n42 plus.t7 159.405
R292 plus.n10 plus.n9 45.0031
R293 plus.n44 plus.n43 45.0031
R294 plus.n32 plus.n31 41.6278
R295 plus.n66 plus.n65 41.6278
R296 plus.n30 plus.n29 37.246
R297 plus.n11 plus.n8 37.246
R298 plus.n64 plus.n63 37.246
R299 plus.n45 plus.n42 37.246
R300 plus.n25 plus.n2 32.8641
R301 plus.n13 plus.n12 32.8641
R302 plus.n59 plus.n36 32.8641
R303 plus.n47 plus.n46 32.8641
R304 plus plus.n67 31.0558
R305 plus.n24 plus.n23 28.4823
R306 plus.n17 plus.n6 28.4823
R307 plus.n58 plus.n57 28.4823
R308 plus.n51 plus.n40 28.4823
R309 plus.n19 plus.n18 24.1005
R310 plus.n19 plus.n4 24.1005
R311 plus.n53 plus.n38 24.1005
R312 plus.n53 plus.n52 24.1005
R313 plus.n23 plus.n4 19.7187
R314 plus.n18 plus.n17 19.7187
R315 plus.n57 plus.n38 19.7187
R316 plus.n52 plus.n51 19.7187
R317 plus.n9 plus.n8 15.6319
R318 plus.n43 plus.n42 15.6319
R319 plus.n25 plus.n24 15.3369
R320 plus.n13 plus.n6 15.3369
R321 plus.n59 plus.n58 15.3369
R322 plus.n47 plus.n40 15.3369
R323 plus.n29 plus.n2 10.955
R324 plus.n12 plus.n11 10.955
R325 plus.n63 plus.n36 10.955
R326 plus.n46 plus.n45 10.955
R327 plus plus.n33 8.90202
R328 plus.n31 plus.n30 6.57323
R329 plus.n65 plus.n64 6.57323
R330 plus.n10 plus.n7 0.189894
R331 plus.n14 plus.n7 0.189894
R332 plus.n15 plus.n14 0.189894
R333 plus.n16 plus.n15 0.189894
R334 plus.n16 plus.n5 0.189894
R335 plus.n20 plus.n5 0.189894
R336 plus.n21 plus.n20 0.189894
R337 plus.n22 plus.n21 0.189894
R338 plus.n22 plus.n3 0.189894
R339 plus.n26 plus.n3 0.189894
R340 plus.n27 plus.n26 0.189894
R341 plus.n28 plus.n27 0.189894
R342 plus.n28 plus.n1 0.189894
R343 plus.n1 plus.n0 0.189894
R344 plus.n33 plus.n0 0.189894
R345 plus.n67 plus.n34 0.189894
R346 plus.n35 plus.n34 0.189894
R347 plus.n62 plus.n35 0.189894
R348 plus.n62 plus.n61 0.189894
R349 plus.n61 plus.n60 0.189894
R350 plus.n60 plus.n37 0.189894
R351 plus.n56 plus.n37 0.189894
R352 plus.n56 plus.n55 0.189894
R353 plus.n55 plus.n54 0.189894
R354 plus.n54 plus.n39 0.189894
R355 plus.n50 plus.n39 0.189894
R356 plus.n50 plus.n49 0.189894
R357 plus.n49 plus.n48 0.189894
R358 plus.n48 plus.n41 0.189894
R359 plus.n44 plus.n41 0.189894
R360 drain_left.n10 drain_left.n8 80.661
R361 drain_left.n6 drain_left.n4 80.6609
R362 drain_left.n2 drain_left.n0 80.6609
R363 drain_left.n16 drain_left.n15 79.7731
R364 drain_left.n14 drain_left.n13 79.7731
R365 drain_left.n12 drain_left.n11 79.7731
R366 drain_left.n10 drain_left.n9 79.7731
R367 drain_left.n7 drain_left.n3 79.773
R368 drain_left.n6 drain_left.n5 79.773
R369 drain_left.n2 drain_left.n1 79.773
R370 drain_left drain_left.n7 27.6523
R371 drain_left.n3 drain_left.t1 6.6005
R372 drain_left.n3 drain_left.t4 6.6005
R373 drain_left.n4 drain_left.t12 6.6005
R374 drain_left.n4 drain_left.t13 6.6005
R375 drain_left.n5 drain_left.t3 6.6005
R376 drain_left.n5 drain_left.t8 6.6005
R377 drain_left.n1 drain_left.t16 6.6005
R378 drain_left.n1 drain_left.t2 6.6005
R379 drain_left.n0 drain_left.t10 6.6005
R380 drain_left.n0 drain_left.t11 6.6005
R381 drain_left.n15 drain_left.t0 6.6005
R382 drain_left.n15 drain_left.t17 6.6005
R383 drain_left.n13 drain_left.t19 6.6005
R384 drain_left.n13 drain_left.t9 6.6005
R385 drain_left.n11 drain_left.t15 6.6005
R386 drain_left.n11 drain_left.t6 6.6005
R387 drain_left.n9 drain_left.t18 6.6005
R388 drain_left.n9 drain_left.t7 6.6005
R389 drain_left.n8 drain_left.t14 6.6005
R390 drain_left.n8 drain_left.t5 6.6005
R391 drain_left drain_left.n16 6.54115
R392 drain_left.n12 drain_left.n10 0.888431
R393 drain_left.n14 drain_left.n12 0.888431
R394 drain_left.n16 drain_left.n14 0.888431
R395 drain_left.n7 drain_left.n6 0.833085
R396 drain_left.n7 drain_left.n2 0.833085
C0 drain_right source 9.09751f
C1 plus minus 5.20567f
C2 drain_right drain_left 1.59887f
C3 drain_left source 9.09514f
C4 drain_right minus 3.6682f
C5 drain_right plus 0.46039f
C6 source minus 4.32983f
C7 source plus 4.34383f
C8 drain_left minus 0.178628f
C9 drain_left plus 3.96566f
C10 drain_right a_n2982_n1488# 5.60505f
C11 drain_left a_n2982_n1488# 6.03955f
C12 source a_n2982_n1488# 4.097922f
C13 minus a_n2982_n1488# 11.232555f
C14 plus a_n2982_n1488# 12.64236f
C15 drain_left.t10 a_n2982_n1488# 0.064947f
C16 drain_left.t11 a_n2982_n1488# 0.064947f
C17 drain_left.n0 a_n2982_n1488# 0.472649f
C18 drain_left.t16 a_n2982_n1488# 0.064947f
C19 drain_left.t2 a_n2982_n1488# 0.064947f
C20 drain_left.n1 a_n2982_n1488# 0.468388f
C21 drain_left.n2 a_n2982_n1488# 0.754774f
C22 drain_left.t1 a_n2982_n1488# 0.064947f
C23 drain_left.t4 a_n2982_n1488# 0.064947f
C24 drain_left.n3 a_n2982_n1488# 0.468388f
C25 drain_left.t12 a_n2982_n1488# 0.064947f
C26 drain_left.t13 a_n2982_n1488# 0.064947f
C27 drain_left.n4 a_n2982_n1488# 0.472649f
C28 drain_left.t3 a_n2982_n1488# 0.064947f
C29 drain_left.t8 a_n2982_n1488# 0.064947f
C30 drain_left.n5 a_n2982_n1488# 0.468388f
C31 drain_left.n6 a_n2982_n1488# 0.754774f
C32 drain_left.n7 a_n2982_n1488# 1.46552f
C33 drain_left.t14 a_n2982_n1488# 0.064947f
C34 drain_left.t5 a_n2982_n1488# 0.064947f
C35 drain_left.n8 a_n2982_n1488# 0.472652f
C36 drain_left.t18 a_n2982_n1488# 0.064947f
C37 drain_left.t7 a_n2982_n1488# 0.064947f
C38 drain_left.n9 a_n2982_n1488# 0.46839f
C39 drain_left.n10 a_n2982_n1488# 0.758892f
C40 drain_left.t15 a_n2982_n1488# 0.064947f
C41 drain_left.t6 a_n2982_n1488# 0.064947f
C42 drain_left.n11 a_n2982_n1488# 0.46839f
C43 drain_left.n12 a_n2982_n1488# 0.37606f
C44 drain_left.t19 a_n2982_n1488# 0.064947f
C45 drain_left.t9 a_n2982_n1488# 0.064947f
C46 drain_left.n13 a_n2982_n1488# 0.46839f
C47 drain_left.n14 a_n2982_n1488# 0.37606f
C48 drain_left.t0 a_n2982_n1488# 0.064947f
C49 drain_left.t17 a_n2982_n1488# 0.064947f
C50 drain_left.n15 a_n2982_n1488# 0.46839f
C51 drain_left.n16 a_n2982_n1488# 0.618375f
C52 plus.n0 a_n2982_n1488# 0.042721f
C53 plus.t2 a_n2982_n1488# 0.26902f
C54 plus.t19 a_n2982_n1488# 0.26902f
C55 plus.n1 a_n2982_n1488# 0.042721f
C56 plus.t10 a_n2982_n1488# 0.26902f
C57 plus.n2 a_n2982_n1488# 0.156683f
C58 plus.n3 a_n2982_n1488# 0.042721f
C59 plus.t0 a_n2982_n1488# 0.26902f
C60 plus.t13 a_n2982_n1488# 0.26902f
C61 plus.n4 a_n2982_n1488# 0.156683f
C62 plus.n5 a_n2982_n1488# 0.042721f
C63 plus.t4 a_n2982_n1488# 0.26902f
C64 plus.t12 a_n2982_n1488# 0.26902f
C65 plus.n6 a_n2982_n1488# 0.156683f
C66 plus.n7 a_n2982_n1488# 0.042721f
C67 plus.t1 a_n2982_n1488# 0.26902f
C68 plus.t14 a_n2982_n1488# 0.26902f
C69 plus.n8 a_n2982_n1488# 0.163829f
C70 plus.t5 a_n2982_n1488# 0.29061f
C71 plus.n9 a_n2982_n1488# 0.13816f
C72 plus.n10 a_n2982_n1488# 0.18235f
C73 plus.n11 a_n2982_n1488# 0.009694f
C74 plus.n12 a_n2982_n1488# 0.156683f
C75 plus.n13 a_n2982_n1488# 0.009694f
C76 plus.n14 a_n2982_n1488# 0.042721f
C77 plus.n15 a_n2982_n1488# 0.042721f
C78 plus.n16 a_n2982_n1488# 0.042721f
C79 plus.n17 a_n2982_n1488# 0.009694f
C80 plus.n18 a_n2982_n1488# 0.156683f
C81 plus.n19 a_n2982_n1488# 0.009694f
C82 plus.n20 a_n2982_n1488# 0.042721f
C83 plus.n21 a_n2982_n1488# 0.042721f
C84 plus.n22 a_n2982_n1488# 0.042721f
C85 plus.n23 a_n2982_n1488# 0.009694f
C86 plus.n24 a_n2982_n1488# 0.156683f
C87 plus.n25 a_n2982_n1488# 0.009694f
C88 plus.n26 a_n2982_n1488# 0.042721f
C89 plus.n27 a_n2982_n1488# 0.042721f
C90 plus.n28 a_n2982_n1488# 0.042721f
C91 plus.n29 a_n2982_n1488# 0.009694f
C92 plus.n30 a_n2982_n1488# 0.156683f
C93 plus.n31 a_n2982_n1488# 0.009694f
C94 plus.n32 a_n2982_n1488# 0.156288f
C95 plus.n33 a_n2982_n1488# 0.336712f
C96 plus.n34 a_n2982_n1488# 0.042721f
C97 plus.t9 a_n2982_n1488# 0.26902f
C98 plus.n35 a_n2982_n1488# 0.042721f
C99 plus.t8 a_n2982_n1488# 0.26902f
C100 plus.t3 a_n2982_n1488# 0.26902f
C101 plus.n36 a_n2982_n1488# 0.156683f
C102 plus.n37 a_n2982_n1488# 0.042721f
C103 plus.t17 a_n2982_n1488# 0.26902f
C104 plus.t18 a_n2982_n1488# 0.26902f
C105 plus.n38 a_n2982_n1488# 0.156683f
C106 plus.n39 a_n2982_n1488# 0.042721f
C107 plus.t15 a_n2982_n1488# 0.26902f
C108 plus.t16 a_n2982_n1488# 0.26902f
C109 plus.n40 a_n2982_n1488# 0.156683f
C110 plus.n41 a_n2982_n1488# 0.042721f
C111 plus.t11 a_n2982_n1488# 0.26902f
C112 plus.t7 a_n2982_n1488# 0.26902f
C113 plus.n42 a_n2982_n1488# 0.163829f
C114 plus.t6 a_n2982_n1488# 0.29061f
C115 plus.n43 a_n2982_n1488# 0.13816f
C116 plus.n44 a_n2982_n1488# 0.18235f
C117 plus.n45 a_n2982_n1488# 0.009694f
C118 plus.n46 a_n2982_n1488# 0.156683f
C119 plus.n47 a_n2982_n1488# 0.009694f
C120 plus.n48 a_n2982_n1488# 0.042721f
C121 plus.n49 a_n2982_n1488# 0.042721f
C122 plus.n50 a_n2982_n1488# 0.042721f
C123 plus.n51 a_n2982_n1488# 0.009694f
C124 plus.n52 a_n2982_n1488# 0.156683f
C125 plus.n53 a_n2982_n1488# 0.009694f
C126 plus.n54 a_n2982_n1488# 0.042721f
C127 plus.n55 a_n2982_n1488# 0.042721f
C128 plus.n56 a_n2982_n1488# 0.042721f
C129 plus.n57 a_n2982_n1488# 0.009694f
C130 plus.n58 a_n2982_n1488# 0.156683f
C131 plus.n59 a_n2982_n1488# 0.009694f
C132 plus.n60 a_n2982_n1488# 0.042721f
C133 plus.n61 a_n2982_n1488# 0.042721f
C134 plus.n62 a_n2982_n1488# 0.042721f
C135 plus.n63 a_n2982_n1488# 0.009694f
C136 plus.n64 a_n2982_n1488# 0.156683f
C137 plus.n65 a_n2982_n1488# 0.009694f
C138 plus.n66 a_n2982_n1488# 0.156288f
C139 plus.n67 a_n2982_n1488# 1.27503f
C140 drain_right.t18 a_n2982_n1488# 0.063983f
C141 drain_right.t19 a_n2982_n1488# 0.063983f
C142 drain_right.n0 a_n2982_n1488# 0.465634f
C143 drain_right.t15 a_n2982_n1488# 0.063983f
C144 drain_right.t16 a_n2982_n1488# 0.063983f
C145 drain_right.n1 a_n2982_n1488# 0.461436f
C146 drain_right.n2 a_n2982_n1488# 0.743572f
C147 drain_right.t13 a_n2982_n1488# 0.063983f
C148 drain_right.t8 a_n2982_n1488# 0.063983f
C149 drain_right.n3 a_n2982_n1488# 0.461436f
C150 drain_right.t5 a_n2982_n1488# 0.063983f
C151 drain_right.t14 a_n2982_n1488# 0.063983f
C152 drain_right.n4 a_n2982_n1488# 0.465634f
C153 drain_right.t9 a_n2982_n1488# 0.063983f
C154 drain_right.t4 a_n2982_n1488# 0.063983f
C155 drain_right.n5 a_n2982_n1488# 0.461436f
C156 drain_right.n6 a_n2982_n1488# 0.743572f
C157 drain_right.n7 a_n2982_n1488# 1.39099f
C158 drain_right.t17 a_n2982_n1488# 0.063983f
C159 drain_right.t6 a_n2982_n1488# 0.063983f
C160 drain_right.n8 a_n2982_n1488# 0.465637f
C161 drain_right.t1 a_n2982_n1488# 0.063983f
C162 drain_right.t7 a_n2982_n1488# 0.063983f
C163 drain_right.n9 a_n2982_n1488# 0.461439f
C164 drain_right.n10 a_n2982_n1488# 0.747629f
C165 drain_right.t0 a_n2982_n1488# 0.063983f
C166 drain_right.t10 a_n2982_n1488# 0.063983f
C167 drain_right.n11 a_n2982_n1488# 0.461439f
C168 drain_right.n12 a_n2982_n1488# 0.370478f
C169 drain_right.t2 a_n2982_n1488# 0.063983f
C170 drain_right.t11 a_n2982_n1488# 0.063983f
C171 drain_right.n13 a_n2982_n1488# 0.461439f
C172 drain_right.n14 a_n2982_n1488# 0.370478f
C173 drain_right.t3 a_n2982_n1488# 0.063983f
C174 drain_right.t12 a_n2982_n1488# 0.063983f
C175 drain_right.n15 a_n2982_n1488# 0.461439f
C176 drain_right.n16 a_n2982_n1488# 0.609198f
C177 source.t2 a_n2982_n1488# 0.570486f
C178 source.n0 a_n2982_n1488# 0.834893f
C179 source.t5 a_n2982_n1488# 0.068702f
C180 source.t39 a_n2982_n1488# 0.068702f
C181 source.n1 a_n2982_n1488# 0.435607f
C182 source.n2 a_n2982_n1488# 0.418277f
C183 source.t27 a_n2982_n1488# 0.068702f
C184 source.t28 a_n2982_n1488# 0.068702f
C185 source.n3 a_n2982_n1488# 0.435607f
C186 source.n4 a_n2982_n1488# 0.418277f
C187 source.t34 a_n2982_n1488# 0.068702f
C188 source.t1 a_n2982_n1488# 0.068702f
C189 source.n5 a_n2982_n1488# 0.435607f
C190 source.n6 a_n2982_n1488# 0.418277f
C191 source.t30 a_n2982_n1488# 0.068702f
C192 source.t31 a_n2982_n1488# 0.068702f
C193 source.n7 a_n2982_n1488# 0.435607f
C194 source.n8 a_n2982_n1488# 0.418277f
C195 source.t3 a_n2982_n1488# 0.570486f
C196 source.n9 a_n2982_n1488# 0.431725f
C197 source.t24 a_n2982_n1488# 0.570486f
C198 source.n10 a_n2982_n1488# 0.431725f
C199 source.t10 a_n2982_n1488# 0.068702f
C200 source.t16 a_n2982_n1488# 0.068702f
C201 source.n11 a_n2982_n1488# 0.435607f
C202 source.n12 a_n2982_n1488# 0.418277f
C203 source.t26 a_n2982_n1488# 0.068702f
C204 source.t12 a_n2982_n1488# 0.068702f
C205 source.n13 a_n2982_n1488# 0.435607f
C206 source.n14 a_n2982_n1488# 0.418277f
C207 source.t9 a_n2982_n1488# 0.068702f
C208 source.t25 a_n2982_n1488# 0.068702f
C209 source.n15 a_n2982_n1488# 0.435607f
C210 source.n16 a_n2982_n1488# 0.418277f
C211 source.t8 a_n2982_n1488# 0.068702f
C212 source.t18 a_n2982_n1488# 0.068702f
C213 source.n17 a_n2982_n1488# 0.435607f
C214 source.n18 a_n2982_n1488# 0.418277f
C215 source.t23 a_n2982_n1488# 0.570486f
C216 source.n19 a_n2982_n1488# 1.14481f
C217 source.t37 a_n2982_n1488# 0.570483f
C218 source.n20 a_n2982_n1488# 1.14481f
C219 source.t36 a_n2982_n1488# 0.068702f
C220 source.t0 a_n2982_n1488# 0.068702f
C221 source.n21 a_n2982_n1488# 0.435604f
C222 source.n22 a_n2982_n1488# 0.41828f
C223 source.t38 a_n2982_n1488# 0.068702f
C224 source.t33 a_n2982_n1488# 0.068702f
C225 source.n23 a_n2982_n1488# 0.435604f
C226 source.n24 a_n2982_n1488# 0.41828f
C227 source.t4 a_n2982_n1488# 0.068702f
C228 source.t35 a_n2982_n1488# 0.068702f
C229 source.n25 a_n2982_n1488# 0.435604f
C230 source.n26 a_n2982_n1488# 0.41828f
C231 source.t32 a_n2982_n1488# 0.068702f
C232 source.t6 a_n2982_n1488# 0.068702f
C233 source.n27 a_n2982_n1488# 0.435604f
C234 source.n28 a_n2982_n1488# 0.41828f
C235 source.t29 a_n2982_n1488# 0.570483f
C236 source.n29 a_n2982_n1488# 0.431728f
C237 source.t13 a_n2982_n1488# 0.570483f
C238 source.n30 a_n2982_n1488# 0.431728f
C239 source.t17 a_n2982_n1488# 0.068702f
C240 source.t15 a_n2982_n1488# 0.068702f
C241 source.n31 a_n2982_n1488# 0.435604f
C242 source.n32 a_n2982_n1488# 0.41828f
C243 source.t14 a_n2982_n1488# 0.068702f
C244 source.t19 a_n2982_n1488# 0.068702f
C245 source.n33 a_n2982_n1488# 0.435604f
C246 source.n34 a_n2982_n1488# 0.41828f
C247 source.t21 a_n2982_n1488# 0.068702f
C248 source.t7 a_n2982_n1488# 0.068702f
C249 source.n35 a_n2982_n1488# 0.435604f
C250 source.n36 a_n2982_n1488# 0.41828f
C251 source.t11 a_n2982_n1488# 0.068702f
C252 source.t22 a_n2982_n1488# 0.068702f
C253 source.n37 a_n2982_n1488# 0.435604f
C254 source.n38 a_n2982_n1488# 0.41828f
C255 source.t20 a_n2982_n1488# 0.570483f
C256 source.n39 a_n2982_n1488# 0.620762f
C257 source.n40 a_n2982_n1488# 0.854571f
C258 minus.n0 a_n2982_n1488# 0.041506f
C259 minus.n1 a_n2982_n1488# 0.009419f
C260 minus.t7 a_n2982_n1488# 0.261369f
C261 minus.n2 a_n2982_n1488# 0.041506f
C262 minus.n3 a_n2982_n1488# 0.009419f
C263 minus.t8 a_n2982_n1488# 0.261369f
C264 minus.n4 a_n2982_n1488# 0.041506f
C265 minus.n5 a_n2982_n1488# 0.009419f
C266 minus.t9 a_n2982_n1488# 0.261369f
C267 minus.n6 a_n2982_n1488# 0.041506f
C268 minus.n7 a_n2982_n1488# 0.009419f
C269 minus.t12 a_n2982_n1488# 0.261369f
C270 minus.t13 a_n2982_n1488# 0.282345f
C271 minus.t2 a_n2982_n1488# 0.261369f
C272 minus.n8 a_n2982_n1488# 0.15917f
C273 minus.n9 a_n2982_n1488# 0.134231f
C274 minus.n10 a_n2982_n1488# 0.177164f
C275 minus.n11 a_n2982_n1488# 0.041506f
C276 minus.n12 a_n2982_n1488# 0.152227f
C277 minus.n13 a_n2982_n1488# 0.009419f
C278 minus.t18 a_n2982_n1488# 0.261369f
C279 minus.n14 a_n2982_n1488# 0.152227f
C280 minus.n15 a_n2982_n1488# 0.041506f
C281 minus.n16 a_n2982_n1488# 0.041506f
C282 minus.n17 a_n2982_n1488# 0.041506f
C283 minus.n18 a_n2982_n1488# 0.152227f
C284 minus.n19 a_n2982_n1488# 0.009419f
C285 minus.t19 a_n2982_n1488# 0.261369f
C286 minus.n20 a_n2982_n1488# 0.152227f
C287 minus.n21 a_n2982_n1488# 0.041506f
C288 minus.n22 a_n2982_n1488# 0.041506f
C289 minus.n23 a_n2982_n1488# 0.041506f
C290 minus.n24 a_n2982_n1488# 0.152227f
C291 minus.n25 a_n2982_n1488# 0.009419f
C292 minus.t17 a_n2982_n1488# 0.261369f
C293 minus.n26 a_n2982_n1488# 0.152227f
C294 minus.n27 a_n2982_n1488# 0.041506f
C295 minus.n28 a_n2982_n1488# 0.041506f
C296 minus.n29 a_n2982_n1488# 0.041506f
C297 minus.n30 a_n2982_n1488# 0.152227f
C298 minus.n31 a_n2982_n1488# 0.009419f
C299 minus.t16 a_n2982_n1488# 0.261369f
C300 minus.n32 a_n2982_n1488# 0.151844f
C301 minus.n33 a_n2982_n1488# 1.31947f
C302 minus.n34 a_n2982_n1488# 0.041506f
C303 minus.n35 a_n2982_n1488# 0.009419f
C304 minus.n36 a_n2982_n1488# 0.041506f
C305 minus.n37 a_n2982_n1488# 0.009419f
C306 minus.n38 a_n2982_n1488# 0.041506f
C307 minus.n39 a_n2982_n1488# 0.009419f
C308 minus.n40 a_n2982_n1488# 0.041506f
C309 minus.n41 a_n2982_n1488# 0.009419f
C310 minus.t1 a_n2982_n1488# 0.282345f
C311 minus.t0 a_n2982_n1488# 0.261369f
C312 minus.n42 a_n2982_n1488# 0.15917f
C313 minus.n43 a_n2982_n1488# 0.134231f
C314 minus.n44 a_n2982_n1488# 0.177164f
C315 minus.n45 a_n2982_n1488# 0.041506f
C316 minus.t4 a_n2982_n1488# 0.261369f
C317 minus.n46 a_n2982_n1488# 0.152227f
C318 minus.n47 a_n2982_n1488# 0.009419f
C319 minus.t3 a_n2982_n1488# 0.261369f
C320 minus.n48 a_n2982_n1488# 0.152227f
C321 minus.n49 a_n2982_n1488# 0.041506f
C322 minus.n50 a_n2982_n1488# 0.041506f
C323 minus.n51 a_n2982_n1488# 0.041506f
C324 minus.t6 a_n2982_n1488# 0.261369f
C325 minus.n52 a_n2982_n1488# 0.152227f
C326 minus.n53 a_n2982_n1488# 0.009419f
C327 minus.t11 a_n2982_n1488# 0.261369f
C328 minus.n54 a_n2982_n1488# 0.152227f
C329 minus.n55 a_n2982_n1488# 0.041506f
C330 minus.n56 a_n2982_n1488# 0.041506f
C331 minus.n57 a_n2982_n1488# 0.041506f
C332 minus.t10 a_n2982_n1488# 0.261369f
C333 minus.n58 a_n2982_n1488# 0.152227f
C334 minus.n59 a_n2982_n1488# 0.009419f
C335 minus.t15 a_n2982_n1488# 0.261369f
C336 minus.n60 a_n2982_n1488# 0.152227f
C337 minus.n61 a_n2982_n1488# 0.041506f
C338 minus.n62 a_n2982_n1488# 0.041506f
C339 minus.n63 a_n2982_n1488# 0.041506f
C340 minus.t14 a_n2982_n1488# 0.261369f
C341 minus.n64 a_n2982_n1488# 0.152227f
C342 minus.n65 a_n2982_n1488# 0.009419f
C343 minus.t5 a_n2982_n1488# 0.261369f
C344 minus.n66 a_n2982_n1488# 0.151844f
C345 minus.n67 a_n2982_n1488# 0.287575f
C346 minus.n68 a_n2982_n1488# 1.6075f
.ends

