* NGSPICE file created from diffpair396.ext - technology: sky130A

.subckt diffpair396 minus drain_right drain_left source plus
X0 a_n2524_n2688# a_n2524_n2688# a_n2524_n2688# a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.8
X1 source.t27 minus.t0 drain_right.t11 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X2 source.t26 minus.t1 drain_right.t12 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X3 source.t2 plus.t0 drain_left.t13 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X4 a_n2524_n2688# a_n2524_n2688# a_n2524_n2688# a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X5 source.t8 plus.t1 drain_left.t12 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X6 a_n2524_n2688# a_n2524_n2688# a_n2524_n2688# a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X7 source.t25 minus.t2 drain_right.t8 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X8 drain_left.t11 plus.t2 source.t12 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X9 drain_right.t7 minus.t3 source.t24 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X10 drain_left.t10 plus.t3 source.t13 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X11 drain_left.t9 plus.t4 source.t6 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X12 source.t23 minus.t4 drain_right.t13 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X13 drain_right.t2 minus.t5 source.t22 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X14 drain_right.t0 minus.t6 source.t21 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X15 drain_right.t9 minus.t7 source.t20 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X16 drain_right.t3 minus.t8 source.t19 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X17 source.t18 minus.t9 drain_right.t5 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X18 source.t17 minus.t10 drain_right.t1 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X19 drain_left.t8 plus.t5 source.t5 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X20 drain_right.t10 minus.t11 source.t16 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X21 drain_left.t7 plus.t6 source.t10 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X22 drain_right.t4 minus.t12 source.t15 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X23 source.t4 plus.t7 drain_left.t6 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X24 source.t7 plus.t8 drain_left.t5 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X25 drain_right.t6 minus.t13 source.t14 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X26 source.t1 plus.t9 drain_left.t4 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X27 drain_left.t3 plus.t10 source.t0 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X28 drain_left.t2 plus.t11 source.t11 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X29 source.t9 plus.t12 drain_left.t1 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X30 a_n2524_n2688# a_n2524_n2688# a_n2524_n2688# a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X31 drain_left.t0 plus.t13 source.t3 a_n2524_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
R0 minus.n5 minus.t8 344.075
R1 minus.n23 minus.t13 344.075
R2 minus.n4 minus.t4 320.229
R3 minus.n8 minus.t3 320.229
R4 minus.n9 minus.t10 320.229
R5 minus.n10 minus.t11 320.229
R6 minus.n14 minus.t9 320.229
R7 minus.n16 minus.t6 320.229
R8 minus.n22 minus.t2 320.229
R9 minus.n26 minus.t7 320.229
R10 minus.n27 minus.t1 320.229
R11 minus.n28 minus.t12 320.229
R12 minus.n32 minus.t0 320.229
R13 minus.n34 minus.t5 320.229
R14 minus.n17 minus.n16 161.3
R15 minus.n15 minus.n0 161.3
R16 minus.n14 minus.n13 161.3
R17 minus.n12 minus.n1 161.3
R18 minus.n6 minus.n3 161.3
R19 minus.n35 minus.n34 161.3
R20 minus.n33 minus.n18 161.3
R21 minus.n32 minus.n31 161.3
R22 minus.n30 minus.n19 161.3
R23 minus.n24 minus.n21 161.3
R24 minus.n11 minus.n10 80.6037
R25 minus.n9 minus.n2 80.6037
R26 minus.n8 minus.n7 80.6037
R27 minus.n29 minus.n28 80.6037
R28 minus.n27 minus.n20 80.6037
R29 minus.n26 minus.n25 80.6037
R30 minus.n9 minus.n8 48.2005
R31 minus.n10 minus.n9 48.2005
R32 minus.n27 minus.n26 48.2005
R33 minus.n28 minus.n27 48.2005
R34 minus.n6 minus.n5 44.9119
R35 minus.n24 minus.n23 44.9119
R36 minus.n36 minus.n17 36.635
R37 minus.n16 minus.n15 35.055
R38 minus.n34 minus.n33 35.055
R39 minus.n8 minus.n3 32.1338
R40 minus.n10 minus.n1 32.1338
R41 minus.n26 minus.n21 32.1338
R42 minus.n28 minus.n19 32.1338
R43 minus.n5 minus.n4 17.739
R44 minus.n23 minus.n22 17.739
R45 minus.n4 minus.n3 16.0672
R46 minus.n14 minus.n1 16.0672
R47 minus.n22 minus.n21 16.0672
R48 minus.n32 minus.n19 16.0672
R49 minus.n15 minus.n14 13.146
R50 minus.n33 minus.n32 13.146
R51 minus.n36 minus.n35 6.72588
R52 minus.n11 minus.n2 0.380177
R53 minus.n7 minus.n2 0.380177
R54 minus.n25 minus.n20 0.380177
R55 minus.n29 minus.n20 0.380177
R56 minus.n12 minus.n11 0.285035
R57 minus.n7 minus.n6 0.285035
R58 minus.n25 minus.n24 0.285035
R59 minus.n30 minus.n29 0.285035
R60 minus.n17 minus.n0 0.189894
R61 minus.n13 minus.n0 0.189894
R62 minus.n13 minus.n12 0.189894
R63 minus.n31 minus.n30 0.189894
R64 minus.n31 minus.n18 0.189894
R65 minus.n35 minus.n18 0.189894
R66 minus minus.n36 0.188
R67 drain_right.n1 drain_right.t6 68.7115
R68 drain_right.n11 drain_right.t0 67.7376
R69 drain_right.n8 drain_right.n6 66.5116
R70 drain_right.n4 drain_right.n2 66.5115
R71 drain_right.n8 drain_right.n7 65.5376
R72 drain_right.n10 drain_right.n9 65.5376
R73 drain_right.n4 drain_right.n3 65.5373
R74 drain_right.n1 drain_right.n0 65.5373
R75 drain_right drain_right.n5 30.1424
R76 drain_right drain_right.n11 6.14028
R77 drain_right.n2 drain_right.t11 2.2005
R78 drain_right.n2 drain_right.t2 2.2005
R79 drain_right.n3 drain_right.t12 2.2005
R80 drain_right.n3 drain_right.t4 2.2005
R81 drain_right.n0 drain_right.t8 2.2005
R82 drain_right.n0 drain_right.t9 2.2005
R83 drain_right.n6 drain_right.t13 2.2005
R84 drain_right.n6 drain_right.t3 2.2005
R85 drain_right.n7 drain_right.t1 2.2005
R86 drain_right.n7 drain_right.t7 2.2005
R87 drain_right.n9 drain_right.t5 2.2005
R88 drain_right.n9 drain_right.t10 2.2005
R89 drain_right.n11 drain_right.n10 0.974638
R90 drain_right.n10 drain_right.n8 0.974638
R91 drain_right.n5 drain_right.n1 0.675757
R92 drain_right.n5 drain_right.n4 0.188688
R93 source.n7 source.t19 51.0588
R94 source.n27 source.t22 51.0586
R95 source.n20 source.t5 51.0586
R96 source.n0 source.t10 51.0586
R97 source.n2 source.n1 48.8588
R98 source.n4 source.n3 48.8588
R99 source.n6 source.n5 48.8588
R100 source.n9 source.n8 48.8588
R101 source.n11 source.n10 48.8588
R102 source.n13 source.n12 48.8588
R103 source.n26 source.n25 48.8586
R104 source.n24 source.n23 48.8586
R105 source.n22 source.n21 48.8586
R106 source.n19 source.n18 48.8586
R107 source.n17 source.n16 48.8586
R108 source.n15 source.n14 48.8586
R109 source.n15 source.n13 20.9633
R110 source.n28 source.n0 14.2391
R111 source.n28 source.n27 5.7505
R112 source.n25 source.t15 2.2005
R113 source.n25 source.t27 2.2005
R114 source.n23 source.t20 2.2005
R115 source.n23 source.t26 2.2005
R116 source.n21 source.t14 2.2005
R117 source.n21 source.t25 2.2005
R118 source.n18 source.t6 2.2005
R119 source.n18 source.t8 2.2005
R120 source.n16 source.t13 2.2005
R121 source.n16 source.t2 2.2005
R122 source.n14 source.t12 2.2005
R123 source.n14 source.t1 2.2005
R124 source.n1 source.t11 2.2005
R125 source.n1 source.t4 2.2005
R126 source.n3 source.t0 2.2005
R127 source.n3 source.t7 2.2005
R128 source.n5 source.t3 2.2005
R129 source.n5 source.t9 2.2005
R130 source.n8 source.t24 2.2005
R131 source.n8 source.t23 2.2005
R132 source.n10 source.t16 2.2005
R133 source.n10 source.t17 2.2005
R134 source.n12 source.t21 2.2005
R135 source.n12 source.t18 2.2005
R136 source.n13 source.n11 0.974638
R137 source.n11 source.n9 0.974638
R138 source.n9 source.n7 0.974638
R139 source.n6 source.n4 0.974638
R140 source.n4 source.n2 0.974638
R141 source.n2 source.n0 0.974638
R142 source.n17 source.n15 0.974638
R143 source.n19 source.n17 0.974638
R144 source.n20 source.n19 0.974638
R145 source.n24 source.n22 0.974638
R146 source.n26 source.n24 0.974638
R147 source.n27 source.n26 0.974638
R148 source.n7 source.n6 0.957397
R149 source.n22 source.n20 0.957397
R150 source source.n28 0.188
R151 plus.n5 plus.t13 344.075
R152 plus.n23 plus.t5 344.075
R153 plus.n16 plus.t6 320.229
R154 plus.n14 plus.t7 320.229
R155 plus.n2 plus.t11 320.229
R156 plus.n9 plus.t8 320.229
R157 plus.n8 plus.t10 320.229
R158 plus.n4 plus.t12 320.229
R159 plus.n34 plus.t2 320.229
R160 plus.n32 plus.t9 320.229
R161 plus.n20 plus.t3 320.229
R162 plus.n27 plus.t0 320.229
R163 plus.n26 plus.t4 320.229
R164 plus.n22 plus.t1 320.229
R165 plus.n7 plus.n6 161.3
R166 plus.n13 plus.n12 161.3
R167 plus.n14 plus.n1 161.3
R168 plus.n15 plus.n0 161.3
R169 plus.n17 plus.n16 161.3
R170 plus.n25 plus.n24 161.3
R171 plus.n31 plus.n30 161.3
R172 plus.n32 plus.n19 161.3
R173 plus.n33 plus.n18 161.3
R174 plus.n35 plus.n34 161.3
R175 plus.n8 plus.n3 80.6037
R176 plus.n10 plus.n9 80.6037
R177 plus.n11 plus.n2 80.6037
R178 plus.n26 plus.n21 80.6037
R179 plus.n28 plus.n27 80.6037
R180 plus.n29 plus.n20 80.6037
R181 plus.n9 plus.n2 48.2005
R182 plus.n9 plus.n8 48.2005
R183 plus.n27 plus.n20 48.2005
R184 plus.n27 plus.n26 48.2005
R185 plus.n24 plus.n23 44.9119
R186 plus.n6 plus.n5 44.9119
R187 plus.n16 plus.n15 35.055
R188 plus.n34 plus.n33 35.055
R189 plus.n13 plus.n2 32.1338
R190 plus.n8 plus.n7 32.1338
R191 plus.n31 plus.n20 32.1338
R192 plus.n26 plus.n25 32.1338
R193 plus plus.n35 31.6524
R194 plus.n23 plus.n22 17.739
R195 plus.n5 plus.n4 17.739
R196 plus.n14 plus.n13 16.0672
R197 plus.n7 plus.n4 16.0672
R198 plus.n32 plus.n31 16.0672
R199 plus.n25 plus.n22 16.0672
R200 plus.n15 plus.n14 13.146
R201 plus.n33 plus.n32 13.146
R202 plus plus.n17 11.2335
R203 plus.n10 plus.n3 0.380177
R204 plus.n11 plus.n10 0.380177
R205 plus.n29 plus.n28 0.380177
R206 plus.n28 plus.n21 0.380177
R207 plus.n6 plus.n3 0.285035
R208 plus.n12 plus.n11 0.285035
R209 plus.n30 plus.n29 0.285035
R210 plus.n24 plus.n21 0.285035
R211 plus.n12 plus.n1 0.189894
R212 plus.n1 plus.n0 0.189894
R213 plus.n17 plus.n0 0.189894
R214 plus.n35 plus.n18 0.189894
R215 plus.n19 plus.n18 0.189894
R216 plus.n30 plus.n19 0.189894
R217 drain_left.n7 drain_left.t0 68.7117
R218 drain_left.n1 drain_left.t11 68.7115
R219 drain_left.n4 drain_left.n2 66.5115
R220 drain_left.n9 drain_left.n8 65.5376
R221 drain_left.n7 drain_left.n6 65.5376
R222 drain_left.n11 drain_left.n10 65.5374
R223 drain_left.n4 drain_left.n3 65.5373
R224 drain_left.n1 drain_left.n0 65.5373
R225 drain_left drain_left.n5 30.6956
R226 drain_left drain_left.n11 6.62735
R227 drain_left.n2 drain_left.t12 2.2005
R228 drain_left.n2 drain_left.t8 2.2005
R229 drain_left.n3 drain_left.t13 2.2005
R230 drain_left.n3 drain_left.t9 2.2005
R231 drain_left.n0 drain_left.t4 2.2005
R232 drain_left.n0 drain_left.t10 2.2005
R233 drain_left.n10 drain_left.t6 2.2005
R234 drain_left.n10 drain_left.t7 2.2005
R235 drain_left.n8 drain_left.t5 2.2005
R236 drain_left.n8 drain_left.t2 2.2005
R237 drain_left.n6 drain_left.t1 2.2005
R238 drain_left.n6 drain_left.t3 2.2005
R239 drain_left.n9 drain_left.n7 0.974638
R240 drain_left.n11 drain_left.n9 0.974638
R241 drain_left.n5 drain_left.n1 0.675757
R242 drain_left.n5 drain_left.n4 0.188688
C0 source minus 7.57496f
C1 drain_left minus 0.173289f
C2 source drain_left 14.003599f
C3 drain_right plus 0.407865f
C4 plus minus 5.73109f
C5 source plus 7.58935f
C6 drain_left plus 7.6755f
C7 drain_right minus 7.42735f
C8 source drain_right 14f
C9 drain_left drain_right 1.31613f
C10 drain_right a_n2524_n2688# 6.862401f
C11 drain_left a_n2524_n2688# 7.24347f
C12 source a_n2524_n2688# 5.706505f
C13 minus a_n2524_n2688# 9.83227f
C14 plus a_n2524_n2688# 11.373989f
C15 drain_left.t11 a_n2524_n2688# 1.95556f
C16 drain_left.t4 a_n2524_n2688# 0.175204f
C17 drain_left.t10 a_n2524_n2688# 0.175204f
C18 drain_left.n0 a_n2524_n2688# 1.53245f
C19 drain_left.n1 a_n2524_n2688# 0.668397f
C20 drain_left.t12 a_n2524_n2688# 0.175204f
C21 drain_left.t8 a_n2524_n2688# 0.175204f
C22 drain_left.n2 a_n2524_n2688# 1.53775f
C23 drain_left.t13 a_n2524_n2688# 0.175204f
C24 drain_left.t9 a_n2524_n2688# 0.175204f
C25 drain_left.n3 a_n2524_n2688# 1.53245f
C26 drain_left.n4 a_n2524_n2688# 0.649227f
C27 drain_left.n5 a_n2524_n2688# 1.23975f
C28 drain_left.t0 a_n2524_n2688# 1.95556f
C29 drain_left.t1 a_n2524_n2688# 0.175204f
C30 drain_left.t3 a_n2524_n2688# 0.175204f
C31 drain_left.n6 a_n2524_n2688# 1.53246f
C32 drain_left.n7 a_n2524_n2688# 0.69127f
C33 drain_left.t5 a_n2524_n2688# 0.175204f
C34 drain_left.t2 a_n2524_n2688# 0.175204f
C35 drain_left.n8 a_n2524_n2688# 1.53246f
C36 drain_left.n9 a_n2524_n2688# 0.351976f
C37 drain_left.t6 a_n2524_n2688# 0.175204f
C38 drain_left.t7 a_n2524_n2688# 0.175204f
C39 drain_left.n10 a_n2524_n2688# 1.53245f
C40 drain_left.n11 a_n2524_n2688# 0.572881f
C41 plus.n0 a_n2524_n2688# 0.039995f
C42 plus.t6 a_n2524_n2688# 0.825831f
C43 plus.t7 a_n2524_n2688# 0.825831f
C44 plus.n1 a_n2524_n2688# 0.039995f
C45 plus.t11 a_n2524_n2688# 0.825831f
C46 plus.n2 a_n2524_n2688# 0.352885f
C47 plus.n3 a_n2524_n2688# 0.066616f
C48 plus.t8 a_n2524_n2688# 0.825831f
C49 plus.t10 a_n2524_n2688# 0.825831f
C50 plus.t12 a_n2524_n2688# 0.825831f
C51 plus.n4 a_n2524_n2688# 0.34827f
C52 plus.t13 a_n2524_n2688# 0.849799f
C53 plus.n5 a_n2524_n2688# 0.325329f
C54 plus.n6 a_n2524_n2688# 0.18678f
C55 plus.n7 a_n2524_n2688# 0.009076f
C56 plus.n8 a_n2524_n2688# 0.352885f
C57 plus.n9 a_n2524_n2688# 0.355597f
C58 plus.n10 a_n2524_n2688# 0.079989f
C59 plus.n11 a_n2524_n2688# 0.066616f
C60 plus.n12 a_n2524_n2688# 0.053368f
C61 plus.n13 a_n2524_n2688# 0.009076f
C62 plus.n14 a_n2524_n2688# 0.343316f
C63 plus.n15 a_n2524_n2688# 0.009076f
C64 plus.n16 a_n2524_n2688# 0.344302f
C65 plus.n17 a_n2524_n2688# 0.414635f
C66 plus.n18 a_n2524_n2688# 0.039995f
C67 plus.t2 a_n2524_n2688# 0.825831f
C68 plus.n19 a_n2524_n2688# 0.039995f
C69 plus.t9 a_n2524_n2688# 0.825831f
C70 plus.t3 a_n2524_n2688# 0.825831f
C71 plus.n20 a_n2524_n2688# 0.352885f
C72 plus.n21 a_n2524_n2688# 0.066616f
C73 plus.t0 a_n2524_n2688# 0.825831f
C74 plus.t4 a_n2524_n2688# 0.825831f
C75 plus.t1 a_n2524_n2688# 0.825831f
C76 plus.n22 a_n2524_n2688# 0.34827f
C77 plus.t5 a_n2524_n2688# 0.849799f
C78 plus.n23 a_n2524_n2688# 0.325329f
C79 plus.n24 a_n2524_n2688# 0.18678f
C80 plus.n25 a_n2524_n2688# 0.009076f
C81 plus.n26 a_n2524_n2688# 0.352885f
C82 plus.n27 a_n2524_n2688# 0.355597f
C83 plus.n28 a_n2524_n2688# 0.079989f
C84 plus.n29 a_n2524_n2688# 0.066616f
C85 plus.n30 a_n2524_n2688# 0.053368f
C86 plus.n31 a_n2524_n2688# 0.009076f
C87 plus.n32 a_n2524_n2688# 0.343316f
C88 plus.n33 a_n2524_n2688# 0.009076f
C89 plus.n34 a_n2524_n2688# 0.344302f
C90 plus.n35 a_n2524_n2688# 1.26974f
C91 source.t10 a_n2524_n2688# 2.0127f
C92 source.n0 a_n2524_n2688# 1.21897f
C93 source.t11 a_n2524_n2688# 0.188747f
C94 source.t4 a_n2524_n2688# 0.188747f
C95 source.n1 a_n2524_n2688# 1.58007f
C96 source.n2 a_n2524_n2688# 0.413954f
C97 source.t0 a_n2524_n2688# 0.188747f
C98 source.t7 a_n2524_n2688# 0.188747f
C99 source.n3 a_n2524_n2688# 1.58007f
C100 source.n4 a_n2524_n2688# 0.413954f
C101 source.t3 a_n2524_n2688# 0.188747f
C102 source.t9 a_n2524_n2688# 0.188747f
C103 source.n5 a_n2524_n2688# 1.58007f
C104 source.n6 a_n2524_n2688# 0.412479f
C105 source.t19 a_n2524_n2688# 2.0127f
C106 source.n7 a_n2524_n2688# 0.494609f
C107 source.t24 a_n2524_n2688# 0.188747f
C108 source.t23 a_n2524_n2688# 0.188747f
C109 source.n8 a_n2524_n2688# 1.58007f
C110 source.n9 a_n2524_n2688# 0.413954f
C111 source.t16 a_n2524_n2688# 0.188747f
C112 source.t17 a_n2524_n2688# 0.188747f
C113 source.n10 a_n2524_n2688# 1.58007f
C114 source.n11 a_n2524_n2688# 0.413954f
C115 source.t21 a_n2524_n2688# 0.188747f
C116 source.t18 a_n2524_n2688# 0.188747f
C117 source.n12 a_n2524_n2688# 1.58007f
C118 source.n13 a_n2524_n2688# 1.61786f
C119 source.t12 a_n2524_n2688# 0.188747f
C120 source.t1 a_n2524_n2688# 0.188747f
C121 source.n14 a_n2524_n2688# 1.58006f
C122 source.n15 a_n2524_n2688# 1.61786f
C123 source.t13 a_n2524_n2688# 0.188747f
C124 source.t2 a_n2524_n2688# 0.188747f
C125 source.n16 a_n2524_n2688# 1.58006f
C126 source.n17 a_n2524_n2688# 0.413959f
C127 source.t6 a_n2524_n2688# 0.188747f
C128 source.t8 a_n2524_n2688# 0.188747f
C129 source.n18 a_n2524_n2688# 1.58006f
C130 source.n19 a_n2524_n2688# 0.413959f
C131 source.t5 a_n2524_n2688# 2.0127f
C132 source.n20 a_n2524_n2688# 0.494614f
C133 source.t14 a_n2524_n2688# 0.188747f
C134 source.t25 a_n2524_n2688# 0.188747f
C135 source.n21 a_n2524_n2688# 1.58006f
C136 source.n22 a_n2524_n2688# 0.412484f
C137 source.t20 a_n2524_n2688# 0.188747f
C138 source.t26 a_n2524_n2688# 0.188747f
C139 source.n23 a_n2524_n2688# 1.58006f
C140 source.n24 a_n2524_n2688# 0.413959f
C141 source.t15 a_n2524_n2688# 0.188747f
C142 source.t27 a_n2524_n2688# 0.188747f
C143 source.n25 a_n2524_n2688# 1.58006f
C144 source.n26 a_n2524_n2688# 0.413959f
C145 source.t22 a_n2524_n2688# 2.0127f
C146 source.n27 a_n2524_n2688# 0.631823f
C147 source.n28 a_n2524_n2688# 1.40146f
C148 drain_right.t6 a_n2524_n2688# 1.93713f
C149 drain_right.t8 a_n2524_n2688# 0.173553f
C150 drain_right.t9 a_n2524_n2688# 0.173553f
C151 drain_right.n0 a_n2524_n2688# 1.51801f
C152 drain_right.n1 a_n2524_n2688# 0.662096f
C153 drain_right.t11 a_n2524_n2688# 0.173553f
C154 drain_right.t2 a_n2524_n2688# 0.173553f
C155 drain_right.n2 a_n2524_n2688# 1.52326f
C156 drain_right.t12 a_n2524_n2688# 0.173553f
C157 drain_right.t4 a_n2524_n2688# 0.173553f
C158 drain_right.n3 a_n2524_n2688# 1.51801f
C159 drain_right.n4 a_n2524_n2688# 0.643107f
C160 drain_right.n5 a_n2524_n2688# 1.17839f
C161 drain_right.t13 a_n2524_n2688# 0.173553f
C162 drain_right.t3 a_n2524_n2688# 0.173553f
C163 drain_right.n6 a_n2524_n2688# 1.52325f
C164 drain_right.t1 a_n2524_n2688# 0.173553f
C165 drain_right.t7 a_n2524_n2688# 0.173553f
C166 drain_right.n7 a_n2524_n2688# 1.51801f
C167 drain_right.n8 a_n2524_n2688# 0.701901f
C168 drain_right.t5 a_n2524_n2688# 0.173553f
C169 drain_right.t10 a_n2524_n2688# 0.173553f
C170 drain_right.n9 a_n2524_n2688# 1.51801f
C171 drain_right.n10 a_n2524_n2688# 0.348658f
C172 drain_right.t0 a_n2524_n2688# 1.9323f
C173 drain_right.n11 a_n2524_n2688# 0.570313f
C174 minus.n0 a_n2524_n2688# 0.039272f
C175 minus.n1 a_n2524_n2688# 0.008912f
C176 minus.t9 a_n2524_n2688# 0.81091f
C177 minus.n2 a_n2524_n2688# 0.078544f
C178 minus.n3 a_n2524_n2688# 0.008912f
C179 minus.t3 a_n2524_n2688# 0.81091f
C180 minus.t8 a_n2524_n2688# 0.834445f
C181 minus.t4 a_n2524_n2688# 0.81091f
C182 minus.n4 a_n2524_n2688# 0.341978f
C183 minus.n5 a_n2524_n2688# 0.319451f
C184 minus.n6 a_n2524_n2688# 0.183405f
C185 minus.n7 a_n2524_n2688# 0.065412f
C186 minus.n8 a_n2524_n2688# 0.346509f
C187 minus.t10 a_n2524_n2688# 0.81091f
C188 minus.n9 a_n2524_n2688# 0.349172f
C189 minus.t11 a_n2524_n2688# 0.81091f
C190 minus.n10 a_n2524_n2688# 0.346509f
C191 minus.n11 a_n2524_n2688# 0.065412f
C192 minus.n12 a_n2524_n2688# 0.052403f
C193 minus.n13 a_n2524_n2688# 0.039272f
C194 minus.n14 a_n2524_n2688# 0.337113f
C195 minus.n15 a_n2524_n2688# 0.008912f
C196 minus.t6 a_n2524_n2688# 0.81091f
C197 minus.n16 a_n2524_n2688# 0.338082f
C198 minus.n17 a_n2524_n2688# 1.42115f
C199 minus.n18 a_n2524_n2688# 0.039272f
C200 minus.n19 a_n2524_n2688# 0.008912f
C201 minus.n20 a_n2524_n2688# 0.078544f
C202 minus.n21 a_n2524_n2688# 0.008912f
C203 minus.t13 a_n2524_n2688# 0.834445f
C204 minus.t2 a_n2524_n2688# 0.81091f
C205 minus.n22 a_n2524_n2688# 0.341978f
C206 minus.n23 a_n2524_n2688# 0.319451f
C207 minus.n24 a_n2524_n2688# 0.183405f
C208 minus.n25 a_n2524_n2688# 0.065412f
C209 minus.t7 a_n2524_n2688# 0.81091f
C210 minus.n26 a_n2524_n2688# 0.346509f
C211 minus.t1 a_n2524_n2688# 0.81091f
C212 minus.n27 a_n2524_n2688# 0.349172f
C213 minus.t12 a_n2524_n2688# 0.81091f
C214 minus.n28 a_n2524_n2688# 0.346509f
C215 minus.n29 a_n2524_n2688# 0.065412f
C216 minus.n30 a_n2524_n2688# 0.052403f
C217 minus.n31 a_n2524_n2688# 0.039272f
C218 minus.t0 a_n2524_n2688# 0.81091f
C219 minus.n32 a_n2524_n2688# 0.337113f
C220 minus.n33 a_n2524_n2688# 0.008912f
C221 minus.t5 a_n2524_n2688# 0.81091f
C222 minus.n34 a_n2524_n2688# 0.338082f
C223 minus.n35 a_n2524_n2688# 0.277431f
C224 minus.n36 a_n2524_n2688# 1.71728f
.ends

