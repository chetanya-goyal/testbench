* NGSPICE file created from diffpair517.ext - technology: sky130A

.subckt diffpair517 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t29 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X1 source.t13 minus.t0 drain_right.t15 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X2 drain_left.t14 plus.t1 source.t19 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X3 drain_left.t13 plus.t2 source.t24 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X4 drain_right.t14 minus.t1 source.t1 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X5 a_n1850_n3888# a_n1850_n3888# a_n1850_n3888# a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.3
X6 source.t16 plus.t3 drain_left.t12 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X7 source.t8 minus.t2 drain_right.t13 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X8 source.t11 minus.t3 drain_right.t12 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X9 drain_right.t11 minus.t4 source.t6 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X10 drain_left.t11 plus.t4 source.t21 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X11 drain_left.t10 plus.t5 source.t26 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X12 source.t27 plus.t6 drain_left.t9 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X13 drain_left.t8 plus.t7 source.t22 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X14 a_n1850_n3888# a_n1850_n3888# a_n1850_n3888# a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X15 source.t9 minus.t5 drain_right.t10 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X16 source.t5 minus.t6 drain_right.t9 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X17 source.t10 minus.t7 drain_right.t8 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X18 drain_right.t7 minus.t8 source.t12 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X19 drain_left.t7 plus.t8 source.t31 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X20 a_n1850_n3888# a_n1850_n3888# a_n1850_n3888# a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X21 source.t25 plus.t9 drain_left.t6 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X22 source.t17 plus.t10 drain_left.t5 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X23 source.t18 plus.t11 drain_left.t4 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X24 source.t23 plus.t12 drain_left.t3 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X25 a_n1850_n3888# a_n1850_n3888# a_n1850_n3888# a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X26 drain_right.t6 minus.t9 source.t3 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X27 drain_right.t5 minus.t10 source.t0 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X28 drain_right.t4 minus.t11 source.t2 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X29 source.t4 minus.t12 drain_right.t3 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X30 source.t14 minus.t13 drain_right.t2 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X31 source.t20 plus.t13 drain_left.t2 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X32 drain_right.t1 minus.t14 source.t7 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X33 drain_right.t0 minus.t15 source.t15 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X34 source.t30 plus.t14 drain_left.t1 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X35 drain_left.t0 plus.t15 source.t28 a_n1850_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
R0 plus.n5 plus.t3 1339.38
R1 plus.n21 plus.t0 1339.38
R2 plus.n28 plus.t1 1339.38
R3 plus.n44 plus.t14 1339.38
R4 plus.n6 plus.t7 1309.43
R5 plus.n3 plus.t10 1309.43
R6 plus.n12 plus.t15 1309.43
R7 plus.n14 plus.t6 1309.43
R8 plus.n1 plus.t8 1309.43
R9 plus.n20 plus.t13 1309.43
R10 plus.n29 plus.t9 1309.43
R11 plus.n26 plus.t2 1309.43
R12 plus.n35 plus.t11 1309.43
R13 plus.n37 plus.t4 1309.43
R14 plus.n24 plus.t12 1309.43
R15 plus.n43 plus.t5 1309.43
R16 plus.n5 plus.n4 161.489
R17 plus.n28 plus.n27 161.489
R18 plus.n7 plus.n4 161.3
R19 plus.n9 plus.n8 161.3
R20 plus.n11 plus.n10 161.3
R21 plus.n13 plus.n2 161.3
R22 plus.n16 plus.n15 161.3
R23 plus.n18 plus.n17 161.3
R24 plus.n19 plus.n0 161.3
R25 plus.n22 plus.n21 161.3
R26 plus.n30 plus.n27 161.3
R27 plus.n32 plus.n31 161.3
R28 plus.n34 plus.n33 161.3
R29 plus.n36 plus.n25 161.3
R30 plus.n39 plus.n38 161.3
R31 plus.n41 plus.n40 161.3
R32 plus.n42 plus.n23 161.3
R33 plus.n45 plus.n44 161.3
R34 plus.n8 plus.n7 73.0308
R35 plus.n19 plus.n18 73.0308
R36 plus.n42 plus.n41 73.0308
R37 plus.n31 plus.n30 73.0308
R38 plus.n11 plus.n3 64.9975
R39 plus.n15 plus.n1 64.9975
R40 plus.n38 plus.n24 64.9975
R41 plus.n34 plus.n26 64.9975
R42 plus.n6 plus.n5 62.0763
R43 plus.n21 plus.n20 62.0763
R44 plus.n44 plus.n43 62.0763
R45 plus.n29 plus.n28 62.0763
R46 plus.n13 plus.n12 46.0096
R47 plus.n14 plus.n13 46.0096
R48 plus.n37 plus.n36 46.0096
R49 plus.n36 plus.n35 46.0096
R50 plus plus.n45 31.1127
R51 plus.n12 plus.n11 27.0217
R52 plus.n15 plus.n14 27.0217
R53 plus.n38 plus.n37 27.0217
R54 plus.n35 plus.n34 27.0217
R55 plus plus.n22 13.2467
R56 plus.n7 plus.n6 10.955
R57 plus.n20 plus.n19 10.955
R58 plus.n43 plus.n42 10.955
R59 plus.n30 plus.n29 10.955
R60 plus.n8 plus.n3 8.03383
R61 plus.n18 plus.n1 8.03383
R62 plus.n41 plus.n24 8.03383
R63 plus.n31 plus.n26 8.03383
R64 plus.n9 plus.n4 0.189894
R65 plus.n10 plus.n9 0.189894
R66 plus.n10 plus.n2 0.189894
R67 plus.n16 plus.n2 0.189894
R68 plus.n17 plus.n16 0.189894
R69 plus.n17 plus.n0 0.189894
R70 plus.n22 plus.n0 0.189894
R71 plus.n45 plus.n23 0.189894
R72 plus.n40 plus.n23 0.189894
R73 plus.n40 plus.n39 0.189894
R74 plus.n39 plus.n25 0.189894
R75 plus.n33 plus.n25 0.189894
R76 plus.n33 plus.n32 0.189894
R77 plus.n32 plus.n27 0.189894
R78 source.n7 source.t16 45.521
R79 source.n8 source.t12 45.521
R80 source.n15 source.t14 45.521
R81 source.n31 source.t7 45.5208
R82 source.n24 source.t11 45.5208
R83 source.n23 source.t19 45.5208
R84 source.n16 source.t30 45.5208
R85 source.n0 source.t29 45.5208
R86 source.n2 source.n1 44.201
R87 source.n4 source.n3 44.201
R88 source.n6 source.n5 44.201
R89 source.n10 source.n9 44.201
R90 source.n12 source.n11 44.201
R91 source.n14 source.n13 44.201
R92 source.n30 source.n29 44.2008
R93 source.n28 source.n27 44.2008
R94 source.n26 source.n25 44.2008
R95 source.n22 source.n21 44.2008
R96 source.n20 source.n19 44.2008
R97 source.n18 source.n17 44.2008
R98 source.n16 source.n15 24.1036
R99 source.n32 source.n0 18.5691
R100 source.n32 source.n31 5.53498
R101 source.n29 source.t15 1.3205
R102 source.n29 source.t5 1.3205
R103 source.n27 source.t0 1.3205
R104 source.n27 source.t10 1.3205
R105 source.n25 source.t2 1.3205
R106 source.n25 source.t8 1.3205
R107 source.n21 source.t24 1.3205
R108 source.n21 source.t25 1.3205
R109 source.n19 source.t21 1.3205
R110 source.n19 source.t18 1.3205
R111 source.n17 source.t26 1.3205
R112 source.n17 source.t23 1.3205
R113 source.n1 source.t31 1.3205
R114 source.n1 source.t20 1.3205
R115 source.n3 source.t28 1.3205
R116 source.n3 source.t27 1.3205
R117 source.n5 source.t22 1.3205
R118 source.n5 source.t17 1.3205
R119 source.n9 source.t1 1.3205
R120 source.n9 source.t4 1.3205
R121 source.n11 source.t3 1.3205
R122 source.n11 source.t9 1.3205
R123 source.n13 source.t6 1.3205
R124 source.n13 source.t13 1.3205
R125 source.n15 source.n14 0.543603
R126 source.n14 source.n12 0.543603
R127 source.n12 source.n10 0.543603
R128 source.n10 source.n8 0.543603
R129 source.n7 source.n6 0.543603
R130 source.n6 source.n4 0.543603
R131 source.n4 source.n2 0.543603
R132 source.n2 source.n0 0.543603
R133 source.n18 source.n16 0.543603
R134 source.n20 source.n18 0.543603
R135 source.n22 source.n20 0.543603
R136 source.n23 source.n22 0.543603
R137 source.n26 source.n24 0.543603
R138 source.n28 source.n26 0.543603
R139 source.n30 source.n28 0.543603
R140 source.n31 source.n30 0.543603
R141 source.n8 source.n7 0.470328
R142 source.n24 source.n23 0.470328
R143 source source.n32 0.188
R144 drain_left.n9 drain_left.n7 61.4229
R145 drain_left.n5 drain_left.n3 61.4227
R146 drain_left.n2 drain_left.n0 61.4227
R147 drain_left.n11 drain_left.n10 60.8798
R148 drain_left.n9 drain_left.n8 60.8798
R149 drain_left.n13 drain_left.n12 60.8796
R150 drain_left.n5 drain_left.n4 60.8796
R151 drain_left.n2 drain_left.n1 60.8796
R152 drain_left drain_left.n6 33.17
R153 drain_left drain_left.n13 6.19632
R154 drain_left.n3 drain_left.t6 1.3205
R155 drain_left.n3 drain_left.t14 1.3205
R156 drain_left.n4 drain_left.t4 1.3205
R157 drain_left.n4 drain_left.t13 1.3205
R158 drain_left.n1 drain_left.t3 1.3205
R159 drain_left.n1 drain_left.t11 1.3205
R160 drain_left.n0 drain_left.t1 1.3205
R161 drain_left.n0 drain_left.t10 1.3205
R162 drain_left.n12 drain_left.t2 1.3205
R163 drain_left.n12 drain_left.t15 1.3205
R164 drain_left.n10 drain_left.t9 1.3205
R165 drain_left.n10 drain_left.t7 1.3205
R166 drain_left.n8 drain_left.t5 1.3205
R167 drain_left.n8 drain_left.t0 1.3205
R168 drain_left.n7 drain_left.t12 1.3205
R169 drain_left.n7 drain_left.t8 1.3205
R170 drain_left.n11 drain_left.n9 0.543603
R171 drain_left.n13 drain_left.n11 0.543603
R172 drain_left.n6 drain_left.n5 0.216706
R173 drain_left.n6 drain_left.n2 0.216706
R174 minus.n21 minus.t13 1339.38
R175 minus.n5 minus.t8 1339.38
R176 minus.n44 minus.t14 1339.38
R177 minus.n28 minus.t3 1339.38
R178 minus.n20 minus.t4 1309.43
R179 minus.n1 minus.t0 1309.43
R180 minus.n14 minus.t9 1309.43
R181 minus.n12 minus.t5 1309.43
R182 minus.n3 minus.t1 1309.43
R183 minus.n6 minus.t12 1309.43
R184 minus.n43 minus.t6 1309.43
R185 minus.n24 minus.t15 1309.43
R186 minus.n37 minus.t7 1309.43
R187 minus.n35 minus.t10 1309.43
R188 minus.n26 minus.t2 1309.43
R189 minus.n29 minus.t11 1309.43
R190 minus.n5 minus.n4 161.489
R191 minus.n28 minus.n27 161.489
R192 minus.n22 minus.n21 161.3
R193 minus.n19 minus.n0 161.3
R194 minus.n18 minus.n17 161.3
R195 minus.n16 minus.n15 161.3
R196 minus.n13 minus.n2 161.3
R197 minus.n11 minus.n10 161.3
R198 minus.n9 minus.n8 161.3
R199 minus.n7 minus.n4 161.3
R200 minus.n45 minus.n44 161.3
R201 minus.n42 minus.n23 161.3
R202 minus.n41 minus.n40 161.3
R203 minus.n39 minus.n38 161.3
R204 minus.n36 minus.n25 161.3
R205 minus.n34 minus.n33 161.3
R206 minus.n32 minus.n31 161.3
R207 minus.n30 minus.n27 161.3
R208 minus.n19 minus.n18 73.0308
R209 minus.n8 minus.n7 73.0308
R210 minus.n31 minus.n30 73.0308
R211 minus.n42 minus.n41 73.0308
R212 minus.n15 minus.n1 64.9975
R213 minus.n11 minus.n3 64.9975
R214 minus.n34 minus.n26 64.9975
R215 minus.n38 minus.n24 64.9975
R216 minus.n21 minus.n20 62.0763
R217 minus.n6 minus.n5 62.0763
R218 minus.n29 minus.n28 62.0763
R219 minus.n44 minus.n43 62.0763
R220 minus.n14 minus.n13 46.0096
R221 minus.n13 minus.n12 46.0096
R222 minus.n36 minus.n35 46.0096
R223 minus.n37 minus.n36 46.0096
R224 minus.n46 minus.n22 38.3679
R225 minus.n15 minus.n14 27.0217
R226 minus.n12 minus.n11 27.0217
R227 minus.n35 minus.n34 27.0217
R228 minus.n38 minus.n37 27.0217
R229 minus.n20 minus.n19 10.955
R230 minus.n7 minus.n6 10.955
R231 minus.n30 minus.n29 10.955
R232 minus.n43 minus.n42 10.955
R233 minus.n18 minus.n1 8.03383
R234 minus.n8 minus.n3 8.03383
R235 minus.n31 minus.n26 8.03383
R236 minus.n41 minus.n24 8.03383
R237 minus.n46 minus.n45 6.46641
R238 minus.n22 minus.n0 0.189894
R239 minus.n17 minus.n0 0.189894
R240 minus.n17 minus.n16 0.189894
R241 minus.n16 minus.n2 0.189894
R242 minus.n10 minus.n2 0.189894
R243 minus.n10 minus.n9 0.189894
R244 minus.n9 minus.n4 0.189894
R245 minus.n32 minus.n27 0.189894
R246 minus.n33 minus.n32 0.189894
R247 minus.n33 minus.n25 0.189894
R248 minus.n39 minus.n25 0.189894
R249 minus.n40 minus.n39 0.189894
R250 minus.n40 minus.n23 0.189894
R251 minus.n45 minus.n23 0.189894
R252 minus minus.n46 0.188
R253 drain_right.n9 drain_right.n7 61.4227
R254 drain_right.n5 drain_right.n3 61.4227
R255 drain_right.n2 drain_right.n0 61.4227
R256 drain_right.n9 drain_right.n8 60.8798
R257 drain_right.n11 drain_right.n10 60.8798
R258 drain_right.n13 drain_right.n12 60.8798
R259 drain_right.n5 drain_right.n4 60.8796
R260 drain_right.n2 drain_right.n1 60.8796
R261 drain_right drain_right.n6 32.6167
R262 drain_right drain_right.n13 6.19632
R263 drain_right.n3 drain_right.t9 1.3205
R264 drain_right.n3 drain_right.t1 1.3205
R265 drain_right.n4 drain_right.t8 1.3205
R266 drain_right.n4 drain_right.t0 1.3205
R267 drain_right.n1 drain_right.t13 1.3205
R268 drain_right.n1 drain_right.t5 1.3205
R269 drain_right.n0 drain_right.t12 1.3205
R270 drain_right.n0 drain_right.t4 1.3205
R271 drain_right.n7 drain_right.t3 1.3205
R272 drain_right.n7 drain_right.t7 1.3205
R273 drain_right.n8 drain_right.t10 1.3205
R274 drain_right.n8 drain_right.t14 1.3205
R275 drain_right.n10 drain_right.t15 1.3205
R276 drain_right.n10 drain_right.t6 1.3205
R277 drain_right.n12 drain_right.t2 1.3205
R278 drain_right.n12 drain_right.t11 1.3205
R279 drain_right.n13 drain_right.n11 0.543603
R280 drain_right.n11 drain_right.n9 0.543603
R281 drain_right.n6 drain_right.n5 0.216706
R282 drain_right.n6 drain_right.n2 0.216706
C0 drain_right drain_left 0.948737f
C1 plus minus 6.01864f
C2 plus drain_left 7.425271f
C3 drain_left minus 0.171647f
C4 drain_right source 37.417603f
C5 plus source 6.83162f
C6 minus source 6.81758f
C7 drain_right plus 0.334364f
C8 drain_left source 37.4173f
C9 drain_right minus 7.24557f
C10 drain_right a_n1850_n3888# 7.222049f
C11 drain_left a_n1850_n3888# 7.509969f
C12 source a_n1850_n3888# 10.338611f
C13 minus a_n1850_n3888# 7.433937f
C14 plus a_n1850_n3888# 9.60645f
C15 drain_right.t12 a_n1850_n3888# 0.403362f
C16 drain_right.t4 a_n1850_n3888# 0.403362f
C17 drain_right.n0 a_n1850_n3888# 3.64956f
C18 drain_right.t13 a_n1850_n3888# 0.403362f
C19 drain_right.t5 a_n1850_n3888# 0.403362f
C20 drain_right.n1 a_n1850_n3888# 3.64592f
C21 drain_right.n2 a_n1850_n3888# 0.773513f
C22 drain_right.t9 a_n1850_n3888# 0.403362f
C23 drain_right.t1 a_n1850_n3888# 0.403362f
C24 drain_right.n3 a_n1850_n3888# 3.64956f
C25 drain_right.t8 a_n1850_n3888# 0.403362f
C26 drain_right.t0 a_n1850_n3888# 0.403362f
C27 drain_right.n4 a_n1850_n3888# 3.64592f
C28 drain_right.n5 a_n1850_n3888# 0.773513f
C29 drain_right.n6 a_n1850_n3888# 1.83971f
C30 drain_right.t3 a_n1850_n3888# 0.403362f
C31 drain_right.t7 a_n1850_n3888# 0.403362f
C32 drain_right.n7 a_n1850_n3888# 3.64955f
C33 drain_right.t10 a_n1850_n3888# 0.403362f
C34 drain_right.t14 a_n1850_n3888# 0.403362f
C35 drain_right.n8 a_n1850_n3888# 3.64592f
C36 drain_right.n9 a_n1850_n3888# 0.805715f
C37 drain_right.t15 a_n1850_n3888# 0.403362f
C38 drain_right.t6 a_n1850_n3888# 0.403362f
C39 drain_right.n10 a_n1850_n3888# 3.64592f
C40 drain_right.n11 a_n1850_n3888# 0.397817f
C41 drain_right.t2 a_n1850_n3888# 0.403362f
C42 drain_right.t11 a_n1850_n3888# 0.403362f
C43 drain_right.n12 a_n1850_n3888# 3.64592f
C44 drain_right.n13 a_n1850_n3888# 0.681062f
C45 minus.n0 a_n1850_n3888# 0.050385f
C46 minus.t13 a_n1850_n3888# 0.645146f
C47 minus.t4 a_n1850_n3888# 0.63965f
C48 minus.t0 a_n1850_n3888# 0.63965f
C49 minus.n1 a_n1850_n3888# 0.245693f
C50 minus.n2 a_n1850_n3888# 0.050385f
C51 minus.t9 a_n1850_n3888# 0.63965f
C52 minus.t5 a_n1850_n3888# 0.63965f
C53 minus.t1 a_n1850_n3888# 0.63965f
C54 minus.n3 a_n1850_n3888# 0.245693f
C55 minus.n4 a_n1850_n3888# 0.107227f
C56 minus.t12 a_n1850_n3888# 0.63965f
C57 minus.t8 a_n1850_n3888# 0.645146f
C58 minus.n5 a_n1850_n3888# 0.261172f
C59 minus.n6 a_n1850_n3888# 0.245693f
C60 minus.n7 a_n1850_n3888# 0.019044f
C61 minus.n8 a_n1850_n3888# 0.018423f
C62 minus.n9 a_n1850_n3888# 0.050385f
C63 minus.n10 a_n1850_n3888# 0.050385f
C64 minus.n11 a_n1850_n3888# 0.020753f
C65 minus.n12 a_n1850_n3888# 0.245693f
C66 minus.n13 a_n1850_n3888# 0.020753f
C67 minus.n14 a_n1850_n3888# 0.245693f
C68 minus.n15 a_n1850_n3888# 0.020753f
C69 minus.n16 a_n1850_n3888# 0.050385f
C70 minus.n17 a_n1850_n3888# 0.050385f
C71 minus.n18 a_n1850_n3888# 0.018423f
C72 minus.n19 a_n1850_n3888# 0.019044f
C73 minus.n20 a_n1850_n3888# 0.245693f
C74 minus.n21 a_n1850_n3888# 0.261106f
C75 minus.n22 a_n1850_n3888# 1.94731f
C76 minus.n23 a_n1850_n3888# 0.050385f
C77 minus.t6 a_n1850_n3888# 0.63965f
C78 minus.t15 a_n1850_n3888# 0.63965f
C79 minus.n24 a_n1850_n3888# 0.245693f
C80 minus.n25 a_n1850_n3888# 0.050385f
C81 minus.t7 a_n1850_n3888# 0.63965f
C82 minus.t10 a_n1850_n3888# 0.63965f
C83 minus.t2 a_n1850_n3888# 0.63965f
C84 minus.n26 a_n1850_n3888# 0.245693f
C85 minus.n27 a_n1850_n3888# 0.107227f
C86 minus.t11 a_n1850_n3888# 0.63965f
C87 minus.t3 a_n1850_n3888# 0.645146f
C88 minus.n28 a_n1850_n3888# 0.261172f
C89 minus.n29 a_n1850_n3888# 0.245693f
C90 minus.n30 a_n1850_n3888# 0.019044f
C91 minus.n31 a_n1850_n3888# 0.018423f
C92 minus.n32 a_n1850_n3888# 0.050385f
C93 minus.n33 a_n1850_n3888# 0.050385f
C94 minus.n34 a_n1850_n3888# 0.020753f
C95 minus.n35 a_n1850_n3888# 0.245693f
C96 minus.n36 a_n1850_n3888# 0.020753f
C97 minus.n37 a_n1850_n3888# 0.245693f
C98 minus.n38 a_n1850_n3888# 0.020753f
C99 minus.n39 a_n1850_n3888# 0.050385f
C100 minus.n40 a_n1850_n3888# 0.050385f
C101 minus.n41 a_n1850_n3888# 0.018423f
C102 minus.n42 a_n1850_n3888# 0.019044f
C103 minus.n43 a_n1850_n3888# 0.245693f
C104 minus.t14 a_n1850_n3888# 0.645146f
C105 minus.n44 a_n1850_n3888# 0.261106f
C106 minus.n45 a_n1850_n3888# 0.325412f
C107 minus.n46 a_n1850_n3888# 2.35146f
C108 drain_left.t1 a_n1850_n3888# 0.403965f
C109 drain_left.t10 a_n1850_n3888# 0.403965f
C110 drain_left.n0 a_n1850_n3888# 3.65502f
C111 drain_left.t3 a_n1850_n3888# 0.403965f
C112 drain_left.t11 a_n1850_n3888# 0.403965f
C113 drain_left.n1 a_n1850_n3888# 3.65137f
C114 drain_left.n2 a_n1850_n3888# 0.77467f
C115 drain_left.t6 a_n1850_n3888# 0.403965f
C116 drain_left.t14 a_n1850_n3888# 0.403965f
C117 drain_left.n3 a_n1850_n3888# 3.65502f
C118 drain_left.t4 a_n1850_n3888# 0.403965f
C119 drain_left.t13 a_n1850_n3888# 0.403965f
C120 drain_left.n4 a_n1850_n3888# 3.65137f
C121 drain_left.n5 a_n1850_n3888# 0.77467f
C122 drain_left.n6 a_n1850_n3888# 1.91338f
C123 drain_left.t12 a_n1850_n3888# 0.403965f
C124 drain_left.t8 a_n1850_n3888# 0.403965f
C125 drain_left.n7 a_n1850_n3888# 3.65502f
C126 drain_left.t5 a_n1850_n3888# 0.403965f
C127 drain_left.t0 a_n1850_n3888# 0.403965f
C128 drain_left.n8 a_n1850_n3888# 3.65137f
C129 drain_left.n9 a_n1850_n3888# 0.806907f
C130 drain_left.t9 a_n1850_n3888# 0.403965f
C131 drain_left.t7 a_n1850_n3888# 0.403965f
C132 drain_left.n10 a_n1850_n3888# 3.65137f
C133 drain_left.n11 a_n1850_n3888# 0.398412f
C134 drain_left.t2 a_n1850_n3888# 0.403965f
C135 drain_left.t15 a_n1850_n3888# 0.403965f
C136 drain_left.n12 a_n1850_n3888# 3.65136f
C137 drain_left.n13 a_n1850_n3888# 0.682093f
C138 source.t29 a_n1850_n3888# 3.74121f
C139 source.n0 a_n1850_n3888# 1.73285f
C140 source.t31 a_n1850_n3888# 0.33384f
C141 source.t20 a_n1850_n3888# 0.33384f
C142 source.n1 a_n1850_n3888# 2.9325f
C143 source.n2 a_n1850_n3888# 0.375991f
C144 source.t28 a_n1850_n3888# 0.33384f
C145 source.t27 a_n1850_n3888# 0.33384f
C146 source.n3 a_n1850_n3888# 2.9325f
C147 source.n4 a_n1850_n3888# 0.375991f
C148 source.t22 a_n1850_n3888# 0.33384f
C149 source.t17 a_n1850_n3888# 0.33384f
C150 source.n5 a_n1850_n3888# 2.9325f
C151 source.n6 a_n1850_n3888# 0.375991f
C152 source.t16 a_n1850_n3888# 3.74121f
C153 source.n7 a_n1850_n3888# 0.471099f
C154 source.t12 a_n1850_n3888# 3.74121f
C155 source.n8 a_n1850_n3888# 0.471099f
C156 source.t1 a_n1850_n3888# 0.33384f
C157 source.t4 a_n1850_n3888# 0.33384f
C158 source.n9 a_n1850_n3888# 2.9325f
C159 source.n10 a_n1850_n3888# 0.375991f
C160 source.t3 a_n1850_n3888# 0.33384f
C161 source.t9 a_n1850_n3888# 0.33384f
C162 source.n11 a_n1850_n3888# 2.9325f
C163 source.n12 a_n1850_n3888# 0.375991f
C164 source.t6 a_n1850_n3888# 0.33384f
C165 source.t13 a_n1850_n3888# 0.33384f
C166 source.n13 a_n1850_n3888# 2.9325f
C167 source.n14 a_n1850_n3888# 0.375991f
C168 source.t14 a_n1850_n3888# 3.74121f
C169 source.n15 a_n1850_n3888# 2.2011f
C170 source.t30 a_n1850_n3888# 3.74121f
C171 source.n16 a_n1850_n3888# 2.20111f
C172 source.t26 a_n1850_n3888# 0.33384f
C173 source.t23 a_n1850_n3888# 0.33384f
C174 source.n17 a_n1850_n3888# 2.9325f
C175 source.n18 a_n1850_n3888# 0.375995f
C176 source.t21 a_n1850_n3888# 0.33384f
C177 source.t18 a_n1850_n3888# 0.33384f
C178 source.n19 a_n1850_n3888# 2.9325f
C179 source.n20 a_n1850_n3888# 0.375995f
C180 source.t24 a_n1850_n3888# 0.33384f
C181 source.t25 a_n1850_n3888# 0.33384f
C182 source.n21 a_n1850_n3888# 2.9325f
C183 source.n22 a_n1850_n3888# 0.375995f
C184 source.t19 a_n1850_n3888# 3.74121f
C185 source.n23 a_n1850_n3888# 0.471104f
C186 source.t11 a_n1850_n3888# 3.74121f
C187 source.n24 a_n1850_n3888# 0.471104f
C188 source.t2 a_n1850_n3888# 0.33384f
C189 source.t8 a_n1850_n3888# 0.33384f
C190 source.n25 a_n1850_n3888# 2.9325f
C191 source.n26 a_n1850_n3888# 0.375995f
C192 source.t0 a_n1850_n3888# 0.33384f
C193 source.t10 a_n1850_n3888# 0.33384f
C194 source.n27 a_n1850_n3888# 2.9325f
C195 source.n28 a_n1850_n3888# 0.375995f
C196 source.t15 a_n1850_n3888# 0.33384f
C197 source.t5 a_n1850_n3888# 0.33384f
C198 source.n29 a_n1850_n3888# 2.9325f
C199 source.n30 a_n1850_n3888# 0.375995f
C200 source.t7 a_n1850_n3888# 3.74121f
C201 source.n31 a_n1850_n3888# 0.630089f
C202 source.n32 a_n1850_n3888# 2.0593f
C203 plus.n0 a_n1850_n3888# 0.05115f
C204 plus.t13 a_n1850_n3888# 0.649355f
C205 plus.t8 a_n1850_n3888# 0.649355f
C206 plus.n1 a_n1850_n3888# 0.249421f
C207 plus.n2 a_n1850_n3888# 0.05115f
C208 plus.t6 a_n1850_n3888# 0.649355f
C209 plus.t15 a_n1850_n3888# 0.649355f
C210 plus.t10 a_n1850_n3888# 0.649355f
C211 plus.n3 a_n1850_n3888# 0.249421f
C212 plus.n4 a_n1850_n3888# 0.108854f
C213 plus.t7 a_n1850_n3888# 0.649355f
C214 plus.t3 a_n1850_n3888# 0.654935f
C215 plus.n5 a_n1850_n3888# 0.265135f
C216 plus.n6 a_n1850_n3888# 0.249421f
C217 plus.n7 a_n1850_n3888# 0.019333f
C218 plus.n8 a_n1850_n3888# 0.018702f
C219 plus.n9 a_n1850_n3888# 0.05115f
C220 plus.n10 a_n1850_n3888# 0.05115f
C221 plus.n11 a_n1850_n3888# 0.021068f
C222 plus.n12 a_n1850_n3888# 0.249421f
C223 plus.n13 a_n1850_n3888# 0.021068f
C224 plus.n14 a_n1850_n3888# 0.249421f
C225 plus.n15 a_n1850_n3888# 0.021068f
C226 plus.n16 a_n1850_n3888# 0.05115f
C227 plus.n17 a_n1850_n3888# 0.05115f
C228 plus.n18 a_n1850_n3888# 0.018702f
C229 plus.n19 a_n1850_n3888# 0.019333f
C230 plus.n20 a_n1850_n3888# 0.249421f
C231 plus.t0 a_n1850_n3888# 0.654935f
C232 plus.n21 a_n1850_n3888# 0.265067f
C233 plus.n22 a_n1850_n3888# 0.64232f
C234 plus.n23 a_n1850_n3888# 0.05115f
C235 plus.t14 a_n1850_n3888# 0.654935f
C236 plus.t5 a_n1850_n3888# 0.649355f
C237 plus.t12 a_n1850_n3888# 0.649355f
C238 plus.n24 a_n1850_n3888# 0.249421f
C239 plus.n25 a_n1850_n3888# 0.05115f
C240 plus.t4 a_n1850_n3888# 0.649355f
C241 plus.t11 a_n1850_n3888# 0.649355f
C242 plus.t2 a_n1850_n3888# 0.649355f
C243 plus.n26 a_n1850_n3888# 0.249421f
C244 plus.n27 a_n1850_n3888# 0.108854f
C245 plus.t9 a_n1850_n3888# 0.649355f
C246 plus.t1 a_n1850_n3888# 0.654935f
C247 plus.n28 a_n1850_n3888# 0.265135f
C248 plus.n29 a_n1850_n3888# 0.249421f
C249 plus.n30 a_n1850_n3888# 0.019333f
C250 plus.n31 a_n1850_n3888# 0.018702f
C251 plus.n32 a_n1850_n3888# 0.05115f
C252 plus.n33 a_n1850_n3888# 0.05115f
C253 plus.n34 a_n1850_n3888# 0.021068f
C254 plus.n35 a_n1850_n3888# 0.249421f
C255 plus.n36 a_n1850_n3888# 0.021068f
C256 plus.n37 a_n1850_n3888# 0.249421f
C257 plus.n38 a_n1850_n3888# 0.021068f
C258 plus.n39 a_n1850_n3888# 0.05115f
C259 plus.n40 a_n1850_n3888# 0.05115f
C260 plus.n41 a_n1850_n3888# 0.018702f
C261 plus.n42 a_n1850_n3888# 0.019333f
C262 plus.n43 a_n1850_n3888# 0.249421f
C263 plus.n44 a_n1850_n3888# 0.265067f
C264 plus.n45 a_n1850_n3888# 1.62581f
.ends

