* NGSPICE file created from diffpair587.ext - technology: sky130A

.subckt diffpair587 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t16 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X1 drain_left.t14 plus.t1 source.t25 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X2 drain_left.t13 plus.t2 source.t20 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X3 drain_right.t15 minus.t0 source.t3 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X4 a_n1760_n4888# a_n1760_n4888# a_n1760_n4888# a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.25
X5 source.t8 minus.t1 drain_right.t14 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X6 source.t1 minus.t2 drain_right.t13 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X7 drain_left.t12 plus.t3 source.t30 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X8 source.t10 minus.t3 drain_right.t12 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X9 source.t28 plus.t4 drain_left.t11 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X10 a_n1760_n4888# a_n1760_n4888# a_n1760_n4888# a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X11 source.t27 plus.t5 drain_left.t10 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X12 source.t13 minus.t4 drain_right.t11 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X13 drain_right.t10 minus.t5 source.t7 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X14 source.t9 minus.t6 drain_right.t9 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X15 drain_left.t9 plus.t6 source.t19 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X16 source.t12 minus.t7 drain_right.t8 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X17 source.t31 plus.t7 drain_left.t8 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X18 source.t23 plus.t8 drain_left.t7 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X19 source.t24 plus.t9 drain_left.t6 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X20 source.t17 plus.t10 drain_left.t5 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X21 a_n1760_n4888# a_n1760_n4888# a_n1760_n4888# a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X22 drain_left.t4 plus.t11 source.t26 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X23 drain_right.t7 minus.t8 source.t6 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X24 drain_right.t6 minus.t9 source.t15 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X25 a_n1760_n4888# a_n1760_n4888# a_n1760_n4888# a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X26 drain_right.t5 minus.t10 source.t4 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X27 drain_left.t3 plus.t12 source.t21 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X28 drain_right.t4 minus.t11 source.t0 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X29 drain_right.t3 minus.t12 source.t2 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X30 drain_right.t2 minus.t13 source.t5 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X31 source.t29 plus.t13 drain_left.t2 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X32 source.t11 minus.t14 drain_right.t1 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X33 source.t14 minus.t15 drain_right.t0 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X34 drain_left.t1 plus.t14 source.t18 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X35 source.t22 plus.t15 drain_left.t0 a_n1760_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
R0 plus.n4 plus.t5 2094.22
R1 plus.n19 plus.t3 2094.22
R2 plus.n25 plus.t2 2094.22
R3 plus.n40 plus.t7 2094.22
R4 plus.n5 plus.t1 2053.32
R5 plus.n3 plus.t10 2053.32
R6 plus.n10 plus.t0 2053.32
R7 plus.n1 plus.t9 2053.32
R8 plus.n16 plus.t14 2053.32
R9 plus.n18 plus.t8 2053.32
R10 plus.n26 plus.t13 2053.32
R11 plus.n24 plus.t11 2053.32
R12 plus.n31 plus.t4 2053.32
R13 plus.n22 plus.t6 2053.32
R14 plus.n37 plus.t15 2053.32
R15 plus.n39 plus.t12 2053.32
R16 plus.n7 plus.n4 161.489
R17 plus.n28 plus.n25 161.489
R18 plus.n7 plus.n6 161.3
R19 plus.n9 plus.n8 161.3
R20 plus.n11 plus.n2 161.3
R21 plus.n13 plus.n12 161.3
R22 plus.n15 plus.n14 161.3
R23 plus.n17 plus.n0 161.3
R24 plus.n20 plus.n19 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n29 161.3
R27 plus.n32 plus.n23 161.3
R28 plus.n34 plus.n33 161.3
R29 plus.n36 plus.n35 161.3
R30 plus.n38 plus.n21 161.3
R31 plus.n41 plus.n40 161.3
R32 plus.n12 plus.n11 73.0308
R33 plus.n33 plus.n32 73.0308
R34 plus.n10 plus.n9 67.1884
R35 plus.n15 plus.n1 67.1884
R36 plus.n36 plus.n22 67.1884
R37 plus.n31 plus.n30 67.1884
R38 plus.n6 plus.n3 55.5035
R39 plus.n17 plus.n16 55.5035
R40 plus.n38 plus.n37 55.5035
R41 plus.n27 plus.n24 55.5035
R42 plus.n5 plus.n4 43.8187
R43 plus.n19 plus.n18 43.8187
R44 plus.n40 plus.n39 43.8187
R45 plus.n26 plus.n25 43.8187
R46 plus plus.n41 32.6657
R47 plus.n6 plus.n5 29.2126
R48 plus.n18 plus.n17 29.2126
R49 plus.n39 plus.n38 29.2126
R50 plus.n27 plus.n26 29.2126
R51 plus.n9 plus.n3 17.5278
R52 plus.n16 plus.n15 17.5278
R53 plus.n37 plus.n36 17.5278
R54 plus.n30 plus.n24 17.5278
R55 plus plus.n20 15.1407
R56 plus.n11 plus.n10 5.84292
R57 plus.n12 plus.n1 5.84292
R58 plus.n33 plus.n22 5.84292
R59 plus.n32 plus.n31 5.84292
R60 plus.n8 plus.n7 0.189894
R61 plus.n8 plus.n2 0.189894
R62 plus.n13 plus.n2 0.189894
R63 plus.n14 plus.n13 0.189894
R64 plus.n14 plus.n0 0.189894
R65 plus.n20 plus.n0 0.189894
R66 plus.n41 plus.n21 0.189894
R67 plus.n35 plus.n21 0.189894
R68 plus.n35 plus.n34 0.189894
R69 plus.n34 plus.n23 0.189894
R70 plus.n29 plus.n23 0.189894
R71 plus.n29 plus.n28 0.189894
R72 source.n0 source.t30 44.1297
R73 source.n7 source.t27 44.1296
R74 source.n8 source.t15 44.1296
R75 source.n15 source.t13 44.1296
R76 source.n31 source.t5 44.1295
R77 source.n24 source.t1 44.1295
R78 source.n23 source.t20 44.1295
R79 source.n16 source.t31 44.1295
R80 source.n2 source.n1 43.1397
R81 source.n4 source.n3 43.1397
R82 source.n6 source.n5 43.1397
R83 source.n10 source.n9 43.1397
R84 source.n12 source.n11 43.1397
R85 source.n14 source.n13 43.1397
R86 source.n30 source.n29 43.1396
R87 source.n28 source.n27 43.1396
R88 source.n26 source.n25 43.1396
R89 source.n22 source.n21 43.1396
R90 source.n20 source.n19 43.1396
R91 source.n18 source.n17 43.1396
R92 source.n16 source.n15 27.8483
R93 source.n32 source.n0 22.3354
R94 source.n32 source.n31 5.51343
R95 source.n29 source.t3 0.9905
R96 source.n29 source.t11 0.9905
R97 source.n27 source.t4 0.9905
R98 source.n27 source.t12 0.9905
R99 source.n25 source.t7 0.9905
R100 source.n25 source.t14 0.9905
R101 source.n21 source.t26 0.9905
R102 source.n21 source.t29 0.9905
R103 source.n19 source.t19 0.9905
R104 source.n19 source.t28 0.9905
R105 source.n17 source.t21 0.9905
R106 source.n17 source.t22 0.9905
R107 source.n1 source.t18 0.9905
R108 source.n1 source.t23 0.9905
R109 source.n3 source.t16 0.9905
R110 source.n3 source.t24 0.9905
R111 source.n5 source.t25 0.9905
R112 source.n5 source.t17 0.9905
R113 source.n9 source.t6 0.9905
R114 source.n9 source.t10 0.9905
R115 source.n11 source.t0 0.9905
R116 source.n11 source.t8 0.9905
R117 source.n13 source.t2 0.9905
R118 source.n13 source.t9 0.9905
R119 source.n15 source.n14 0.5005
R120 source.n14 source.n12 0.5005
R121 source.n12 source.n10 0.5005
R122 source.n10 source.n8 0.5005
R123 source.n7 source.n6 0.5005
R124 source.n6 source.n4 0.5005
R125 source.n4 source.n2 0.5005
R126 source.n2 source.n0 0.5005
R127 source.n18 source.n16 0.5005
R128 source.n20 source.n18 0.5005
R129 source.n22 source.n20 0.5005
R130 source.n23 source.n22 0.5005
R131 source.n26 source.n24 0.5005
R132 source.n28 source.n26 0.5005
R133 source.n30 source.n28 0.5005
R134 source.n31 source.n30 0.5005
R135 source.n8 source.n7 0.470328
R136 source.n24 source.n23 0.470328
R137 source source.n32 0.188
R138 drain_left.n9 drain_left.n7 60.3185
R139 drain_left.n5 drain_left.n3 60.3184
R140 drain_left.n2 drain_left.n0 60.3184
R141 drain_left.n13 drain_left.n12 59.8185
R142 drain_left.n11 drain_left.n10 59.8185
R143 drain_left.n9 drain_left.n8 59.8185
R144 drain_left.n5 drain_left.n4 59.8184
R145 drain_left.n2 drain_left.n1 59.8184
R146 drain_left drain_left.n6 36.6777
R147 drain_left drain_left.n13 6.15322
R148 drain_left.n3 drain_left.t2 0.9905
R149 drain_left.n3 drain_left.t13 0.9905
R150 drain_left.n4 drain_left.t11 0.9905
R151 drain_left.n4 drain_left.t4 0.9905
R152 drain_left.n1 drain_left.t0 0.9905
R153 drain_left.n1 drain_left.t9 0.9905
R154 drain_left.n0 drain_left.t8 0.9905
R155 drain_left.n0 drain_left.t3 0.9905
R156 drain_left.n12 drain_left.t7 0.9905
R157 drain_left.n12 drain_left.t12 0.9905
R158 drain_left.n10 drain_left.t6 0.9905
R159 drain_left.n10 drain_left.t1 0.9905
R160 drain_left.n8 drain_left.t5 0.9905
R161 drain_left.n8 drain_left.t15 0.9905
R162 drain_left.n7 drain_left.t10 0.9905
R163 drain_left.n7 drain_left.t14 0.9905
R164 drain_left.n11 drain_left.n9 0.5005
R165 drain_left.n13 drain_left.n11 0.5005
R166 drain_left.n6 drain_left.n5 0.195154
R167 drain_left.n6 drain_left.n2 0.195154
R168 minus.n19 minus.t4 2094.22
R169 minus.n4 minus.t9 2094.22
R170 minus.n40 minus.t13 2094.22
R171 minus.n25 minus.t2 2094.22
R172 minus.n18 minus.t12 2053.32
R173 minus.n16 minus.t6 2053.32
R174 minus.n1 minus.t11 2053.32
R175 minus.n10 minus.t1 2053.32
R176 minus.n3 minus.t8 2053.32
R177 minus.n5 minus.t3 2053.32
R178 minus.n39 minus.t14 2053.32
R179 minus.n37 minus.t0 2053.32
R180 minus.n22 minus.t7 2053.32
R181 minus.n31 minus.t10 2053.32
R182 minus.n24 minus.t15 2053.32
R183 minus.n26 minus.t5 2053.32
R184 minus.n7 minus.n4 161.489
R185 minus.n28 minus.n25 161.489
R186 minus.n20 minus.n19 161.3
R187 minus.n17 minus.n0 161.3
R188 minus.n15 minus.n14 161.3
R189 minus.n13 minus.n12 161.3
R190 minus.n11 minus.n2 161.3
R191 minus.n9 minus.n8 161.3
R192 minus.n7 minus.n6 161.3
R193 minus.n41 minus.n40 161.3
R194 minus.n38 minus.n21 161.3
R195 minus.n36 minus.n35 161.3
R196 minus.n34 minus.n33 161.3
R197 minus.n32 minus.n23 161.3
R198 minus.n30 minus.n29 161.3
R199 minus.n28 minus.n27 161.3
R200 minus.n12 minus.n11 73.0308
R201 minus.n33 minus.n32 73.0308
R202 minus.n15 minus.n1 67.1884
R203 minus.n10 minus.n9 67.1884
R204 minus.n31 minus.n30 67.1884
R205 minus.n36 minus.n22 67.1884
R206 minus.n17 minus.n16 55.5035
R207 minus.n6 minus.n3 55.5035
R208 minus.n27 minus.n24 55.5035
R209 minus.n38 minus.n37 55.5035
R210 minus.n19 minus.n18 43.8187
R211 minus.n5 minus.n4 43.8187
R212 minus.n26 minus.n25 43.8187
R213 minus.n40 minus.n39 43.8187
R214 minus.n42 minus.n20 41.8149
R215 minus.n18 minus.n17 29.2126
R216 minus.n6 minus.n5 29.2126
R217 minus.n27 minus.n26 29.2126
R218 minus.n39 minus.n38 29.2126
R219 minus.n16 minus.n15 17.5278
R220 minus.n9 minus.n3 17.5278
R221 minus.n30 minus.n24 17.5278
R222 minus.n37 minus.n36 17.5278
R223 minus.n42 minus.n41 6.46641
R224 minus.n12 minus.n1 5.84292
R225 minus.n11 minus.n10 5.84292
R226 minus.n32 minus.n31 5.84292
R227 minus.n33 minus.n22 5.84292
R228 minus.n20 minus.n0 0.189894
R229 minus.n14 minus.n0 0.189894
R230 minus.n14 minus.n13 0.189894
R231 minus.n13 minus.n2 0.189894
R232 minus.n8 minus.n2 0.189894
R233 minus.n8 minus.n7 0.189894
R234 minus.n29 minus.n28 0.189894
R235 minus.n29 minus.n23 0.189894
R236 minus.n34 minus.n23 0.189894
R237 minus.n35 minus.n34 0.189894
R238 minus.n35 minus.n21 0.189894
R239 minus.n41 minus.n21 0.189894
R240 minus minus.n42 0.188
R241 drain_right.n9 drain_right.n7 60.3185
R242 drain_right.n5 drain_right.n3 60.3184
R243 drain_right.n2 drain_right.n0 60.3184
R244 drain_right.n9 drain_right.n8 59.8185
R245 drain_right.n11 drain_right.n10 59.8185
R246 drain_right.n13 drain_right.n12 59.8185
R247 drain_right.n5 drain_right.n4 59.8184
R248 drain_right.n2 drain_right.n1 59.8184
R249 drain_right drain_right.n6 36.1245
R250 drain_right drain_right.n13 6.15322
R251 drain_right.n3 drain_right.t1 0.9905
R252 drain_right.n3 drain_right.t2 0.9905
R253 drain_right.n4 drain_right.t8 0.9905
R254 drain_right.n4 drain_right.t15 0.9905
R255 drain_right.n1 drain_right.t0 0.9905
R256 drain_right.n1 drain_right.t5 0.9905
R257 drain_right.n0 drain_right.t13 0.9905
R258 drain_right.n0 drain_right.t10 0.9905
R259 drain_right.n7 drain_right.t12 0.9905
R260 drain_right.n7 drain_right.t6 0.9905
R261 drain_right.n8 drain_right.t14 0.9905
R262 drain_right.n8 drain_right.t7 0.9905
R263 drain_right.n10 drain_right.t9 0.9905
R264 drain_right.n10 drain_right.t4 0.9905
R265 drain_right.n12 drain_right.t11 0.9905
R266 drain_right.n12 drain_right.t3 0.9905
R267 drain_right.n13 drain_right.n11 0.5005
R268 drain_right.n11 drain_right.n9 0.5005
R269 drain_right.n6 drain_right.n5 0.195154
R270 drain_right.n6 drain_right.n2 0.195154
C0 drain_left source 53.5622f
C1 source plus 7.61285f
C2 drain_left plus 8.47253f
C3 source drain_right 53.5622f
C4 source minus 7.59881f
C5 drain_left drain_right 0.897273f
C6 plus drain_right 0.324551f
C7 drain_left minus 0.171252f
C8 minus plus 6.83165f
C9 minus drain_right 8.30219f
C10 drain_right a_n1760_n4888# 8.43007f
C11 drain_left a_n1760_n4888# 8.71083f
C12 source a_n1760_n4888# 12.93929f
C13 minus a_n1760_n4888# 7.389741f
C14 plus a_n1760_n4888# 9.953871f
C15 drain_right.t13 a_n1760_n4888# 0.574773f
C16 drain_right.t10 a_n1760_n4888# 0.574773f
C17 drain_right.n0 a_n1760_n4888# 5.25834f
C18 drain_right.t0 a_n1760_n4888# 0.574773f
C19 drain_right.t5 a_n1760_n4888# 0.574773f
C20 drain_right.n1 a_n1760_n4888# 5.2547f
C21 drain_right.n2 a_n1760_n4888# 0.827707f
C22 drain_right.t1 a_n1760_n4888# 0.574773f
C23 drain_right.t2 a_n1760_n4888# 0.574773f
C24 drain_right.n3 a_n1760_n4888# 5.25834f
C25 drain_right.t8 a_n1760_n4888# 0.574773f
C26 drain_right.t15 a_n1760_n4888# 0.574773f
C27 drain_right.n4 a_n1760_n4888# 5.2547f
C28 drain_right.n5 a_n1760_n4888# 0.827707f
C29 drain_right.n6 a_n1760_n4888# 2.38283f
C30 drain_right.t12 a_n1760_n4888# 0.574773f
C31 drain_right.t6 a_n1760_n4888# 0.574773f
C32 drain_right.n7 a_n1760_n4888# 5.25833f
C33 drain_right.t14 a_n1760_n4888# 0.574773f
C34 drain_right.t7 a_n1760_n4888# 0.574773f
C35 drain_right.n8 a_n1760_n4888# 5.2547f
C36 drain_right.n9 a_n1760_n4888# 0.859172f
C37 drain_right.t9 a_n1760_n4888# 0.574773f
C38 drain_right.t4 a_n1760_n4888# 0.574773f
C39 drain_right.n10 a_n1760_n4888# 5.2547f
C40 drain_right.n11 a_n1760_n4888# 0.424081f
C41 drain_right.t11 a_n1760_n4888# 0.574773f
C42 drain_right.t3 a_n1760_n4888# 0.574773f
C43 drain_right.n12 a_n1760_n4888# 5.2547f
C44 drain_right.n13 a_n1760_n4888# 0.724269f
C45 minus.n0 a_n1760_n4888# 0.05231f
C46 minus.t4 a_n1760_n4888# 0.742069f
C47 minus.t12 a_n1760_n4888# 0.736654f
C48 minus.t6 a_n1760_n4888# 0.736654f
C49 minus.t11 a_n1760_n4888# 0.736654f
C50 minus.n1 a_n1760_n4888# 0.276337f
C51 minus.n2 a_n1760_n4888# 0.05231f
C52 minus.t1 a_n1760_n4888# 0.736654f
C53 minus.t8 a_n1760_n4888# 0.736654f
C54 minus.n3 a_n1760_n4888# 0.276337f
C55 minus.t9 a_n1760_n4888# 0.742069f
C56 minus.n4 a_n1760_n4888# 0.291895f
C57 minus.t3 a_n1760_n4888# 0.736654f
C58 minus.n5 a_n1760_n4888# 0.276337f
C59 minus.n6 a_n1760_n4888# 0.019933f
C60 minus.n7 a_n1760_n4888# 0.114545f
C61 minus.n8 a_n1760_n4888# 0.05231f
C62 minus.n9 a_n1760_n4888# 0.019933f
C63 minus.n10 a_n1760_n4888# 0.276337f
C64 minus.n11 a_n1760_n4888# 0.018643f
C65 minus.n12 a_n1760_n4888# 0.018643f
C66 minus.n13 a_n1760_n4888# 0.05231f
C67 minus.n14 a_n1760_n4888# 0.05231f
C68 minus.n15 a_n1760_n4888# 0.019933f
C69 minus.n16 a_n1760_n4888# 0.276337f
C70 minus.n17 a_n1760_n4888# 0.019933f
C71 minus.n18 a_n1760_n4888# 0.276337f
C72 minus.n19 a_n1760_n4888# 0.291822f
C73 minus.n20 a_n1760_n4888# 2.30043f
C74 minus.n21 a_n1760_n4888# 0.05231f
C75 minus.t14 a_n1760_n4888# 0.736654f
C76 minus.t0 a_n1760_n4888# 0.736654f
C77 minus.t7 a_n1760_n4888# 0.736654f
C78 minus.n22 a_n1760_n4888# 0.276337f
C79 minus.n23 a_n1760_n4888# 0.05231f
C80 minus.t10 a_n1760_n4888# 0.736654f
C81 minus.t15 a_n1760_n4888# 0.736654f
C82 minus.n24 a_n1760_n4888# 0.276337f
C83 minus.t2 a_n1760_n4888# 0.742069f
C84 minus.n25 a_n1760_n4888# 0.291895f
C85 minus.t5 a_n1760_n4888# 0.736654f
C86 minus.n26 a_n1760_n4888# 0.276337f
C87 minus.n27 a_n1760_n4888# 0.019933f
C88 minus.n28 a_n1760_n4888# 0.114545f
C89 minus.n29 a_n1760_n4888# 0.05231f
C90 minus.n30 a_n1760_n4888# 0.019933f
C91 minus.n31 a_n1760_n4888# 0.276337f
C92 minus.n32 a_n1760_n4888# 0.018643f
C93 minus.n33 a_n1760_n4888# 0.018643f
C94 minus.n34 a_n1760_n4888# 0.05231f
C95 minus.n35 a_n1760_n4888# 0.05231f
C96 minus.n36 a_n1760_n4888# 0.019933f
C97 minus.n37 a_n1760_n4888# 0.276337f
C98 minus.n38 a_n1760_n4888# 0.019933f
C99 minus.n39 a_n1760_n4888# 0.276337f
C100 minus.t13 a_n1760_n4888# 0.742069f
C101 minus.n40 a_n1760_n4888# 0.291822f
C102 minus.n41 a_n1760_n4888# 0.337845f
C103 minus.n42 a_n1760_n4888# 2.74954f
C104 drain_left.t8 a_n1760_n4888# 0.575308f
C105 drain_left.t3 a_n1760_n4888# 0.575308f
C106 drain_left.n0 a_n1760_n4888# 5.26323f
C107 drain_left.t0 a_n1760_n4888# 0.575308f
C108 drain_left.t9 a_n1760_n4888# 0.575308f
C109 drain_left.n1 a_n1760_n4888# 5.25959f
C110 drain_left.n2 a_n1760_n4888# 0.828478f
C111 drain_left.t2 a_n1760_n4888# 0.575308f
C112 drain_left.t13 a_n1760_n4888# 0.575308f
C113 drain_left.n3 a_n1760_n4888# 5.26323f
C114 drain_left.t11 a_n1760_n4888# 0.575308f
C115 drain_left.t4 a_n1760_n4888# 0.575308f
C116 drain_left.n4 a_n1760_n4888# 5.25959f
C117 drain_left.n5 a_n1760_n4888# 0.828477f
C118 drain_left.n6 a_n1760_n4888# 2.4609f
C119 drain_left.t10 a_n1760_n4888# 0.575308f
C120 drain_left.t14 a_n1760_n4888# 0.575308f
C121 drain_left.n7 a_n1760_n4888# 5.26323f
C122 drain_left.t5 a_n1760_n4888# 0.575308f
C123 drain_left.t15 a_n1760_n4888# 0.575308f
C124 drain_left.n8 a_n1760_n4888# 5.25959f
C125 drain_left.n9 a_n1760_n4888# 0.859972f
C126 drain_left.t6 a_n1760_n4888# 0.575308f
C127 drain_left.t1 a_n1760_n4888# 0.575308f
C128 drain_left.n10 a_n1760_n4888# 5.25959f
C129 drain_left.n11 a_n1760_n4888# 0.424475f
C130 drain_left.t7 a_n1760_n4888# 0.575308f
C131 drain_left.t12 a_n1760_n4888# 0.575308f
C132 drain_left.n12 a_n1760_n4888# 5.25959f
C133 drain_left.n13 a_n1760_n4888# 0.724943f
C134 source.t30 a_n1760_n4888# 5.35311f
C135 source.n0 a_n1760_n4888# 2.27037f
C136 source.t18 a_n1760_n4888# 0.468405f
C137 source.t23 a_n1760_n4888# 0.468405f
C138 source.n1 a_n1760_n4888# 4.18774f
C139 source.n2 a_n1760_n4888# 0.399831f
C140 source.t16 a_n1760_n4888# 0.468405f
C141 source.t24 a_n1760_n4888# 0.468405f
C142 source.n3 a_n1760_n4888# 4.18774f
C143 source.n4 a_n1760_n4888# 0.399831f
C144 source.t25 a_n1760_n4888# 0.468405f
C145 source.t17 a_n1760_n4888# 0.468405f
C146 source.n5 a_n1760_n4888# 4.18774f
C147 source.n6 a_n1760_n4888# 0.399831f
C148 source.t27 a_n1760_n4888# 5.35312f
C149 source.n7 a_n1760_n4888# 0.509037f
C150 source.t15 a_n1760_n4888# 5.35312f
C151 source.n8 a_n1760_n4888# 0.509037f
C152 source.t6 a_n1760_n4888# 0.468405f
C153 source.t10 a_n1760_n4888# 0.468405f
C154 source.n9 a_n1760_n4888# 4.18774f
C155 source.n10 a_n1760_n4888# 0.399831f
C156 source.t0 a_n1760_n4888# 0.468405f
C157 source.t8 a_n1760_n4888# 0.468405f
C158 source.n11 a_n1760_n4888# 4.18774f
C159 source.n12 a_n1760_n4888# 0.399831f
C160 source.t2 a_n1760_n4888# 0.468405f
C161 source.t9 a_n1760_n4888# 0.468405f
C162 source.n13 a_n1760_n4888# 4.18774f
C163 source.n14 a_n1760_n4888# 0.399831f
C164 source.t13 a_n1760_n4888# 5.35312f
C165 source.n15 a_n1760_n4888# 2.79383f
C166 source.t31 a_n1760_n4888# 5.35309f
C167 source.n16 a_n1760_n4888# 2.79386f
C168 source.t21 a_n1760_n4888# 0.468405f
C169 source.t22 a_n1760_n4888# 0.468405f
C170 source.n17 a_n1760_n4888# 4.18775f
C171 source.n18 a_n1760_n4888# 0.399823f
C172 source.t19 a_n1760_n4888# 0.468405f
C173 source.t28 a_n1760_n4888# 0.468405f
C174 source.n19 a_n1760_n4888# 4.18775f
C175 source.n20 a_n1760_n4888# 0.399823f
C176 source.t26 a_n1760_n4888# 0.468405f
C177 source.t29 a_n1760_n4888# 0.468405f
C178 source.n21 a_n1760_n4888# 4.18775f
C179 source.n22 a_n1760_n4888# 0.399823f
C180 source.t20 a_n1760_n4888# 5.35309f
C181 source.n23 a_n1760_n4888# 0.509067f
C182 source.t1 a_n1760_n4888# 5.35309f
C183 source.n24 a_n1760_n4888# 0.509067f
C184 source.t7 a_n1760_n4888# 0.468405f
C185 source.t14 a_n1760_n4888# 0.468405f
C186 source.n25 a_n1760_n4888# 4.18775f
C187 source.n26 a_n1760_n4888# 0.399823f
C188 source.t4 a_n1760_n4888# 0.468405f
C189 source.t12 a_n1760_n4888# 0.468405f
C190 source.n27 a_n1760_n4888# 4.18775f
C191 source.n28 a_n1760_n4888# 0.399823f
C192 source.t3 a_n1760_n4888# 0.468405f
C193 source.t11 a_n1760_n4888# 0.468405f
C194 source.n29 a_n1760_n4888# 4.18775f
C195 source.n30 a_n1760_n4888# 0.399823f
C196 source.t5 a_n1760_n4888# 5.35309f
C197 source.n31 a_n1760_n4888# 0.673074f
C198 source.n32 a_n1760_n4888# 2.66534f
C199 plus.n0 a_n1760_n4888# 0.053018f
C200 plus.t8 a_n1760_n4888# 0.746624f
C201 plus.t14 a_n1760_n4888# 0.746624f
C202 plus.t9 a_n1760_n4888# 0.746624f
C203 plus.n1 a_n1760_n4888# 0.280077f
C204 plus.n2 a_n1760_n4888# 0.053018f
C205 plus.t0 a_n1760_n4888# 0.746624f
C206 plus.t10 a_n1760_n4888# 0.746624f
C207 plus.n3 a_n1760_n4888# 0.280077f
C208 plus.t5 a_n1760_n4888# 0.752112f
C209 plus.n4 a_n1760_n4888# 0.295846f
C210 plus.t1 a_n1760_n4888# 0.746624f
C211 plus.n5 a_n1760_n4888# 0.280077f
C212 plus.n6 a_n1760_n4888# 0.020203f
C213 plus.n7 a_n1760_n4888# 0.116096f
C214 plus.n8 a_n1760_n4888# 0.053018f
C215 plus.n9 a_n1760_n4888# 0.020203f
C216 plus.n10 a_n1760_n4888# 0.280077f
C217 plus.n11 a_n1760_n4888# 0.018895f
C218 plus.n12 a_n1760_n4888# 0.018895f
C219 plus.n13 a_n1760_n4888# 0.053018f
C220 plus.n14 a_n1760_n4888# 0.053018f
C221 plus.n15 a_n1760_n4888# 0.020203f
C222 plus.n16 a_n1760_n4888# 0.280077f
C223 plus.n17 a_n1760_n4888# 0.020203f
C224 plus.n18 a_n1760_n4888# 0.280077f
C225 plus.t3 a_n1760_n4888# 0.752112f
C226 plus.n19 a_n1760_n4888# 0.295772f
C227 plus.n20 a_n1760_n4888# 0.800946f
C228 plus.n21 a_n1760_n4888# 0.053018f
C229 plus.t7 a_n1760_n4888# 0.752112f
C230 plus.t12 a_n1760_n4888# 0.746624f
C231 plus.t15 a_n1760_n4888# 0.746624f
C232 plus.t6 a_n1760_n4888# 0.746624f
C233 plus.n22 a_n1760_n4888# 0.280077f
C234 plus.n23 a_n1760_n4888# 0.053018f
C235 plus.t4 a_n1760_n4888# 0.746624f
C236 plus.t11 a_n1760_n4888# 0.746624f
C237 plus.n24 a_n1760_n4888# 0.280077f
C238 plus.t2 a_n1760_n4888# 0.752112f
C239 plus.n25 a_n1760_n4888# 0.295846f
C240 plus.t13 a_n1760_n4888# 0.746624f
C241 plus.n26 a_n1760_n4888# 0.280077f
C242 plus.n27 a_n1760_n4888# 0.020203f
C243 plus.n28 a_n1760_n4888# 0.116096f
C244 plus.n29 a_n1760_n4888# 0.053018f
C245 plus.n30 a_n1760_n4888# 0.020203f
C246 plus.n31 a_n1760_n4888# 0.280077f
C247 plus.n32 a_n1760_n4888# 0.018895f
C248 plus.n33 a_n1760_n4888# 0.018895f
C249 plus.n34 a_n1760_n4888# 0.053018f
C250 plus.n35 a_n1760_n4888# 0.053018f
C251 plus.n36 a_n1760_n4888# 0.020203f
C252 plus.n37 a_n1760_n4888# 0.280077f
C253 plus.n38 a_n1760_n4888# 0.020203f
C254 plus.n39 a_n1760_n4888# 0.280077f
C255 plus.n40 a_n1760_n4888# 0.295772f
C256 plus.n41 a_n1760_n4888# 1.84103f
.ends

