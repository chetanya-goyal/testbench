* NGSPICE file created from diffpair352.ext - technology: sky130A

.subckt diffpair352 minus drain_right drain_left source plus
X0 drain_right.t5 minus.t0 source.t7 a_n1220_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X1 a_n1220_n2688# a_n1220_n2688# a_n1220_n2688# a_n1220_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.3
X2 drain_left.t5 plus.t0 source.t1 a_n1220_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X3 source.t2 plus.t1 drain_left.t4 a_n1220_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X4 a_n1220_n2688# a_n1220_n2688# a_n1220_n2688# a_n1220_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X5 a_n1220_n2688# a_n1220_n2688# a_n1220_n2688# a_n1220_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X6 source.t0 plus.t2 drain_left.t3 a_n1220_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X7 source.t8 minus.t1 drain_right.t4 a_n1220_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X8 a_n1220_n2688# a_n1220_n2688# a_n1220_n2688# a_n1220_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X9 drain_right.t3 minus.t2 source.t6 a_n1220_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X10 drain_left.t2 plus.t3 source.t5 a_n1220_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X11 drain_left.t1 plus.t4 source.t4 a_n1220_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X12 drain_left.t0 plus.t5 source.t3 a_n1220_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X13 source.t9 minus.t3 drain_right.t2 a_n1220_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X14 drain_right.t1 minus.t4 source.t10 a_n1220_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X15 drain_right.t0 minus.t5 source.t11 a_n1220_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
R0 minus.n2 minus.t0 882.937
R1 minus.n0 minus.t2 882.937
R2 minus.n6 minus.t4 882.937
R3 minus.n4 minus.t5 882.937
R4 minus.n1 minus.t3 827.433
R5 minus.n5 minus.t1 827.433
R6 minus.n3 minus.n0 161.489
R7 minus.n7 minus.n4 161.489
R8 minus.n3 minus.n2 161.3
R9 minus.n7 minus.n6 161.3
R10 minus.n2 minus.n1 36.5157
R11 minus.n1 minus.n0 36.5157
R12 minus.n5 minus.n4 36.5157
R13 minus.n6 minus.n5 36.5157
R14 minus.n8 minus.n3 31.5024
R15 minus.n8 minus.n7 6.5327
R16 minus minus.n8 0.188
R17 source.n3 source.t6 51.0588
R18 source.n11 source.t10 51.0586
R19 source.n8 source.t5 51.0586
R20 source.n0 source.t4 51.0586
R21 source.n2 source.n1 48.8588
R22 source.n5 source.n4 48.8588
R23 source.n10 source.n9 48.8586
R24 source.n7 source.n6 48.8586
R25 source.n7 source.n5 20.1012
R26 source.n12 source.n0 14.0236
R27 source.n12 source.n11 5.53498
R28 source.n9 source.t11 2.2005
R29 source.n9 source.t8 2.2005
R30 source.n6 source.t3 2.2005
R31 source.n6 source.t2 2.2005
R32 source.n1 source.t1 2.2005
R33 source.n1 source.t0 2.2005
R34 source.n4 source.t7 2.2005
R35 source.n4 source.t9 2.2005
R36 source.n3 source.n2 0.741879
R37 source.n10 source.n8 0.741879
R38 source.n5 source.n3 0.543603
R39 source.n2 source.n0 0.543603
R40 source.n8 source.n7 0.543603
R41 source.n11 source.n10 0.543603
R42 source source.n12 0.188
R43 drain_right.n1 drain_right.t0 68.0893
R44 drain_right.n3 drain_right.t5 67.7376
R45 drain_right.n3 drain_right.n2 66.0805
R46 drain_right.n1 drain_right.n0 65.6178
R47 drain_right drain_right.n1 26.0347
R48 drain_right drain_right.n3 5.92477
R49 drain_right.n0 drain_right.t4 2.2005
R50 drain_right.n0 drain_right.t1 2.2005
R51 drain_right.n2 drain_right.t2 2.2005
R52 drain_right.n2 drain_right.t3 2.2005
R53 plus.n0 plus.t0 882.937
R54 plus.n2 plus.t4 882.937
R55 plus.n4 plus.t3 882.937
R56 plus.n6 plus.t5 882.937
R57 plus.n1 plus.t2 827.433
R58 plus.n5 plus.t1 827.433
R59 plus.n3 plus.n0 161.489
R60 plus.n7 plus.n4 161.489
R61 plus.n3 plus.n2 161.3
R62 plus.n7 plus.n6 161.3
R63 plus.n1 plus.n0 36.5157
R64 plus.n2 plus.n1 36.5157
R65 plus.n6 plus.n5 36.5157
R66 plus.n5 plus.n4 36.5157
R67 plus plus.n7 26.5199
R68 plus plus.n3 11.0403
R69 drain_left.n3 drain_left.t5 68.2807
R70 drain_left.n1 drain_left.t0 68.0893
R71 drain_left.n1 drain_left.n0 65.6178
R72 drain_left.n3 drain_left.n2 65.5374
R73 drain_left drain_left.n1 26.5879
R74 drain_left drain_left.n3 6.19632
R75 drain_left.n0 drain_left.t4 2.2005
R76 drain_left.n0 drain_left.t2 2.2005
R77 drain_left.n2 drain_left.t3 2.2005
R78 drain_left.n2 drain_left.t1 2.2005
C0 drain_left source 10.975901f
C1 drain_right plus 0.26923f
C2 minus drain_left 0.17071f
C3 source plus 1.79966f
C4 minus plus 4.11274f
C5 source drain_right 10.9667f
C6 minus drain_right 2.1247f
C7 minus source 1.78514f
C8 drain_left plus 2.23673f
C9 drain_left drain_right 0.56775f
C10 drain_right a_n1220_n2688# 5.45674f
C11 drain_left a_n1220_n2688# 5.643099f
C12 source a_n1220_n2688# 4.984919f
C13 minus a_n1220_n2688# 4.44913f
C14 plus a_n1220_n2688# 5.828361f
C15 drain_left.t0 a_n1220_n2688# 2.17114f
C16 drain_left.t4 a_n1220_n2688# 0.194852f
C17 drain_left.t2 a_n1220_n2688# 0.194852f
C18 drain_left.n0 a_n1220_n2688# 1.70466f
C19 drain_left.n1 a_n1220_n2688# 1.59701f
C20 drain_left.t5 a_n1220_n2688# 2.17218f
C21 drain_left.t3 a_n1220_n2688# 0.194852f
C22 drain_left.t1 a_n1220_n2688# 0.194852f
C23 drain_left.n2 a_n1220_n2688# 1.7043f
C24 drain_left.n3 a_n1220_n2688# 0.88537f
C25 plus.t0 a_n1220_n2688# 0.358416f
C26 plus.n0 a_n1220_n2688# 0.160152f
C27 plus.t2 a_n1220_n2688# 0.348939f
C28 plus.n1 a_n1220_n2688# 0.145711f
C29 plus.t4 a_n1220_n2688# 0.358416f
C30 plus.n2 a_n1220_n2688# 0.16008f
C31 plus.n3 a_n1220_n2688# 0.512909f
C32 plus.t3 a_n1220_n2688# 0.358416f
C33 plus.n4 a_n1220_n2688# 0.160152f
C34 plus.t5 a_n1220_n2688# 0.358416f
C35 plus.t1 a_n1220_n2688# 0.348939f
C36 plus.n5 a_n1220_n2688# 0.145711f
C37 plus.n6 a_n1220_n2688# 0.16008f
C38 plus.n7 a_n1220_n2688# 1.18475f
C39 drain_right.t0 a_n1220_n2688# 2.17233f
C40 drain_right.t4 a_n1220_n2688# 0.194959f
C41 drain_right.t1 a_n1220_n2688# 0.194959f
C42 drain_right.n0 a_n1220_n2688# 1.7056f
C43 drain_right.n1 a_n1220_n2688# 1.54078f
C44 drain_right.t2 a_n1220_n2688# 0.194959f
C45 drain_right.t3 a_n1220_n2688# 0.194959f
C46 drain_right.n2 a_n1220_n2688# 1.70792f
C47 drain_right.t5 a_n1220_n2688# 2.17063f
C48 drain_right.n3 a_n1220_n2688# 0.897473f
C49 source.t4 a_n1220_n2688# 1.87322f
C50 source.n0 a_n1220_n2688# 1.07715f
C51 source.t1 a_n1220_n2688# 0.175667f
C52 source.t0 a_n1220_n2688# 0.175667f
C53 source.n1 a_n1220_n2688# 1.47057f
C54 source.n2 a_n1220_n2688# 0.332437f
C55 source.t6 a_n1220_n2688# 1.87322f
C56 source.n3 a_n1220_n2688# 0.408875f
C57 source.t7 a_n1220_n2688# 0.175667f
C58 source.t9 a_n1220_n2688# 0.175667f
C59 source.n4 a_n1220_n2688# 1.47057f
C60 source.n5 a_n1220_n2688# 1.40282f
C61 source.t3 a_n1220_n2688# 0.175667f
C62 source.t2 a_n1220_n2688# 0.175667f
C63 source.n6 a_n1220_n2688# 1.47057f
C64 source.n7 a_n1220_n2688# 1.40283f
C65 source.t5 a_n1220_n2688# 1.87322f
C66 source.n8 a_n1220_n2688# 0.408879f
C67 source.t11 a_n1220_n2688# 0.175667f
C68 source.t8 a_n1220_n2688# 0.175667f
C69 source.n9 a_n1220_n2688# 1.47057f
C70 source.n10 a_n1220_n2688# 0.332441f
C71 source.t10 a_n1220_n2688# 1.87322f
C72 source.n11 a_n1220_n2688# 0.526697f
C73 source.n12 a_n1220_n2688# 1.2858f
C74 minus.t2 a_n1220_n2688# 0.347638f
C75 minus.n0 a_n1220_n2688# 0.155336f
C76 minus.t0 a_n1220_n2688# 0.347638f
C77 minus.t3 a_n1220_n2688# 0.338445f
C78 minus.n1 a_n1220_n2688# 0.141329f
C79 minus.n2 a_n1220_n2688# 0.155266f
C80 minus.n3 a_n1220_n2688# 1.31039f
C81 minus.t5 a_n1220_n2688# 0.347638f
C82 minus.n4 a_n1220_n2688# 0.155336f
C83 minus.t1 a_n1220_n2688# 0.338445f
C84 minus.n5 a_n1220_n2688# 0.141329f
C85 minus.t4 a_n1220_n2688# 0.347638f
C86 minus.n6 a_n1220_n2688# 0.155266f
C87 minus.n7 a_n1220_n2688# 0.352052f
C88 minus.n8 a_n1220_n2688# 1.53721f
.ends

