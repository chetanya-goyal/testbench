* NGSPICE file created from diffpair455.ext - technology: sky130A

.subckt diffpair455 minus drain_right drain_left source plus
X0 drain_right.t11 minus.t0 source.t17 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.6
X1 drain_left.t11 plus.t0 source.t4 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X2 source.t13 minus.t1 drain_right.t10 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X3 drain_right.t9 minus.t2 source.t10 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X4 source.t6 plus.t1 drain_left.t10 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.6
X5 drain_left.t9 plus.t2 source.t2 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.6
X6 drain_right.t8 minus.t3 source.t19 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X7 source.t11 minus.t4 drain_right.t7 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.6
X8 source.t15 minus.t5 drain_right.t6 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X9 source.t20 plus.t3 drain_left.t8 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X10 a_n2018_n3288# a_n2018_n3288# a_n2018_n3288# a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.6
X11 source.t21 plus.t4 drain_left.t7 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X12 source.t16 minus.t6 drain_right.t5 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X13 drain_right.t4 minus.t7 source.t14 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X14 source.t12 minus.t8 drain_right.t3 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.6
X15 a_n2018_n3288# a_n2018_n3288# a_n2018_n3288# a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.6
X16 drain_left.t6 plus.t5 source.t22 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X17 source.t18 minus.t9 drain_right.t2 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X18 source.t23 plus.t6 drain_left.t5 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X19 drain_right.t1 minus.t10 source.t8 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.6
X20 drain_left.t4 plus.t7 source.t1 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X21 a_n2018_n3288# a_n2018_n3288# a_n2018_n3288# a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.6
X22 drain_left.t3 plus.t8 source.t0 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X23 source.t3 plus.t9 drain_left.t2 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.6
X24 a_n2018_n3288# a_n2018_n3288# a_n2018_n3288# a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.6
X25 drain_right.t0 minus.t11 source.t9 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
X26 drain_left.t1 plus.t10 source.t5 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.6
X27 source.t7 plus.t11 drain_left.t0 a_n2018_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.6
R0 minus.n2 minus.t10 572.532
R1 minus.n14 minus.t8 572.532
R2 minus.n3 minus.t9 547.472
R3 minus.n4 minus.t7 547.472
R4 minus.n1 minus.t6 547.472
R5 minus.n8 minus.t3 547.472
R6 minus.n10 minus.t4 547.472
R7 minus.n15 minus.t2 547.472
R8 minus.n16 minus.t5 547.472
R9 minus.n13 minus.t11 547.472
R10 minus.n20 minus.t1 547.472
R11 minus.n22 minus.t0 547.472
R12 minus.n11 minus.n10 161.3
R13 minus.n9 minus.n0 161.3
R14 minus.n8 minus.n7 161.3
R15 minus.n23 minus.n22 161.3
R16 minus.n21 minus.n12 161.3
R17 minus.n20 minus.n19 161.3
R18 minus.n6 minus.n1 80.6037
R19 minus.n5 minus.n4 80.6037
R20 minus.n18 minus.n13 80.6037
R21 minus.n17 minus.n16 80.6037
R22 minus.n4 minus.n3 48.2005
R23 minus.n4 minus.n1 48.2005
R24 minus.n8 minus.n1 48.2005
R25 minus.n16 minus.n15 48.2005
R26 minus.n16 minus.n13 48.2005
R27 minus.n20 minus.n13 48.2005
R28 minus.n5 minus.n2 45.0744
R29 minus.n17 minus.n14 45.0744
R30 minus.n10 minus.n9 40.1672
R31 minus.n22 minus.n21 40.1672
R32 minus.n24 minus.n11 36.8528
R33 minus.n3 minus.n2 16.1124
R34 minus.n15 minus.n14 16.1124
R35 minus.n9 minus.n8 8.03383
R36 minus.n21 minus.n20 8.03383
R37 minus.n24 minus.n23 6.58762
R38 minus.n6 minus.n5 0.380177
R39 minus.n18 minus.n17 0.380177
R40 minus.n7 minus.n6 0.285035
R41 minus.n19 minus.n18 0.285035
R42 minus.n11 minus.n0 0.189894
R43 minus.n7 minus.n0 0.189894
R44 minus.n19 minus.n12 0.189894
R45 minus.n23 minus.n12 0.189894
R46 minus minus.n24 0.188
R47 source.n538 source.n478 289.615
R48 source.n468 source.n408 289.615
R49 source.n402 source.n342 289.615
R50 source.n332 source.n272 289.615
R51 source.n60 source.n0 289.615
R52 source.n130 source.n70 289.615
R53 source.n196 source.n136 289.615
R54 source.n266 source.n206 289.615
R55 source.n498 source.n497 185
R56 source.n503 source.n502 185
R57 source.n505 source.n504 185
R58 source.n494 source.n493 185
R59 source.n511 source.n510 185
R60 source.n513 source.n512 185
R61 source.n490 source.n489 185
R62 source.n520 source.n519 185
R63 source.n521 source.n488 185
R64 source.n523 source.n522 185
R65 source.n486 source.n485 185
R66 source.n529 source.n528 185
R67 source.n531 source.n530 185
R68 source.n482 source.n481 185
R69 source.n537 source.n536 185
R70 source.n539 source.n538 185
R71 source.n428 source.n427 185
R72 source.n433 source.n432 185
R73 source.n435 source.n434 185
R74 source.n424 source.n423 185
R75 source.n441 source.n440 185
R76 source.n443 source.n442 185
R77 source.n420 source.n419 185
R78 source.n450 source.n449 185
R79 source.n451 source.n418 185
R80 source.n453 source.n452 185
R81 source.n416 source.n415 185
R82 source.n459 source.n458 185
R83 source.n461 source.n460 185
R84 source.n412 source.n411 185
R85 source.n467 source.n466 185
R86 source.n469 source.n468 185
R87 source.n362 source.n361 185
R88 source.n367 source.n366 185
R89 source.n369 source.n368 185
R90 source.n358 source.n357 185
R91 source.n375 source.n374 185
R92 source.n377 source.n376 185
R93 source.n354 source.n353 185
R94 source.n384 source.n383 185
R95 source.n385 source.n352 185
R96 source.n387 source.n386 185
R97 source.n350 source.n349 185
R98 source.n393 source.n392 185
R99 source.n395 source.n394 185
R100 source.n346 source.n345 185
R101 source.n401 source.n400 185
R102 source.n403 source.n402 185
R103 source.n292 source.n291 185
R104 source.n297 source.n296 185
R105 source.n299 source.n298 185
R106 source.n288 source.n287 185
R107 source.n305 source.n304 185
R108 source.n307 source.n306 185
R109 source.n284 source.n283 185
R110 source.n314 source.n313 185
R111 source.n315 source.n282 185
R112 source.n317 source.n316 185
R113 source.n280 source.n279 185
R114 source.n323 source.n322 185
R115 source.n325 source.n324 185
R116 source.n276 source.n275 185
R117 source.n331 source.n330 185
R118 source.n333 source.n332 185
R119 source.n61 source.n60 185
R120 source.n59 source.n58 185
R121 source.n4 source.n3 185
R122 source.n53 source.n52 185
R123 source.n51 source.n50 185
R124 source.n8 source.n7 185
R125 source.n45 source.n44 185
R126 source.n43 source.n10 185
R127 source.n42 source.n41 185
R128 source.n13 source.n11 185
R129 source.n36 source.n35 185
R130 source.n34 source.n33 185
R131 source.n17 source.n16 185
R132 source.n28 source.n27 185
R133 source.n26 source.n25 185
R134 source.n21 source.n20 185
R135 source.n131 source.n130 185
R136 source.n129 source.n128 185
R137 source.n74 source.n73 185
R138 source.n123 source.n122 185
R139 source.n121 source.n120 185
R140 source.n78 source.n77 185
R141 source.n115 source.n114 185
R142 source.n113 source.n80 185
R143 source.n112 source.n111 185
R144 source.n83 source.n81 185
R145 source.n106 source.n105 185
R146 source.n104 source.n103 185
R147 source.n87 source.n86 185
R148 source.n98 source.n97 185
R149 source.n96 source.n95 185
R150 source.n91 source.n90 185
R151 source.n197 source.n196 185
R152 source.n195 source.n194 185
R153 source.n140 source.n139 185
R154 source.n189 source.n188 185
R155 source.n187 source.n186 185
R156 source.n144 source.n143 185
R157 source.n181 source.n180 185
R158 source.n179 source.n146 185
R159 source.n178 source.n177 185
R160 source.n149 source.n147 185
R161 source.n172 source.n171 185
R162 source.n170 source.n169 185
R163 source.n153 source.n152 185
R164 source.n164 source.n163 185
R165 source.n162 source.n161 185
R166 source.n157 source.n156 185
R167 source.n267 source.n266 185
R168 source.n265 source.n264 185
R169 source.n210 source.n209 185
R170 source.n259 source.n258 185
R171 source.n257 source.n256 185
R172 source.n214 source.n213 185
R173 source.n251 source.n250 185
R174 source.n249 source.n216 185
R175 source.n248 source.n247 185
R176 source.n219 source.n217 185
R177 source.n242 source.n241 185
R178 source.n240 source.n239 185
R179 source.n223 source.n222 185
R180 source.n234 source.n233 185
R181 source.n232 source.n231 185
R182 source.n227 source.n226 185
R183 source.n499 source.t17 149.524
R184 source.n429 source.t12 149.524
R185 source.n363 source.t5 149.524
R186 source.n293 source.t6 149.524
R187 source.n22 source.t2 149.524
R188 source.n92 source.t3 149.524
R189 source.n158 source.t8 149.524
R190 source.n228 source.t11 149.524
R191 source.n503 source.n497 104.615
R192 source.n504 source.n503 104.615
R193 source.n504 source.n493 104.615
R194 source.n511 source.n493 104.615
R195 source.n512 source.n511 104.615
R196 source.n512 source.n489 104.615
R197 source.n520 source.n489 104.615
R198 source.n521 source.n520 104.615
R199 source.n522 source.n521 104.615
R200 source.n522 source.n485 104.615
R201 source.n529 source.n485 104.615
R202 source.n530 source.n529 104.615
R203 source.n530 source.n481 104.615
R204 source.n537 source.n481 104.615
R205 source.n538 source.n537 104.615
R206 source.n433 source.n427 104.615
R207 source.n434 source.n433 104.615
R208 source.n434 source.n423 104.615
R209 source.n441 source.n423 104.615
R210 source.n442 source.n441 104.615
R211 source.n442 source.n419 104.615
R212 source.n450 source.n419 104.615
R213 source.n451 source.n450 104.615
R214 source.n452 source.n451 104.615
R215 source.n452 source.n415 104.615
R216 source.n459 source.n415 104.615
R217 source.n460 source.n459 104.615
R218 source.n460 source.n411 104.615
R219 source.n467 source.n411 104.615
R220 source.n468 source.n467 104.615
R221 source.n367 source.n361 104.615
R222 source.n368 source.n367 104.615
R223 source.n368 source.n357 104.615
R224 source.n375 source.n357 104.615
R225 source.n376 source.n375 104.615
R226 source.n376 source.n353 104.615
R227 source.n384 source.n353 104.615
R228 source.n385 source.n384 104.615
R229 source.n386 source.n385 104.615
R230 source.n386 source.n349 104.615
R231 source.n393 source.n349 104.615
R232 source.n394 source.n393 104.615
R233 source.n394 source.n345 104.615
R234 source.n401 source.n345 104.615
R235 source.n402 source.n401 104.615
R236 source.n297 source.n291 104.615
R237 source.n298 source.n297 104.615
R238 source.n298 source.n287 104.615
R239 source.n305 source.n287 104.615
R240 source.n306 source.n305 104.615
R241 source.n306 source.n283 104.615
R242 source.n314 source.n283 104.615
R243 source.n315 source.n314 104.615
R244 source.n316 source.n315 104.615
R245 source.n316 source.n279 104.615
R246 source.n323 source.n279 104.615
R247 source.n324 source.n323 104.615
R248 source.n324 source.n275 104.615
R249 source.n331 source.n275 104.615
R250 source.n332 source.n331 104.615
R251 source.n60 source.n59 104.615
R252 source.n59 source.n3 104.615
R253 source.n52 source.n3 104.615
R254 source.n52 source.n51 104.615
R255 source.n51 source.n7 104.615
R256 source.n44 source.n7 104.615
R257 source.n44 source.n43 104.615
R258 source.n43 source.n42 104.615
R259 source.n42 source.n11 104.615
R260 source.n35 source.n11 104.615
R261 source.n35 source.n34 104.615
R262 source.n34 source.n16 104.615
R263 source.n27 source.n16 104.615
R264 source.n27 source.n26 104.615
R265 source.n26 source.n20 104.615
R266 source.n130 source.n129 104.615
R267 source.n129 source.n73 104.615
R268 source.n122 source.n73 104.615
R269 source.n122 source.n121 104.615
R270 source.n121 source.n77 104.615
R271 source.n114 source.n77 104.615
R272 source.n114 source.n113 104.615
R273 source.n113 source.n112 104.615
R274 source.n112 source.n81 104.615
R275 source.n105 source.n81 104.615
R276 source.n105 source.n104 104.615
R277 source.n104 source.n86 104.615
R278 source.n97 source.n86 104.615
R279 source.n97 source.n96 104.615
R280 source.n96 source.n90 104.615
R281 source.n196 source.n195 104.615
R282 source.n195 source.n139 104.615
R283 source.n188 source.n139 104.615
R284 source.n188 source.n187 104.615
R285 source.n187 source.n143 104.615
R286 source.n180 source.n143 104.615
R287 source.n180 source.n179 104.615
R288 source.n179 source.n178 104.615
R289 source.n178 source.n147 104.615
R290 source.n171 source.n147 104.615
R291 source.n171 source.n170 104.615
R292 source.n170 source.n152 104.615
R293 source.n163 source.n152 104.615
R294 source.n163 source.n162 104.615
R295 source.n162 source.n156 104.615
R296 source.n266 source.n265 104.615
R297 source.n265 source.n209 104.615
R298 source.n258 source.n209 104.615
R299 source.n258 source.n257 104.615
R300 source.n257 source.n213 104.615
R301 source.n250 source.n213 104.615
R302 source.n250 source.n249 104.615
R303 source.n249 source.n248 104.615
R304 source.n248 source.n217 104.615
R305 source.n241 source.n217 104.615
R306 source.n241 source.n240 104.615
R307 source.n240 source.n222 104.615
R308 source.n233 source.n222 104.615
R309 source.n233 source.n232 104.615
R310 source.n232 source.n226 104.615
R311 source.t17 source.n497 52.3082
R312 source.t12 source.n427 52.3082
R313 source.t5 source.n361 52.3082
R314 source.t6 source.n291 52.3082
R315 source.t2 source.n20 52.3082
R316 source.t3 source.n90 52.3082
R317 source.t8 source.n156 52.3082
R318 source.t11 source.n226 52.3082
R319 source.n67 source.n66 42.8739
R320 source.n69 source.n68 42.8739
R321 source.n203 source.n202 42.8739
R322 source.n205 source.n204 42.8739
R323 source.n477 source.n476 42.8737
R324 source.n475 source.n474 42.8737
R325 source.n341 source.n340 42.8737
R326 source.n339 source.n338 42.8737
R327 source.n543 source.n542 29.8581
R328 source.n473 source.n472 29.8581
R329 source.n407 source.n406 29.8581
R330 source.n337 source.n336 29.8581
R331 source.n65 source.n64 29.8581
R332 source.n135 source.n134 29.8581
R333 source.n201 source.n200 29.8581
R334 source.n271 source.n270 29.8581
R335 source.n337 source.n271 22.0894
R336 source.n544 source.n65 16.4257
R337 source.n523 source.n488 13.1884
R338 source.n453 source.n418 13.1884
R339 source.n387 source.n352 13.1884
R340 source.n317 source.n282 13.1884
R341 source.n45 source.n10 13.1884
R342 source.n115 source.n80 13.1884
R343 source.n181 source.n146 13.1884
R344 source.n251 source.n216 13.1884
R345 source.n519 source.n518 12.8005
R346 source.n524 source.n486 12.8005
R347 source.n449 source.n448 12.8005
R348 source.n454 source.n416 12.8005
R349 source.n383 source.n382 12.8005
R350 source.n388 source.n350 12.8005
R351 source.n313 source.n312 12.8005
R352 source.n318 source.n280 12.8005
R353 source.n46 source.n8 12.8005
R354 source.n41 source.n12 12.8005
R355 source.n116 source.n78 12.8005
R356 source.n111 source.n82 12.8005
R357 source.n182 source.n144 12.8005
R358 source.n177 source.n148 12.8005
R359 source.n252 source.n214 12.8005
R360 source.n247 source.n218 12.8005
R361 source.n517 source.n490 12.0247
R362 source.n528 source.n527 12.0247
R363 source.n447 source.n420 12.0247
R364 source.n458 source.n457 12.0247
R365 source.n381 source.n354 12.0247
R366 source.n392 source.n391 12.0247
R367 source.n311 source.n284 12.0247
R368 source.n322 source.n321 12.0247
R369 source.n50 source.n49 12.0247
R370 source.n40 source.n13 12.0247
R371 source.n120 source.n119 12.0247
R372 source.n110 source.n83 12.0247
R373 source.n186 source.n185 12.0247
R374 source.n176 source.n149 12.0247
R375 source.n256 source.n255 12.0247
R376 source.n246 source.n219 12.0247
R377 source.n514 source.n513 11.249
R378 source.n531 source.n484 11.249
R379 source.n444 source.n443 11.249
R380 source.n461 source.n414 11.249
R381 source.n378 source.n377 11.249
R382 source.n395 source.n348 11.249
R383 source.n308 source.n307 11.249
R384 source.n325 source.n278 11.249
R385 source.n53 source.n6 11.249
R386 source.n37 source.n36 11.249
R387 source.n123 source.n76 11.249
R388 source.n107 source.n106 11.249
R389 source.n189 source.n142 11.249
R390 source.n173 source.n172 11.249
R391 source.n259 source.n212 11.249
R392 source.n243 source.n242 11.249
R393 source.n510 source.n492 10.4732
R394 source.n532 source.n482 10.4732
R395 source.n440 source.n422 10.4732
R396 source.n462 source.n412 10.4732
R397 source.n374 source.n356 10.4732
R398 source.n396 source.n346 10.4732
R399 source.n304 source.n286 10.4732
R400 source.n326 source.n276 10.4732
R401 source.n54 source.n4 10.4732
R402 source.n33 source.n15 10.4732
R403 source.n124 source.n74 10.4732
R404 source.n103 source.n85 10.4732
R405 source.n190 source.n140 10.4732
R406 source.n169 source.n151 10.4732
R407 source.n260 source.n210 10.4732
R408 source.n239 source.n221 10.4732
R409 source.n499 source.n498 10.2747
R410 source.n429 source.n428 10.2747
R411 source.n363 source.n362 10.2747
R412 source.n293 source.n292 10.2747
R413 source.n22 source.n21 10.2747
R414 source.n92 source.n91 10.2747
R415 source.n158 source.n157 10.2747
R416 source.n228 source.n227 10.2747
R417 source.n509 source.n494 9.69747
R418 source.n536 source.n535 9.69747
R419 source.n439 source.n424 9.69747
R420 source.n466 source.n465 9.69747
R421 source.n373 source.n358 9.69747
R422 source.n400 source.n399 9.69747
R423 source.n303 source.n288 9.69747
R424 source.n330 source.n329 9.69747
R425 source.n58 source.n57 9.69747
R426 source.n32 source.n17 9.69747
R427 source.n128 source.n127 9.69747
R428 source.n102 source.n87 9.69747
R429 source.n194 source.n193 9.69747
R430 source.n168 source.n153 9.69747
R431 source.n264 source.n263 9.69747
R432 source.n238 source.n223 9.69747
R433 source.n542 source.n541 9.45567
R434 source.n472 source.n471 9.45567
R435 source.n406 source.n405 9.45567
R436 source.n336 source.n335 9.45567
R437 source.n64 source.n63 9.45567
R438 source.n134 source.n133 9.45567
R439 source.n200 source.n199 9.45567
R440 source.n270 source.n269 9.45567
R441 source.n541 source.n540 9.3005
R442 source.n480 source.n479 9.3005
R443 source.n535 source.n534 9.3005
R444 source.n533 source.n532 9.3005
R445 source.n484 source.n483 9.3005
R446 source.n527 source.n526 9.3005
R447 source.n525 source.n524 9.3005
R448 source.n501 source.n500 9.3005
R449 source.n496 source.n495 9.3005
R450 source.n507 source.n506 9.3005
R451 source.n509 source.n508 9.3005
R452 source.n492 source.n491 9.3005
R453 source.n515 source.n514 9.3005
R454 source.n517 source.n516 9.3005
R455 source.n518 source.n487 9.3005
R456 source.n471 source.n470 9.3005
R457 source.n410 source.n409 9.3005
R458 source.n465 source.n464 9.3005
R459 source.n463 source.n462 9.3005
R460 source.n414 source.n413 9.3005
R461 source.n457 source.n456 9.3005
R462 source.n455 source.n454 9.3005
R463 source.n431 source.n430 9.3005
R464 source.n426 source.n425 9.3005
R465 source.n437 source.n436 9.3005
R466 source.n439 source.n438 9.3005
R467 source.n422 source.n421 9.3005
R468 source.n445 source.n444 9.3005
R469 source.n447 source.n446 9.3005
R470 source.n448 source.n417 9.3005
R471 source.n405 source.n404 9.3005
R472 source.n344 source.n343 9.3005
R473 source.n399 source.n398 9.3005
R474 source.n397 source.n396 9.3005
R475 source.n348 source.n347 9.3005
R476 source.n391 source.n390 9.3005
R477 source.n389 source.n388 9.3005
R478 source.n365 source.n364 9.3005
R479 source.n360 source.n359 9.3005
R480 source.n371 source.n370 9.3005
R481 source.n373 source.n372 9.3005
R482 source.n356 source.n355 9.3005
R483 source.n379 source.n378 9.3005
R484 source.n381 source.n380 9.3005
R485 source.n382 source.n351 9.3005
R486 source.n335 source.n334 9.3005
R487 source.n274 source.n273 9.3005
R488 source.n329 source.n328 9.3005
R489 source.n327 source.n326 9.3005
R490 source.n278 source.n277 9.3005
R491 source.n321 source.n320 9.3005
R492 source.n319 source.n318 9.3005
R493 source.n295 source.n294 9.3005
R494 source.n290 source.n289 9.3005
R495 source.n301 source.n300 9.3005
R496 source.n303 source.n302 9.3005
R497 source.n286 source.n285 9.3005
R498 source.n309 source.n308 9.3005
R499 source.n311 source.n310 9.3005
R500 source.n312 source.n281 9.3005
R501 source.n24 source.n23 9.3005
R502 source.n19 source.n18 9.3005
R503 source.n30 source.n29 9.3005
R504 source.n32 source.n31 9.3005
R505 source.n15 source.n14 9.3005
R506 source.n38 source.n37 9.3005
R507 source.n40 source.n39 9.3005
R508 source.n12 source.n9 9.3005
R509 source.n63 source.n62 9.3005
R510 source.n2 source.n1 9.3005
R511 source.n57 source.n56 9.3005
R512 source.n55 source.n54 9.3005
R513 source.n6 source.n5 9.3005
R514 source.n49 source.n48 9.3005
R515 source.n47 source.n46 9.3005
R516 source.n94 source.n93 9.3005
R517 source.n89 source.n88 9.3005
R518 source.n100 source.n99 9.3005
R519 source.n102 source.n101 9.3005
R520 source.n85 source.n84 9.3005
R521 source.n108 source.n107 9.3005
R522 source.n110 source.n109 9.3005
R523 source.n82 source.n79 9.3005
R524 source.n133 source.n132 9.3005
R525 source.n72 source.n71 9.3005
R526 source.n127 source.n126 9.3005
R527 source.n125 source.n124 9.3005
R528 source.n76 source.n75 9.3005
R529 source.n119 source.n118 9.3005
R530 source.n117 source.n116 9.3005
R531 source.n160 source.n159 9.3005
R532 source.n155 source.n154 9.3005
R533 source.n166 source.n165 9.3005
R534 source.n168 source.n167 9.3005
R535 source.n151 source.n150 9.3005
R536 source.n174 source.n173 9.3005
R537 source.n176 source.n175 9.3005
R538 source.n148 source.n145 9.3005
R539 source.n199 source.n198 9.3005
R540 source.n138 source.n137 9.3005
R541 source.n193 source.n192 9.3005
R542 source.n191 source.n190 9.3005
R543 source.n142 source.n141 9.3005
R544 source.n185 source.n184 9.3005
R545 source.n183 source.n182 9.3005
R546 source.n230 source.n229 9.3005
R547 source.n225 source.n224 9.3005
R548 source.n236 source.n235 9.3005
R549 source.n238 source.n237 9.3005
R550 source.n221 source.n220 9.3005
R551 source.n244 source.n243 9.3005
R552 source.n246 source.n245 9.3005
R553 source.n218 source.n215 9.3005
R554 source.n269 source.n268 9.3005
R555 source.n208 source.n207 9.3005
R556 source.n263 source.n262 9.3005
R557 source.n261 source.n260 9.3005
R558 source.n212 source.n211 9.3005
R559 source.n255 source.n254 9.3005
R560 source.n253 source.n252 9.3005
R561 source.n506 source.n505 8.92171
R562 source.n539 source.n480 8.92171
R563 source.n436 source.n435 8.92171
R564 source.n469 source.n410 8.92171
R565 source.n370 source.n369 8.92171
R566 source.n403 source.n344 8.92171
R567 source.n300 source.n299 8.92171
R568 source.n333 source.n274 8.92171
R569 source.n61 source.n2 8.92171
R570 source.n29 source.n28 8.92171
R571 source.n131 source.n72 8.92171
R572 source.n99 source.n98 8.92171
R573 source.n197 source.n138 8.92171
R574 source.n165 source.n164 8.92171
R575 source.n267 source.n208 8.92171
R576 source.n235 source.n234 8.92171
R577 source.n502 source.n496 8.14595
R578 source.n540 source.n478 8.14595
R579 source.n432 source.n426 8.14595
R580 source.n470 source.n408 8.14595
R581 source.n366 source.n360 8.14595
R582 source.n404 source.n342 8.14595
R583 source.n296 source.n290 8.14595
R584 source.n334 source.n272 8.14595
R585 source.n62 source.n0 8.14595
R586 source.n25 source.n19 8.14595
R587 source.n132 source.n70 8.14595
R588 source.n95 source.n89 8.14595
R589 source.n198 source.n136 8.14595
R590 source.n161 source.n155 8.14595
R591 source.n268 source.n206 8.14595
R592 source.n231 source.n225 8.14595
R593 source.n501 source.n498 7.3702
R594 source.n431 source.n428 7.3702
R595 source.n365 source.n362 7.3702
R596 source.n295 source.n292 7.3702
R597 source.n24 source.n21 7.3702
R598 source.n94 source.n91 7.3702
R599 source.n160 source.n157 7.3702
R600 source.n230 source.n227 7.3702
R601 source.n502 source.n501 5.81868
R602 source.n542 source.n478 5.81868
R603 source.n432 source.n431 5.81868
R604 source.n472 source.n408 5.81868
R605 source.n366 source.n365 5.81868
R606 source.n406 source.n342 5.81868
R607 source.n296 source.n295 5.81868
R608 source.n336 source.n272 5.81868
R609 source.n64 source.n0 5.81868
R610 source.n25 source.n24 5.81868
R611 source.n134 source.n70 5.81868
R612 source.n95 source.n94 5.81868
R613 source.n200 source.n136 5.81868
R614 source.n161 source.n160 5.81868
R615 source.n270 source.n206 5.81868
R616 source.n231 source.n230 5.81868
R617 source.n544 source.n543 5.66429
R618 source.n505 source.n496 5.04292
R619 source.n540 source.n539 5.04292
R620 source.n435 source.n426 5.04292
R621 source.n470 source.n469 5.04292
R622 source.n369 source.n360 5.04292
R623 source.n404 source.n403 5.04292
R624 source.n299 source.n290 5.04292
R625 source.n334 source.n333 5.04292
R626 source.n62 source.n61 5.04292
R627 source.n28 source.n19 5.04292
R628 source.n132 source.n131 5.04292
R629 source.n98 source.n89 5.04292
R630 source.n198 source.n197 5.04292
R631 source.n164 source.n155 5.04292
R632 source.n268 source.n267 5.04292
R633 source.n234 source.n225 5.04292
R634 source.n506 source.n494 4.26717
R635 source.n536 source.n480 4.26717
R636 source.n436 source.n424 4.26717
R637 source.n466 source.n410 4.26717
R638 source.n370 source.n358 4.26717
R639 source.n400 source.n344 4.26717
R640 source.n300 source.n288 4.26717
R641 source.n330 source.n274 4.26717
R642 source.n58 source.n2 4.26717
R643 source.n29 source.n17 4.26717
R644 source.n128 source.n72 4.26717
R645 source.n99 source.n87 4.26717
R646 source.n194 source.n138 4.26717
R647 source.n165 source.n153 4.26717
R648 source.n264 source.n208 4.26717
R649 source.n235 source.n223 4.26717
R650 source.n510 source.n509 3.49141
R651 source.n535 source.n482 3.49141
R652 source.n440 source.n439 3.49141
R653 source.n465 source.n412 3.49141
R654 source.n374 source.n373 3.49141
R655 source.n399 source.n346 3.49141
R656 source.n304 source.n303 3.49141
R657 source.n329 source.n276 3.49141
R658 source.n57 source.n4 3.49141
R659 source.n33 source.n32 3.49141
R660 source.n127 source.n74 3.49141
R661 source.n103 source.n102 3.49141
R662 source.n193 source.n140 3.49141
R663 source.n169 source.n168 3.49141
R664 source.n263 source.n210 3.49141
R665 source.n239 source.n238 3.49141
R666 source.n500 source.n499 2.84303
R667 source.n430 source.n429 2.84303
R668 source.n364 source.n363 2.84303
R669 source.n294 source.n293 2.84303
R670 source.n23 source.n22 2.84303
R671 source.n93 source.n92 2.84303
R672 source.n159 source.n158 2.84303
R673 source.n229 source.n228 2.84303
R674 source.n513 source.n492 2.71565
R675 source.n532 source.n531 2.71565
R676 source.n443 source.n422 2.71565
R677 source.n462 source.n461 2.71565
R678 source.n377 source.n356 2.71565
R679 source.n396 source.n395 2.71565
R680 source.n307 source.n286 2.71565
R681 source.n326 source.n325 2.71565
R682 source.n54 source.n53 2.71565
R683 source.n36 source.n15 2.71565
R684 source.n124 source.n123 2.71565
R685 source.n106 source.n85 2.71565
R686 source.n190 source.n189 2.71565
R687 source.n172 source.n151 2.71565
R688 source.n260 source.n259 2.71565
R689 source.n242 source.n221 2.71565
R690 source.n514 source.n490 1.93989
R691 source.n528 source.n484 1.93989
R692 source.n444 source.n420 1.93989
R693 source.n458 source.n414 1.93989
R694 source.n378 source.n354 1.93989
R695 source.n392 source.n348 1.93989
R696 source.n308 source.n284 1.93989
R697 source.n322 source.n278 1.93989
R698 source.n50 source.n6 1.93989
R699 source.n37 source.n13 1.93989
R700 source.n120 source.n76 1.93989
R701 source.n107 source.n83 1.93989
R702 source.n186 source.n142 1.93989
R703 source.n173 source.n149 1.93989
R704 source.n256 source.n212 1.93989
R705 source.n243 source.n219 1.93989
R706 source.n476 source.t9 1.6505
R707 source.n476 source.t13 1.6505
R708 source.n474 source.t10 1.6505
R709 source.n474 source.t15 1.6505
R710 source.n340 source.t1 1.6505
R711 source.n340 source.t20 1.6505
R712 source.n338 source.t4 1.6505
R713 source.n338 source.t7 1.6505
R714 source.n66 source.t22 1.6505
R715 source.n66 source.t21 1.6505
R716 source.n68 source.t0 1.6505
R717 source.n68 source.t23 1.6505
R718 source.n202 source.t14 1.6505
R719 source.n202 source.t18 1.6505
R720 source.n204 source.t19 1.6505
R721 source.n204 source.t16 1.6505
R722 source.n519 source.n517 1.16414
R723 source.n527 source.n486 1.16414
R724 source.n449 source.n447 1.16414
R725 source.n457 source.n416 1.16414
R726 source.n383 source.n381 1.16414
R727 source.n391 source.n350 1.16414
R728 source.n313 source.n311 1.16414
R729 source.n321 source.n280 1.16414
R730 source.n49 source.n8 1.16414
R731 source.n41 source.n40 1.16414
R732 source.n119 source.n78 1.16414
R733 source.n111 source.n110 1.16414
R734 source.n185 source.n144 1.16414
R735 source.n177 source.n176 1.16414
R736 source.n255 source.n214 1.16414
R737 source.n247 source.n246 1.16414
R738 source.n271 source.n205 0.802224
R739 source.n205 source.n203 0.802224
R740 source.n203 source.n201 0.802224
R741 source.n135 source.n69 0.802224
R742 source.n69 source.n67 0.802224
R743 source.n67 source.n65 0.802224
R744 source.n339 source.n337 0.802224
R745 source.n341 source.n339 0.802224
R746 source.n407 source.n341 0.802224
R747 source.n475 source.n473 0.802224
R748 source.n477 source.n475 0.802224
R749 source.n543 source.n477 0.802224
R750 source.n201 source.n135 0.470328
R751 source.n473 source.n407 0.470328
R752 source.n518 source.n488 0.388379
R753 source.n524 source.n523 0.388379
R754 source.n448 source.n418 0.388379
R755 source.n454 source.n453 0.388379
R756 source.n382 source.n352 0.388379
R757 source.n388 source.n387 0.388379
R758 source.n312 source.n282 0.388379
R759 source.n318 source.n317 0.388379
R760 source.n46 source.n45 0.388379
R761 source.n12 source.n10 0.388379
R762 source.n116 source.n115 0.388379
R763 source.n82 source.n80 0.388379
R764 source.n182 source.n181 0.388379
R765 source.n148 source.n146 0.388379
R766 source.n252 source.n251 0.388379
R767 source.n218 source.n216 0.388379
R768 source source.n544 0.188
R769 source.n500 source.n495 0.155672
R770 source.n507 source.n495 0.155672
R771 source.n508 source.n507 0.155672
R772 source.n508 source.n491 0.155672
R773 source.n515 source.n491 0.155672
R774 source.n516 source.n515 0.155672
R775 source.n516 source.n487 0.155672
R776 source.n525 source.n487 0.155672
R777 source.n526 source.n525 0.155672
R778 source.n526 source.n483 0.155672
R779 source.n533 source.n483 0.155672
R780 source.n534 source.n533 0.155672
R781 source.n534 source.n479 0.155672
R782 source.n541 source.n479 0.155672
R783 source.n430 source.n425 0.155672
R784 source.n437 source.n425 0.155672
R785 source.n438 source.n437 0.155672
R786 source.n438 source.n421 0.155672
R787 source.n445 source.n421 0.155672
R788 source.n446 source.n445 0.155672
R789 source.n446 source.n417 0.155672
R790 source.n455 source.n417 0.155672
R791 source.n456 source.n455 0.155672
R792 source.n456 source.n413 0.155672
R793 source.n463 source.n413 0.155672
R794 source.n464 source.n463 0.155672
R795 source.n464 source.n409 0.155672
R796 source.n471 source.n409 0.155672
R797 source.n364 source.n359 0.155672
R798 source.n371 source.n359 0.155672
R799 source.n372 source.n371 0.155672
R800 source.n372 source.n355 0.155672
R801 source.n379 source.n355 0.155672
R802 source.n380 source.n379 0.155672
R803 source.n380 source.n351 0.155672
R804 source.n389 source.n351 0.155672
R805 source.n390 source.n389 0.155672
R806 source.n390 source.n347 0.155672
R807 source.n397 source.n347 0.155672
R808 source.n398 source.n397 0.155672
R809 source.n398 source.n343 0.155672
R810 source.n405 source.n343 0.155672
R811 source.n294 source.n289 0.155672
R812 source.n301 source.n289 0.155672
R813 source.n302 source.n301 0.155672
R814 source.n302 source.n285 0.155672
R815 source.n309 source.n285 0.155672
R816 source.n310 source.n309 0.155672
R817 source.n310 source.n281 0.155672
R818 source.n319 source.n281 0.155672
R819 source.n320 source.n319 0.155672
R820 source.n320 source.n277 0.155672
R821 source.n327 source.n277 0.155672
R822 source.n328 source.n327 0.155672
R823 source.n328 source.n273 0.155672
R824 source.n335 source.n273 0.155672
R825 source.n63 source.n1 0.155672
R826 source.n56 source.n1 0.155672
R827 source.n56 source.n55 0.155672
R828 source.n55 source.n5 0.155672
R829 source.n48 source.n5 0.155672
R830 source.n48 source.n47 0.155672
R831 source.n47 source.n9 0.155672
R832 source.n39 source.n9 0.155672
R833 source.n39 source.n38 0.155672
R834 source.n38 source.n14 0.155672
R835 source.n31 source.n14 0.155672
R836 source.n31 source.n30 0.155672
R837 source.n30 source.n18 0.155672
R838 source.n23 source.n18 0.155672
R839 source.n133 source.n71 0.155672
R840 source.n126 source.n71 0.155672
R841 source.n126 source.n125 0.155672
R842 source.n125 source.n75 0.155672
R843 source.n118 source.n75 0.155672
R844 source.n118 source.n117 0.155672
R845 source.n117 source.n79 0.155672
R846 source.n109 source.n79 0.155672
R847 source.n109 source.n108 0.155672
R848 source.n108 source.n84 0.155672
R849 source.n101 source.n84 0.155672
R850 source.n101 source.n100 0.155672
R851 source.n100 source.n88 0.155672
R852 source.n93 source.n88 0.155672
R853 source.n199 source.n137 0.155672
R854 source.n192 source.n137 0.155672
R855 source.n192 source.n191 0.155672
R856 source.n191 source.n141 0.155672
R857 source.n184 source.n141 0.155672
R858 source.n184 source.n183 0.155672
R859 source.n183 source.n145 0.155672
R860 source.n175 source.n145 0.155672
R861 source.n175 source.n174 0.155672
R862 source.n174 source.n150 0.155672
R863 source.n167 source.n150 0.155672
R864 source.n167 source.n166 0.155672
R865 source.n166 source.n154 0.155672
R866 source.n159 source.n154 0.155672
R867 source.n269 source.n207 0.155672
R868 source.n262 source.n207 0.155672
R869 source.n262 source.n261 0.155672
R870 source.n261 source.n211 0.155672
R871 source.n254 source.n211 0.155672
R872 source.n254 source.n253 0.155672
R873 source.n253 source.n215 0.155672
R874 source.n245 source.n215 0.155672
R875 source.n245 source.n244 0.155672
R876 source.n244 source.n220 0.155672
R877 source.n237 source.n220 0.155672
R878 source.n237 source.n236 0.155672
R879 source.n236 source.n224 0.155672
R880 source.n229 source.n224 0.155672
R881 drain_right.n6 drain_right.n4 60.3542
R882 drain_right.n3 drain_right.n2 60.2989
R883 drain_right.n3 drain_right.n0 60.2989
R884 drain_right.n6 drain_right.n5 59.5527
R885 drain_right.n8 drain_right.n7 59.5527
R886 drain_right.n3 drain_right.n1 59.5525
R887 drain_right drain_right.n3 30.8225
R888 drain_right drain_right.n8 6.45494
R889 drain_right.n1 drain_right.t6 1.6505
R890 drain_right.n1 drain_right.t0 1.6505
R891 drain_right.n2 drain_right.t10 1.6505
R892 drain_right.n2 drain_right.t11 1.6505
R893 drain_right.n0 drain_right.t3 1.6505
R894 drain_right.n0 drain_right.t9 1.6505
R895 drain_right.n4 drain_right.t2 1.6505
R896 drain_right.n4 drain_right.t1 1.6505
R897 drain_right.n5 drain_right.t5 1.6505
R898 drain_right.n5 drain_right.t4 1.6505
R899 drain_right.n7 drain_right.t7 1.6505
R900 drain_right.n7 drain_right.t8 1.6505
R901 drain_right.n8 drain_right.n6 0.802224
R902 plus.n4 plus.t9 572.532
R903 plus.n16 plus.t10 572.532
R904 plus.n10 plus.t2 547.472
R905 plus.n8 plus.t4 547.472
R906 plus.n7 plus.t5 547.472
R907 plus.n6 plus.t6 547.472
R908 plus.n5 plus.t8 547.472
R909 plus.n22 plus.t1 547.472
R910 plus.n20 plus.t0 547.472
R911 plus.n19 plus.t11 547.472
R912 plus.n18 plus.t7 547.472
R913 plus.n17 plus.t3 547.472
R914 plus.n8 plus.n1 161.3
R915 plus.n9 plus.n0 161.3
R916 plus.n11 plus.n10 161.3
R917 plus.n20 plus.n13 161.3
R918 plus.n21 plus.n12 161.3
R919 plus.n23 plus.n22 161.3
R920 plus.n6 plus.n3 80.6037
R921 plus.n7 plus.n2 80.6037
R922 plus.n18 plus.n15 80.6037
R923 plus.n19 plus.n14 80.6037
R924 plus.n8 plus.n7 48.2005
R925 plus.n7 plus.n6 48.2005
R926 plus.n6 plus.n5 48.2005
R927 plus.n20 plus.n19 48.2005
R928 plus.n19 plus.n18 48.2005
R929 plus.n18 plus.n17 48.2005
R930 plus.n4 plus.n3 45.0744
R931 plus.n16 plus.n15 45.0744
R932 plus.n10 plus.n9 40.1672
R933 plus.n22 plus.n21 40.1672
R934 plus plus.n23 30.7339
R935 plus.n5 plus.n4 16.1124
R936 plus.n17 plus.n16 16.1124
R937 plus plus.n11 12.2316
R938 plus.n9 plus.n8 8.03383
R939 plus.n21 plus.n20 8.03383
R940 plus.n3 plus.n2 0.380177
R941 plus.n15 plus.n14 0.380177
R942 plus.n2 plus.n1 0.285035
R943 plus.n14 plus.n13 0.285035
R944 plus.n1 plus.n0 0.189894
R945 plus.n11 plus.n0 0.189894
R946 plus.n23 plus.n12 0.189894
R947 plus.n13 plus.n12 0.189894
R948 drain_left.n6 drain_left.n4 60.3544
R949 drain_left.n3 drain_left.n2 60.2989
R950 drain_left.n3 drain_left.n0 60.2989
R951 drain_left.n6 drain_left.n5 59.5527
R952 drain_left.n3 drain_left.n1 59.5525
R953 drain_left.n8 drain_left.n7 59.5525
R954 drain_left drain_left.n3 31.3757
R955 drain_left drain_left.n8 6.45494
R956 drain_left.n1 drain_left.t0 1.6505
R957 drain_left.n1 drain_left.t4 1.6505
R958 drain_left.n2 drain_left.t8 1.6505
R959 drain_left.n2 drain_left.t1 1.6505
R960 drain_left.n0 drain_left.t10 1.6505
R961 drain_left.n0 drain_left.t11 1.6505
R962 drain_left.n7 drain_left.t7 1.6505
R963 drain_left.n7 drain_left.t9 1.6505
R964 drain_left.n5 drain_left.t5 1.6505
R965 drain_left.n5 drain_left.t6 1.6505
R966 drain_left.n4 drain_left.t2 1.6505
R967 drain_left.n4 drain_left.t3 1.6505
R968 drain_left.n8 drain_left.n6 0.802224
C0 minus drain_right 7.22362f
C1 minus source 7.0638f
C2 drain_right source 16.7151f
C3 plus minus 5.66402f
C4 plus drain_right 0.352374f
C5 minus drain_left 0.17204f
C6 drain_right drain_left 1.01253f
C7 plus source 7.07784f
C8 drain_left source 16.7136f
C9 plus drain_left 7.42079f
C10 drain_right a_n2018_n3288# 6.13158f
C11 drain_left a_n2018_n3288# 6.42768f
C12 source a_n2018_n3288# 9.009165f
C13 minus a_n2018_n3288# 7.931088f
C14 plus a_n2018_n3288# 9.698441f
C15 drain_left.t10 a_n2018_n3288# 0.265541f
C16 drain_left.t11 a_n2018_n3288# 0.265541f
C17 drain_left.n0 a_n2018_n3288# 2.3677f
C18 drain_left.t0 a_n2018_n3288# 0.265541f
C19 drain_left.t4 a_n2018_n3288# 0.265541f
C20 drain_left.n1 a_n2018_n3288# 2.36291f
C21 drain_left.t8 a_n2018_n3288# 0.265541f
C22 drain_left.t1 a_n2018_n3288# 0.265541f
C23 drain_left.n2 a_n2018_n3288# 2.3677f
C24 drain_left.n3 a_n2018_n3288# 2.5147f
C25 drain_left.t2 a_n2018_n3288# 0.265541f
C26 drain_left.t3 a_n2018_n3288# 0.265541f
C27 drain_left.n4 a_n2018_n3288# 2.36811f
C28 drain_left.t5 a_n2018_n3288# 0.265541f
C29 drain_left.t6 a_n2018_n3288# 0.265541f
C30 drain_left.n5 a_n2018_n3288# 2.36292f
C31 drain_left.n6 a_n2018_n3288# 0.765451f
C32 drain_left.t7 a_n2018_n3288# 0.265541f
C33 drain_left.t9 a_n2018_n3288# 0.265541f
C34 drain_left.n7 a_n2018_n3288# 2.36291f
C35 drain_left.n8 a_n2018_n3288# 0.623872f
C36 plus.n0 a_n2018_n3288# 0.044769f
C37 plus.t2 a_n2018_n3288# 0.91915f
C38 plus.t4 a_n2018_n3288# 0.91915f
C39 plus.n1 a_n2018_n3288# 0.059739f
C40 plus.t5 a_n2018_n3288# 0.91915f
C41 plus.n2 a_n2018_n3288# 0.074569f
C42 plus.t6 a_n2018_n3288# 0.91915f
C43 plus.n3 a_n2018_n3288# 0.229448f
C44 plus.t8 a_n2018_n3288# 0.91915f
C45 plus.t9 a_n2018_n3288# 0.935268f
C46 plus.n4 a_n2018_n3288# 0.35555f
C47 plus.n5 a_n2018_n3288# 0.37726f
C48 plus.n6 a_n2018_n3288# 0.378894f
C49 plus.n7 a_n2018_n3288# 0.378894f
C50 plus.n8 a_n2018_n3288# 0.370253f
C51 plus.n9 a_n2018_n3288# 0.010159f
C52 plus.n10 a_n2018_n3288# 0.367217f
C53 plus.n11 a_n2018_n3288# 0.510256f
C54 plus.n12 a_n2018_n3288# 0.044769f
C55 plus.t1 a_n2018_n3288# 0.91915f
C56 plus.n13 a_n2018_n3288# 0.059739f
C57 plus.t0 a_n2018_n3288# 0.91915f
C58 plus.n14 a_n2018_n3288# 0.074569f
C59 plus.t11 a_n2018_n3288# 0.91915f
C60 plus.n15 a_n2018_n3288# 0.229448f
C61 plus.t7 a_n2018_n3288# 0.91915f
C62 plus.t10 a_n2018_n3288# 0.935268f
C63 plus.n16 a_n2018_n3288# 0.35555f
C64 plus.t3 a_n2018_n3288# 0.91915f
C65 plus.n17 a_n2018_n3288# 0.37726f
C66 plus.n18 a_n2018_n3288# 0.378894f
C67 plus.n19 a_n2018_n3288# 0.378894f
C68 plus.n20 a_n2018_n3288# 0.370253f
C69 plus.n21 a_n2018_n3288# 0.010159f
C70 plus.n22 a_n2018_n3288# 0.367217f
C71 plus.n23 a_n2018_n3288# 1.38184f
C72 drain_right.t3 a_n2018_n3288# 0.26454f
C73 drain_right.t9 a_n2018_n3288# 0.26454f
C74 drain_right.n0 a_n2018_n3288# 2.35877f
C75 drain_right.t6 a_n2018_n3288# 0.26454f
C76 drain_right.t0 a_n2018_n3288# 0.26454f
C77 drain_right.n1 a_n2018_n3288# 2.354f
C78 drain_right.t10 a_n2018_n3288# 0.26454f
C79 drain_right.t11 a_n2018_n3288# 0.26454f
C80 drain_right.n2 a_n2018_n3288# 2.35877f
C81 drain_right.n3 a_n2018_n3288# 2.44752f
C82 drain_right.t2 a_n2018_n3288# 0.26454f
C83 drain_right.t1 a_n2018_n3288# 0.26454f
C84 drain_right.n4 a_n2018_n3288# 2.35917f
C85 drain_right.t5 a_n2018_n3288# 0.26454f
C86 drain_right.t4 a_n2018_n3288# 0.26454f
C87 drain_right.n5 a_n2018_n3288# 2.35401f
C88 drain_right.n6 a_n2018_n3288# 0.762574f
C89 drain_right.t7 a_n2018_n3288# 0.26454f
C90 drain_right.t8 a_n2018_n3288# 0.26454f
C91 drain_right.n7 a_n2018_n3288# 2.35401f
C92 drain_right.n8 a_n2018_n3288# 0.62151f
C93 source.n0 a_n2018_n3288# 0.029898f
C94 source.n1 a_n2018_n3288# 0.022571f
C95 source.n2 a_n2018_n3288# 0.012129f
C96 source.n3 a_n2018_n3288# 0.028668f
C97 source.n4 a_n2018_n3288# 0.012842f
C98 source.n5 a_n2018_n3288# 0.022571f
C99 source.n6 a_n2018_n3288# 0.012129f
C100 source.n7 a_n2018_n3288# 0.028668f
C101 source.n8 a_n2018_n3288# 0.012842f
C102 source.n9 a_n2018_n3288# 0.022571f
C103 source.n10 a_n2018_n3288# 0.012486f
C104 source.n11 a_n2018_n3288# 0.028668f
C105 source.n12 a_n2018_n3288# 0.012129f
C106 source.n13 a_n2018_n3288# 0.012842f
C107 source.n14 a_n2018_n3288# 0.022571f
C108 source.n15 a_n2018_n3288# 0.012129f
C109 source.n16 a_n2018_n3288# 0.028668f
C110 source.n17 a_n2018_n3288# 0.012842f
C111 source.n18 a_n2018_n3288# 0.022571f
C112 source.n19 a_n2018_n3288# 0.012129f
C113 source.n20 a_n2018_n3288# 0.021501f
C114 source.n21 a_n2018_n3288# 0.020266f
C115 source.t2 a_n2018_n3288# 0.048418f
C116 source.n22 a_n2018_n3288# 0.162736f
C117 source.n23 a_n2018_n3288# 1.13868f
C118 source.n24 a_n2018_n3288# 0.012129f
C119 source.n25 a_n2018_n3288# 0.012842f
C120 source.n26 a_n2018_n3288# 0.028668f
C121 source.n27 a_n2018_n3288# 0.028668f
C122 source.n28 a_n2018_n3288# 0.012842f
C123 source.n29 a_n2018_n3288# 0.012129f
C124 source.n30 a_n2018_n3288# 0.022571f
C125 source.n31 a_n2018_n3288# 0.022571f
C126 source.n32 a_n2018_n3288# 0.012129f
C127 source.n33 a_n2018_n3288# 0.012842f
C128 source.n34 a_n2018_n3288# 0.028668f
C129 source.n35 a_n2018_n3288# 0.028668f
C130 source.n36 a_n2018_n3288# 0.012842f
C131 source.n37 a_n2018_n3288# 0.012129f
C132 source.n38 a_n2018_n3288# 0.022571f
C133 source.n39 a_n2018_n3288# 0.022571f
C134 source.n40 a_n2018_n3288# 0.012129f
C135 source.n41 a_n2018_n3288# 0.012842f
C136 source.n42 a_n2018_n3288# 0.028668f
C137 source.n43 a_n2018_n3288# 0.028668f
C138 source.n44 a_n2018_n3288# 0.028668f
C139 source.n45 a_n2018_n3288# 0.012486f
C140 source.n46 a_n2018_n3288# 0.012129f
C141 source.n47 a_n2018_n3288# 0.022571f
C142 source.n48 a_n2018_n3288# 0.022571f
C143 source.n49 a_n2018_n3288# 0.012129f
C144 source.n50 a_n2018_n3288# 0.012842f
C145 source.n51 a_n2018_n3288# 0.028668f
C146 source.n52 a_n2018_n3288# 0.028668f
C147 source.n53 a_n2018_n3288# 0.012842f
C148 source.n54 a_n2018_n3288# 0.012129f
C149 source.n55 a_n2018_n3288# 0.022571f
C150 source.n56 a_n2018_n3288# 0.022571f
C151 source.n57 a_n2018_n3288# 0.012129f
C152 source.n58 a_n2018_n3288# 0.012842f
C153 source.n59 a_n2018_n3288# 0.028668f
C154 source.n60 a_n2018_n3288# 0.05883f
C155 source.n61 a_n2018_n3288# 0.012842f
C156 source.n62 a_n2018_n3288# 0.012129f
C157 source.n63 a_n2018_n3288# 0.048472f
C158 source.n64 a_n2018_n3288# 0.032468f
C159 source.n65 a_n2018_n3288# 0.939219f
C160 source.t22 a_n2018_n3288# 0.214038f
C161 source.t21 a_n2018_n3288# 0.214038f
C162 source.n66 a_n2018_n3288# 1.83259f
C163 source.n67 a_n2018_n3288# 0.34738f
C164 source.t0 a_n2018_n3288# 0.214038f
C165 source.t23 a_n2018_n3288# 0.214038f
C166 source.n68 a_n2018_n3288# 1.83259f
C167 source.n69 a_n2018_n3288# 0.34738f
C168 source.n70 a_n2018_n3288# 0.029898f
C169 source.n71 a_n2018_n3288# 0.022571f
C170 source.n72 a_n2018_n3288# 0.012129f
C171 source.n73 a_n2018_n3288# 0.028668f
C172 source.n74 a_n2018_n3288# 0.012842f
C173 source.n75 a_n2018_n3288# 0.022571f
C174 source.n76 a_n2018_n3288# 0.012129f
C175 source.n77 a_n2018_n3288# 0.028668f
C176 source.n78 a_n2018_n3288# 0.012842f
C177 source.n79 a_n2018_n3288# 0.022571f
C178 source.n80 a_n2018_n3288# 0.012486f
C179 source.n81 a_n2018_n3288# 0.028668f
C180 source.n82 a_n2018_n3288# 0.012129f
C181 source.n83 a_n2018_n3288# 0.012842f
C182 source.n84 a_n2018_n3288# 0.022571f
C183 source.n85 a_n2018_n3288# 0.012129f
C184 source.n86 a_n2018_n3288# 0.028668f
C185 source.n87 a_n2018_n3288# 0.012842f
C186 source.n88 a_n2018_n3288# 0.022571f
C187 source.n89 a_n2018_n3288# 0.012129f
C188 source.n90 a_n2018_n3288# 0.021501f
C189 source.n91 a_n2018_n3288# 0.020266f
C190 source.t3 a_n2018_n3288# 0.048418f
C191 source.n92 a_n2018_n3288# 0.162736f
C192 source.n93 a_n2018_n3288# 1.13868f
C193 source.n94 a_n2018_n3288# 0.012129f
C194 source.n95 a_n2018_n3288# 0.012842f
C195 source.n96 a_n2018_n3288# 0.028668f
C196 source.n97 a_n2018_n3288# 0.028668f
C197 source.n98 a_n2018_n3288# 0.012842f
C198 source.n99 a_n2018_n3288# 0.012129f
C199 source.n100 a_n2018_n3288# 0.022571f
C200 source.n101 a_n2018_n3288# 0.022571f
C201 source.n102 a_n2018_n3288# 0.012129f
C202 source.n103 a_n2018_n3288# 0.012842f
C203 source.n104 a_n2018_n3288# 0.028668f
C204 source.n105 a_n2018_n3288# 0.028668f
C205 source.n106 a_n2018_n3288# 0.012842f
C206 source.n107 a_n2018_n3288# 0.012129f
C207 source.n108 a_n2018_n3288# 0.022571f
C208 source.n109 a_n2018_n3288# 0.022571f
C209 source.n110 a_n2018_n3288# 0.012129f
C210 source.n111 a_n2018_n3288# 0.012842f
C211 source.n112 a_n2018_n3288# 0.028668f
C212 source.n113 a_n2018_n3288# 0.028668f
C213 source.n114 a_n2018_n3288# 0.028668f
C214 source.n115 a_n2018_n3288# 0.012486f
C215 source.n116 a_n2018_n3288# 0.012129f
C216 source.n117 a_n2018_n3288# 0.022571f
C217 source.n118 a_n2018_n3288# 0.022571f
C218 source.n119 a_n2018_n3288# 0.012129f
C219 source.n120 a_n2018_n3288# 0.012842f
C220 source.n121 a_n2018_n3288# 0.028668f
C221 source.n122 a_n2018_n3288# 0.028668f
C222 source.n123 a_n2018_n3288# 0.012842f
C223 source.n124 a_n2018_n3288# 0.012129f
C224 source.n125 a_n2018_n3288# 0.022571f
C225 source.n126 a_n2018_n3288# 0.022571f
C226 source.n127 a_n2018_n3288# 0.012129f
C227 source.n128 a_n2018_n3288# 0.012842f
C228 source.n129 a_n2018_n3288# 0.028668f
C229 source.n130 a_n2018_n3288# 0.05883f
C230 source.n131 a_n2018_n3288# 0.012842f
C231 source.n132 a_n2018_n3288# 0.012129f
C232 source.n133 a_n2018_n3288# 0.048472f
C233 source.n134 a_n2018_n3288# 0.032468f
C234 source.n135 a_n2018_n3288# 0.109673f
C235 source.n136 a_n2018_n3288# 0.029898f
C236 source.n137 a_n2018_n3288# 0.022571f
C237 source.n138 a_n2018_n3288# 0.012129f
C238 source.n139 a_n2018_n3288# 0.028668f
C239 source.n140 a_n2018_n3288# 0.012842f
C240 source.n141 a_n2018_n3288# 0.022571f
C241 source.n142 a_n2018_n3288# 0.012129f
C242 source.n143 a_n2018_n3288# 0.028668f
C243 source.n144 a_n2018_n3288# 0.012842f
C244 source.n145 a_n2018_n3288# 0.022571f
C245 source.n146 a_n2018_n3288# 0.012486f
C246 source.n147 a_n2018_n3288# 0.028668f
C247 source.n148 a_n2018_n3288# 0.012129f
C248 source.n149 a_n2018_n3288# 0.012842f
C249 source.n150 a_n2018_n3288# 0.022571f
C250 source.n151 a_n2018_n3288# 0.012129f
C251 source.n152 a_n2018_n3288# 0.028668f
C252 source.n153 a_n2018_n3288# 0.012842f
C253 source.n154 a_n2018_n3288# 0.022571f
C254 source.n155 a_n2018_n3288# 0.012129f
C255 source.n156 a_n2018_n3288# 0.021501f
C256 source.n157 a_n2018_n3288# 0.020266f
C257 source.t8 a_n2018_n3288# 0.048418f
C258 source.n158 a_n2018_n3288# 0.162736f
C259 source.n159 a_n2018_n3288# 1.13868f
C260 source.n160 a_n2018_n3288# 0.012129f
C261 source.n161 a_n2018_n3288# 0.012842f
C262 source.n162 a_n2018_n3288# 0.028668f
C263 source.n163 a_n2018_n3288# 0.028668f
C264 source.n164 a_n2018_n3288# 0.012842f
C265 source.n165 a_n2018_n3288# 0.012129f
C266 source.n166 a_n2018_n3288# 0.022571f
C267 source.n167 a_n2018_n3288# 0.022571f
C268 source.n168 a_n2018_n3288# 0.012129f
C269 source.n169 a_n2018_n3288# 0.012842f
C270 source.n170 a_n2018_n3288# 0.028668f
C271 source.n171 a_n2018_n3288# 0.028668f
C272 source.n172 a_n2018_n3288# 0.012842f
C273 source.n173 a_n2018_n3288# 0.012129f
C274 source.n174 a_n2018_n3288# 0.022571f
C275 source.n175 a_n2018_n3288# 0.022571f
C276 source.n176 a_n2018_n3288# 0.012129f
C277 source.n177 a_n2018_n3288# 0.012842f
C278 source.n178 a_n2018_n3288# 0.028668f
C279 source.n179 a_n2018_n3288# 0.028668f
C280 source.n180 a_n2018_n3288# 0.028668f
C281 source.n181 a_n2018_n3288# 0.012486f
C282 source.n182 a_n2018_n3288# 0.012129f
C283 source.n183 a_n2018_n3288# 0.022571f
C284 source.n184 a_n2018_n3288# 0.022571f
C285 source.n185 a_n2018_n3288# 0.012129f
C286 source.n186 a_n2018_n3288# 0.012842f
C287 source.n187 a_n2018_n3288# 0.028668f
C288 source.n188 a_n2018_n3288# 0.028668f
C289 source.n189 a_n2018_n3288# 0.012842f
C290 source.n190 a_n2018_n3288# 0.012129f
C291 source.n191 a_n2018_n3288# 0.022571f
C292 source.n192 a_n2018_n3288# 0.022571f
C293 source.n193 a_n2018_n3288# 0.012129f
C294 source.n194 a_n2018_n3288# 0.012842f
C295 source.n195 a_n2018_n3288# 0.028668f
C296 source.n196 a_n2018_n3288# 0.05883f
C297 source.n197 a_n2018_n3288# 0.012842f
C298 source.n198 a_n2018_n3288# 0.012129f
C299 source.n199 a_n2018_n3288# 0.048472f
C300 source.n200 a_n2018_n3288# 0.032468f
C301 source.n201 a_n2018_n3288# 0.109673f
C302 source.t14 a_n2018_n3288# 0.214038f
C303 source.t18 a_n2018_n3288# 0.214038f
C304 source.n202 a_n2018_n3288# 1.83259f
C305 source.n203 a_n2018_n3288# 0.34738f
C306 source.t19 a_n2018_n3288# 0.214038f
C307 source.t16 a_n2018_n3288# 0.214038f
C308 source.n204 a_n2018_n3288# 1.83259f
C309 source.n205 a_n2018_n3288# 0.34738f
C310 source.n206 a_n2018_n3288# 0.029898f
C311 source.n207 a_n2018_n3288# 0.022571f
C312 source.n208 a_n2018_n3288# 0.012129f
C313 source.n209 a_n2018_n3288# 0.028668f
C314 source.n210 a_n2018_n3288# 0.012842f
C315 source.n211 a_n2018_n3288# 0.022571f
C316 source.n212 a_n2018_n3288# 0.012129f
C317 source.n213 a_n2018_n3288# 0.028668f
C318 source.n214 a_n2018_n3288# 0.012842f
C319 source.n215 a_n2018_n3288# 0.022571f
C320 source.n216 a_n2018_n3288# 0.012486f
C321 source.n217 a_n2018_n3288# 0.028668f
C322 source.n218 a_n2018_n3288# 0.012129f
C323 source.n219 a_n2018_n3288# 0.012842f
C324 source.n220 a_n2018_n3288# 0.022571f
C325 source.n221 a_n2018_n3288# 0.012129f
C326 source.n222 a_n2018_n3288# 0.028668f
C327 source.n223 a_n2018_n3288# 0.012842f
C328 source.n224 a_n2018_n3288# 0.022571f
C329 source.n225 a_n2018_n3288# 0.012129f
C330 source.n226 a_n2018_n3288# 0.021501f
C331 source.n227 a_n2018_n3288# 0.020266f
C332 source.t11 a_n2018_n3288# 0.048418f
C333 source.n228 a_n2018_n3288# 0.162736f
C334 source.n229 a_n2018_n3288# 1.13868f
C335 source.n230 a_n2018_n3288# 0.012129f
C336 source.n231 a_n2018_n3288# 0.012842f
C337 source.n232 a_n2018_n3288# 0.028668f
C338 source.n233 a_n2018_n3288# 0.028668f
C339 source.n234 a_n2018_n3288# 0.012842f
C340 source.n235 a_n2018_n3288# 0.012129f
C341 source.n236 a_n2018_n3288# 0.022571f
C342 source.n237 a_n2018_n3288# 0.022571f
C343 source.n238 a_n2018_n3288# 0.012129f
C344 source.n239 a_n2018_n3288# 0.012842f
C345 source.n240 a_n2018_n3288# 0.028668f
C346 source.n241 a_n2018_n3288# 0.028668f
C347 source.n242 a_n2018_n3288# 0.012842f
C348 source.n243 a_n2018_n3288# 0.012129f
C349 source.n244 a_n2018_n3288# 0.022571f
C350 source.n245 a_n2018_n3288# 0.022571f
C351 source.n246 a_n2018_n3288# 0.012129f
C352 source.n247 a_n2018_n3288# 0.012842f
C353 source.n248 a_n2018_n3288# 0.028668f
C354 source.n249 a_n2018_n3288# 0.028668f
C355 source.n250 a_n2018_n3288# 0.028668f
C356 source.n251 a_n2018_n3288# 0.012486f
C357 source.n252 a_n2018_n3288# 0.012129f
C358 source.n253 a_n2018_n3288# 0.022571f
C359 source.n254 a_n2018_n3288# 0.022571f
C360 source.n255 a_n2018_n3288# 0.012129f
C361 source.n256 a_n2018_n3288# 0.012842f
C362 source.n257 a_n2018_n3288# 0.028668f
C363 source.n258 a_n2018_n3288# 0.028668f
C364 source.n259 a_n2018_n3288# 0.012842f
C365 source.n260 a_n2018_n3288# 0.012129f
C366 source.n261 a_n2018_n3288# 0.022571f
C367 source.n262 a_n2018_n3288# 0.022571f
C368 source.n263 a_n2018_n3288# 0.012129f
C369 source.n264 a_n2018_n3288# 0.012842f
C370 source.n265 a_n2018_n3288# 0.028668f
C371 source.n266 a_n2018_n3288# 0.05883f
C372 source.n267 a_n2018_n3288# 0.012842f
C373 source.n268 a_n2018_n3288# 0.012129f
C374 source.n269 a_n2018_n3288# 0.048472f
C375 source.n270 a_n2018_n3288# 0.032468f
C376 source.n271 a_n2018_n3288# 1.30091f
C377 source.n272 a_n2018_n3288# 0.029898f
C378 source.n273 a_n2018_n3288# 0.022571f
C379 source.n274 a_n2018_n3288# 0.012129f
C380 source.n275 a_n2018_n3288# 0.028668f
C381 source.n276 a_n2018_n3288# 0.012842f
C382 source.n277 a_n2018_n3288# 0.022571f
C383 source.n278 a_n2018_n3288# 0.012129f
C384 source.n279 a_n2018_n3288# 0.028668f
C385 source.n280 a_n2018_n3288# 0.012842f
C386 source.n281 a_n2018_n3288# 0.022571f
C387 source.n282 a_n2018_n3288# 0.012486f
C388 source.n283 a_n2018_n3288# 0.028668f
C389 source.n284 a_n2018_n3288# 0.012842f
C390 source.n285 a_n2018_n3288# 0.022571f
C391 source.n286 a_n2018_n3288# 0.012129f
C392 source.n287 a_n2018_n3288# 0.028668f
C393 source.n288 a_n2018_n3288# 0.012842f
C394 source.n289 a_n2018_n3288# 0.022571f
C395 source.n290 a_n2018_n3288# 0.012129f
C396 source.n291 a_n2018_n3288# 0.021501f
C397 source.n292 a_n2018_n3288# 0.020266f
C398 source.t6 a_n2018_n3288# 0.048418f
C399 source.n293 a_n2018_n3288# 0.162736f
C400 source.n294 a_n2018_n3288# 1.13868f
C401 source.n295 a_n2018_n3288# 0.012129f
C402 source.n296 a_n2018_n3288# 0.012842f
C403 source.n297 a_n2018_n3288# 0.028668f
C404 source.n298 a_n2018_n3288# 0.028668f
C405 source.n299 a_n2018_n3288# 0.012842f
C406 source.n300 a_n2018_n3288# 0.012129f
C407 source.n301 a_n2018_n3288# 0.022571f
C408 source.n302 a_n2018_n3288# 0.022571f
C409 source.n303 a_n2018_n3288# 0.012129f
C410 source.n304 a_n2018_n3288# 0.012842f
C411 source.n305 a_n2018_n3288# 0.028668f
C412 source.n306 a_n2018_n3288# 0.028668f
C413 source.n307 a_n2018_n3288# 0.012842f
C414 source.n308 a_n2018_n3288# 0.012129f
C415 source.n309 a_n2018_n3288# 0.022571f
C416 source.n310 a_n2018_n3288# 0.022571f
C417 source.n311 a_n2018_n3288# 0.012129f
C418 source.n312 a_n2018_n3288# 0.012129f
C419 source.n313 a_n2018_n3288# 0.012842f
C420 source.n314 a_n2018_n3288# 0.028668f
C421 source.n315 a_n2018_n3288# 0.028668f
C422 source.n316 a_n2018_n3288# 0.028668f
C423 source.n317 a_n2018_n3288# 0.012486f
C424 source.n318 a_n2018_n3288# 0.012129f
C425 source.n319 a_n2018_n3288# 0.022571f
C426 source.n320 a_n2018_n3288# 0.022571f
C427 source.n321 a_n2018_n3288# 0.012129f
C428 source.n322 a_n2018_n3288# 0.012842f
C429 source.n323 a_n2018_n3288# 0.028668f
C430 source.n324 a_n2018_n3288# 0.028668f
C431 source.n325 a_n2018_n3288# 0.012842f
C432 source.n326 a_n2018_n3288# 0.012129f
C433 source.n327 a_n2018_n3288# 0.022571f
C434 source.n328 a_n2018_n3288# 0.022571f
C435 source.n329 a_n2018_n3288# 0.012129f
C436 source.n330 a_n2018_n3288# 0.012842f
C437 source.n331 a_n2018_n3288# 0.028668f
C438 source.n332 a_n2018_n3288# 0.05883f
C439 source.n333 a_n2018_n3288# 0.012842f
C440 source.n334 a_n2018_n3288# 0.012129f
C441 source.n335 a_n2018_n3288# 0.048472f
C442 source.n336 a_n2018_n3288# 0.032468f
C443 source.n337 a_n2018_n3288# 1.30091f
C444 source.t4 a_n2018_n3288# 0.214038f
C445 source.t7 a_n2018_n3288# 0.214038f
C446 source.n338 a_n2018_n3288# 1.83258f
C447 source.n339 a_n2018_n3288# 0.347391f
C448 source.t1 a_n2018_n3288# 0.214038f
C449 source.t20 a_n2018_n3288# 0.214038f
C450 source.n340 a_n2018_n3288# 1.83258f
C451 source.n341 a_n2018_n3288# 0.347391f
C452 source.n342 a_n2018_n3288# 0.029898f
C453 source.n343 a_n2018_n3288# 0.022571f
C454 source.n344 a_n2018_n3288# 0.012129f
C455 source.n345 a_n2018_n3288# 0.028668f
C456 source.n346 a_n2018_n3288# 0.012842f
C457 source.n347 a_n2018_n3288# 0.022571f
C458 source.n348 a_n2018_n3288# 0.012129f
C459 source.n349 a_n2018_n3288# 0.028668f
C460 source.n350 a_n2018_n3288# 0.012842f
C461 source.n351 a_n2018_n3288# 0.022571f
C462 source.n352 a_n2018_n3288# 0.012486f
C463 source.n353 a_n2018_n3288# 0.028668f
C464 source.n354 a_n2018_n3288# 0.012842f
C465 source.n355 a_n2018_n3288# 0.022571f
C466 source.n356 a_n2018_n3288# 0.012129f
C467 source.n357 a_n2018_n3288# 0.028668f
C468 source.n358 a_n2018_n3288# 0.012842f
C469 source.n359 a_n2018_n3288# 0.022571f
C470 source.n360 a_n2018_n3288# 0.012129f
C471 source.n361 a_n2018_n3288# 0.021501f
C472 source.n362 a_n2018_n3288# 0.020266f
C473 source.t5 a_n2018_n3288# 0.048418f
C474 source.n363 a_n2018_n3288# 0.162736f
C475 source.n364 a_n2018_n3288# 1.13868f
C476 source.n365 a_n2018_n3288# 0.012129f
C477 source.n366 a_n2018_n3288# 0.012842f
C478 source.n367 a_n2018_n3288# 0.028668f
C479 source.n368 a_n2018_n3288# 0.028668f
C480 source.n369 a_n2018_n3288# 0.012842f
C481 source.n370 a_n2018_n3288# 0.012129f
C482 source.n371 a_n2018_n3288# 0.022571f
C483 source.n372 a_n2018_n3288# 0.022571f
C484 source.n373 a_n2018_n3288# 0.012129f
C485 source.n374 a_n2018_n3288# 0.012842f
C486 source.n375 a_n2018_n3288# 0.028668f
C487 source.n376 a_n2018_n3288# 0.028668f
C488 source.n377 a_n2018_n3288# 0.012842f
C489 source.n378 a_n2018_n3288# 0.012129f
C490 source.n379 a_n2018_n3288# 0.022571f
C491 source.n380 a_n2018_n3288# 0.022571f
C492 source.n381 a_n2018_n3288# 0.012129f
C493 source.n382 a_n2018_n3288# 0.012129f
C494 source.n383 a_n2018_n3288# 0.012842f
C495 source.n384 a_n2018_n3288# 0.028668f
C496 source.n385 a_n2018_n3288# 0.028668f
C497 source.n386 a_n2018_n3288# 0.028668f
C498 source.n387 a_n2018_n3288# 0.012486f
C499 source.n388 a_n2018_n3288# 0.012129f
C500 source.n389 a_n2018_n3288# 0.022571f
C501 source.n390 a_n2018_n3288# 0.022571f
C502 source.n391 a_n2018_n3288# 0.012129f
C503 source.n392 a_n2018_n3288# 0.012842f
C504 source.n393 a_n2018_n3288# 0.028668f
C505 source.n394 a_n2018_n3288# 0.028668f
C506 source.n395 a_n2018_n3288# 0.012842f
C507 source.n396 a_n2018_n3288# 0.012129f
C508 source.n397 a_n2018_n3288# 0.022571f
C509 source.n398 a_n2018_n3288# 0.022571f
C510 source.n399 a_n2018_n3288# 0.012129f
C511 source.n400 a_n2018_n3288# 0.012842f
C512 source.n401 a_n2018_n3288# 0.028668f
C513 source.n402 a_n2018_n3288# 0.05883f
C514 source.n403 a_n2018_n3288# 0.012842f
C515 source.n404 a_n2018_n3288# 0.012129f
C516 source.n405 a_n2018_n3288# 0.048472f
C517 source.n406 a_n2018_n3288# 0.032468f
C518 source.n407 a_n2018_n3288# 0.109673f
C519 source.n408 a_n2018_n3288# 0.029898f
C520 source.n409 a_n2018_n3288# 0.022571f
C521 source.n410 a_n2018_n3288# 0.012129f
C522 source.n411 a_n2018_n3288# 0.028668f
C523 source.n412 a_n2018_n3288# 0.012842f
C524 source.n413 a_n2018_n3288# 0.022571f
C525 source.n414 a_n2018_n3288# 0.012129f
C526 source.n415 a_n2018_n3288# 0.028668f
C527 source.n416 a_n2018_n3288# 0.012842f
C528 source.n417 a_n2018_n3288# 0.022571f
C529 source.n418 a_n2018_n3288# 0.012486f
C530 source.n419 a_n2018_n3288# 0.028668f
C531 source.n420 a_n2018_n3288# 0.012842f
C532 source.n421 a_n2018_n3288# 0.022571f
C533 source.n422 a_n2018_n3288# 0.012129f
C534 source.n423 a_n2018_n3288# 0.028668f
C535 source.n424 a_n2018_n3288# 0.012842f
C536 source.n425 a_n2018_n3288# 0.022571f
C537 source.n426 a_n2018_n3288# 0.012129f
C538 source.n427 a_n2018_n3288# 0.021501f
C539 source.n428 a_n2018_n3288# 0.020266f
C540 source.t12 a_n2018_n3288# 0.048418f
C541 source.n429 a_n2018_n3288# 0.162736f
C542 source.n430 a_n2018_n3288# 1.13868f
C543 source.n431 a_n2018_n3288# 0.012129f
C544 source.n432 a_n2018_n3288# 0.012842f
C545 source.n433 a_n2018_n3288# 0.028668f
C546 source.n434 a_n2018_n3288# 0.028668f
C547 source.n435 a_n2018_n3288# 0.012842f
C548 source.n436 a_n2018_n3288# 0.012129f
C549 source.n437 a_n2018_n3288# 0.022571f
C550 source.n438 a_n2018_n3288# 0.022571f
C551 source.n439 a_n2018_n3288# 0.012129f
C552 source.n440 a_n2018_n3288# 0.012842f
C553 source.n441 a_n2018_n3288# 0.028668f
C554 source.n442 a_n2018_n3288# 0.028668f
C555 source.n443 a_n2018_n3288# 0.012842f
C556 source.n444 a_n2018_n3288# 0.012129f
C557 source.n445 a_n2018_n3288# 0.022571f
C558 source.n446 a_n2018_n3288# 0.022571f
C559 source.n447 a_n2018_n3288# 0.012129f
C560 source.n448 a_n2018_n3288# 0.012129f
C561 source.n449 a_n2018_n3288# 0.012842f
C562 source.n450 a_n2018_n3288# 0.028668f
C563 source.n451 a_n2018_n3288# 0.028668f
C564 source.n452 a_n2018_n3288# 0.028668f
C565 source.n453 a_n2018_n3288# 0.012486f
C566 source.n454 a_n2018_n3288# 0.012129f
C567 source.n455 a_n2018_n3288# 0.022571f
C568 source.n456 a_n2018_n3288# 0.022571f
C569 source.n457 a_n2018_n3288# 0.012129f
C570 source.n458 a_n2018_n3288# 0.012842f
C571 source.n459 a_n2018_n3288# 0.028668f
C572 source.n460 a_n2018_n3288# 0.028668f
C573 source.n461 a_n2018_n3288# 0.012842f
C574 source.n462 a_n2018_n3288# 0.012129f
C575 source.n463 a_n2018_n3288# 0.022571f
C576 source.n464 a_n2018_n3288# 0.022571f
C577 source.n465 a_n2018_n3288# 0.012129f
C578 source.n466 a_n2018_n3288# 0.012842f
C579 source.n467 a_n2018_n3288# 0.028668f
C580 source.n468 a_n2018_n3288# 0.05883f
C581 source.n469 a_n2018_n3288# 0.012842f
C582 source.n470 a_n2018_n3288# 0.012129f
C583 source.n471 a_n2018_n3288# 0.048472f
C584 source.n472 a_n2018_n3288# 0.032468f
C585 source.n473 a_n2018_n3288# 0.109673f
C586 source.t10 a_n2018_n3288# 0.214038f
C587 source.t15 a_n2018_n3288# 0.214038f
C588 source.n474 a_n2018_n3288# 1.83258f
C589 source.n475 a_n2018_n3288# 0.347391f
C590 source.t9 a_n2018_n3288# 0.214038f
C591 source.t13 a_n2018_n3288# 0.214038f
C592 source.n476 a_n2018_n3288# 1.83258f
C593 source.n477 a_n2018_n3288# 0.347391f
C594 source.n478 a_n2018_n3288# 0.029898f
C595 source.n479 a_n2018_n3288# 0.022571f
C596 source.n480 a_n2018_n3288# 0.012129f
C597 source.n481 a_n2018_n3288# 0.028668f
C598 source.n482 a_n2018_n3288# 0.012842f
C599 source.n483 a_n2018_n3288# 0.022571f
C600 source.n484 a_n2018_n3288# 0.012129f
C601 source.n485 a_n2018_n3288# 0.028668f
C602 source.n486 a_n2018_n3288# 0.012842f
C603 source.n487 a_n2018_n3288# 0.022571f
C604 source.n488 a_n2018_n3288# 0.012486f
C605 source.n489 a_n2018_n3288# 0.028668f
C606 source.n490 a_n2018_n3288# 0.012842f
C607 source.n491 a_n2018_n3288# 0.022571f
C608 source.n492 a_n2018_n3288# 0.012129f
C609 source.n493 a_n2018_n3288# 0.028668f
C610 source.n494 a_n2018_n3288# 0.012842f
C611 source.n495 a_n2018_n3288# 0.022571f
C612 source.n496 a_n2018_n3288# 0.012129f
C613 source.n497 a_n2018_n3288# 0.021501f
C614 source.n498 a_n2018_n3288# 0.020266f
C615 source.t17 a_n2018_n3288# 0.048418f
C616 source.n499 a_n2018_n3288# 0.162736f
C617 source.n500 a_n2018_n3288# 1.13868f
C618 source.n501 a_n2018_n3288# 0.012129f
C619 source.n502 a_n2018_n3288# 0.012842f
C620 source.n503 a_n2018_n3288# 0.028668f
C621 source.n504 a_n2018_n3288# 0.028668f
C622 source.n505 a_n2018_n3288# 0.012842f
C623 source.n506 a_n2018_n3288# 0.012129f
C624 source.n507 a_n2018_n3288# 0.022571f
C625 source.n508 a_n2018_n3288# 0.022571f
C626 source.n509 a_n2018_n3288# 0.012129f
C627 source.n510 a_n2018_n3288# 0.012842f
C628 source.n511 a_n2018_n3288# 0.028668f
C629 source.n512 a_n2018_n3288# 0.028668f
C630 source.n513 a_n2018_n3288# 0.012842f
C631 source.n514 a_n2018_n3288# 0.012129f
C632 source.n515 a_n2018_n3288# 0.022571f
C633 source.n516 a_n2018_n3288# 0.022571f
C634 source.n517 a_n2018_n3288# 0.012129f
C635 source.n518 a_n2018_n3288# 0.012129f
C636 source.n519 a_n2018_n3288# 0.012842f
C637 source.n520 a_n2018_n3288# 0.028668f
C638 source.n521 a_n2018_n3288# 0.028668f
C639 source.n522 a_n2018_n3288# 0.028668f
C640 source.n523 a_n2018_n3288# 0.012486f
C641 source.n524 a_n2018_n3288# 0.012129f
C642 source.n525 a_n2018_n3288# 0.022571f
C643 source.n526 a_n2018_n3288# 0.022571f
C644 source.n527 a_n2018_n3288# 0.012129f
C645 source.n528 a_n2018_n3288# 0.012842f
C646 source.n529 a_n2018_n3288# 0.028668f
C647 source.n530 a_n2018_n3288# 0.028668f
C648 source.n531 a_n2018_n3288# 0.012842f
C649 source.n532 a_n2018_n3288# 0.012129f
C650 source.n533 a_n2018_n3288# 0.022571f
C651 source.n534 a_n2018_n3288# 0.022571f
C652 source.n535 a_n2018_n3288# 0.012129f
C653 source.n536 a_n2018_n3288# 0.012842f
C654 source.n537 a_n2018_n3288# 0.028668f
C655 source.n538 a_n2018_n3288# 0.05883f
C656 source.n539 a_n2018_n3288# 0.012842f
C657 source.n540 a_n2018_n3288# 0.012129f
C658 source.n541 a_n2018_n3288# 0.048472f
C659 source.n542 a_n2018_n3288# 0.032468f
C660 source.n543 a_n2018_n3288# 0.251993f
C661 source.n544 a_n2018_n3288# 1.42667f
C662 minus.n0 a_n2018_n3288# 0.044128f
C663 minus.t6 a_n2018_n3288# 0.905989f
C664 minus.n1 a_n2018_n3288# 0.373469f
C665 minus.t3 a_n2018_n3288# 0.905989f
C666 minus.t10 a_n2018_n3288# 0.921876f
C667 minus.n2 a_n2018_n3288# 0.350459f
C668 minus.t9 a_n2018_n3288# 0.905989f
C669 minus.n3 a_n2018_n3288# 0.371858f
C670 minus.t7 a_n2018_n3288# 0.905989f
C671 minus.n4 a_n2018_n3288# 0.373469f
C672 minus.n5 a_n2018_n3288# 0.226163f
C673 minus.n6 a_n2018_n3288# 0.073501f
C674 minus.n7 a_n2018_n3288# 0.058883f
C675 minus.n8 a_n2018_n3288# 0.364952f
C676 minus.n9 a_n2018_n3288# 0.010014f
C677 minus.t4 a_n2018_n3288# 0.905989f
C678 minus.n10 a_n2018_n3288# 0.361959f
C679 minus.n11 a_n2018_n3288# 1.60691f
C680 minus.n12 a_n2018_n3288# 0.044128f
C681 minus.t11 a_n2018_n3288# 0.905989f
C682 minus.n13 a_n2018_n3288# 0.373469f
C683 minus.t8 a_n2018_n3288# 0.921876f
C684 minus.n14 a_n2018_n3288# 0.350459f
C685 minus.t2 a_n2018_n3288# 0.905989f
C686 minus.n15 a_n2018_n3288# 0.371858f
C687 minus.t5 a_n2018_n3288# 0.905989f
C688 minus.n16 a_n2018_n3288# 0.373469f
C689 minus.n17 a_n2018_n3288# 0.226163f
C690 minus.n18 a_n2018_n3288# 0.073501f
C691 minus.n19 a_n2018_n3288# 0.058883f
C692 minus.t1 a_n2018_n3288# 0.905989f
C693 minus.n20 a_n2018_n3288# 0.364952f
C694 minus.n21 a_n2018_n3288# 0.010014f
C695 minus.t0 a_n2018_n3288# 0.905989f
C696 minus.n22 a_n2018_n3288# 0.361959f
C697 minus.n23 a_n2018_n3288# 0.29757f
C698 minus.n24 a_n2018_n3288# 1.94519f
.ends

