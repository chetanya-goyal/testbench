* NGSPICE file created from diffpair47.ext - technology: sky130A

.subckt diffpair47 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t29 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X1 drain_right.t15 minus.t0 source.t1 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X2 source.t8 minus.t1 drain_right.t14 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X3 a_n2210_n1088# a_n2210_n1088# a_n2210_n1088# a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.5
X4 a_n2210_n1088# a_n2210_n1088# a_n2210_n1088# a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X5 source.t22 plus.t1 drain_left.t14 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X6 drain_right.t13 minus.t2 source.t0 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X7 a_n2210_n1088# a_n2210_n1088# a_n2210_n1088# a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X8 source.t30 plus.t2 drain_left.t13 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X9 drain_right.t12 minus.t3 source.t5 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X10 drain_right.t11 minus.t4 source.t15 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X11 source.t14 minus.t5 drain_right.t10 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X12 drain_left.t12 plus.t3 source.t31 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X13 drain_left.t11 plus.t4 source.t23 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X14 source.t7 minus.t6 drain_right.t9 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X15 source.t24 plus.t5 drain_left.t10 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X16 source.t6 minus.t7 drain_right.t8 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X17 drain_right.t7 minus.t8 source.t13 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X18 source.t11 minus.t9 drain_right.t6 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X19 drain_left.t9 plus.t6 source.t17 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X20 drain_right.t5 minus.t10 source.t10 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X21 drain_right.t4 minus.t11 source.t9 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X22 drain_right.t3 minus.t12 source.t2 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X23 a_n2210_n1088# a_n2210_n1088# a_n2210_n1088# a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.5
X24 drain_left.t8 plus.t7 source.t18 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X25 source.t21 plus.t8 drain_left.t7 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X26 source.t28 plus.t9 drain_left.t6 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X27 source.t4 minus.t13 drain_right.t2 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X28 source.t19 plus.t10 drain_left.t5 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X29 source.t26 plus.t11 drain_left.t4 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X30 source.t3 minus.t14 drain_right.t1 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X31 drain_left.t3 plus.t12 source.t25 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X32 drain_left.t2 plus.t13 source.t27 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X33 source.t16 plus.t14 drain_left.t1 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X34 source.t12 minus.t15 drain_right.t0 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X35 drain_left.t0 plus.t15 source.t20 a_n2210_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
R0 plus.n8 plus.n7 161.3
R1 plus.n9 plus.n4 161.3
R2 plus.n11 plus.n10 161.3
R3 plus.n12 plus.n3 161.3
R4 plus.n13 plus.n2 161.3
R5 plus.n15 plus.n14 161.3
R6 plus.n16 plus.n1 161.3
R7 plus.n18 plus.n17 161.3
R8 plus.n19 plus.n0 161.3
R9 plus.n21 plus.n20 161.3
R10 plus.n30 plus.n29 161.3
R11 plus.n31 plus.n26 161.3
R12 plus.n33 plus.n32 161.3
R13 plus.n34 plus.n25 161.3
R14 plus.n35 plus.n24 161.3
R15 plus.n37 plus.n36 161.3
R16 plus.n38 plus.n23 161.3
R17 plus.n40 plus.n39 161.3
R18 plus.n41 plus.n22 161.3
R19 plus.n43 plus.n42 161.3
R20 plus.n5 plus.t1 147.749
R21 plus.n27 plus.t6 147.749
R22 plus.n20 plus.t13 126.766
R23 plus.n19 plus.t5 126.766
R24 plus.n1 plus.t15 126.766
R25 plus.n13 plus.t11 126.766
R26 plus.n12 plus.t3 126.766
R27 plus.n4 plus.t14 126.766
R28 plus.n6 plus.t7 126.766
R29 plus.n42 plus.t2 126.766
R30 plus.n41 plus.t12 126.766
R31 plus.n23 plus.t9 126.766
R32 plus.n35 plus.t0 126.766
R33 plus.n34 plus.t10 126.766
R34 plus.n26 plus.t4 126.766
R35 plus.n28 plus.t8 126.766
R36 plus.n8 plus.n5 70.4033
R37 plus.n30 plus.n27 70.4033
R38 plus.n20 plus.n19 48.2005
R39 plus.n13 plus.n12 48.2005
R40 plus.n42 plus.n41 48.2005
R41 plus.n35 plus.n34 48.2005
R42 plus.n18 plus.n1 37.246
R43 plus.n7 plus.n4 37.246
R44 plus.n40 plus.n23 37.246
R45 plus.n29 plus.n26 37.246
R46 plus.n14 plus.n1 35.7853
R47 plus.n11 plus.n4 35.7853
R48 plus.n36 plus.n23 35.7853
R49 plus.n33 plus.n26 35.7853
R50 plus plus.n43 27.268
R51 plus.n6 plus.n5 20.9576
R52 plus.n28 plus.n27 20.9576
R53 plus.n14 plus.n13 12.4157
R54 plus.n12 plus.n11 12.4157
R55 plus.n36 plus.n35 12.4157
R56 plus.n34 plus.n33 12.4157
R57 plus.n19 plus.n18 10.955
R58 plus.n7 plus.n6 10.955
R59 plus.n41 plus.n40 10.955
R60 plus.n29 plus.n28 10.955
R61 plus plus.n21 8.03838
R62 plus.n9 plus.n8 0.189894
R63 plus.n10 plus.n9 0.189894
R64 plus.n10 plus.n3 0.189894
R65 plus.n3 plus.n2 0.189894
R66 plus.n15 plus.n2 0.189894
R67 plus.n16 plus.n15 0.189894
R68 plus.n17 plus.n16 0.189894
R69 plus.n17 plus.n0 0.189894
R70 plus.n21 plus.n0 0.189894
R71 plus.n43 plus.n22 0.189894
R72 plus.n39 plus.n22 0.189894
R73 plus.n39 plus.n38 0.189894
R74 plus.n38 plus.n37 0.189894
R75 plus.n37 plus.n24 0.189894
R76 plus.n25 plus.n24 0.189894
R77 plus.n32 plus.n25 0.189894
R78 plus.n32 plus.n31 0.189894
R79 plus.n31 plus.n30 0.189894
R80 source.n0 source.t27 243.255
R81 source.n7 source.t22 243.255
R82 source.n8 source.t10 243.255
R83 source.n15 source.t11 243.255
R84 source.n31 source.t5 243.254
R85 source.n24 source.t7 243.254
R86 source.n23 source.t17 243.254
R87 source.n16 source.t30 243.254
R88 source.n2 source.n1 223.454
R89 source.n4 source.n3 223.454
R90 source.n6 source.n5 223.454
R91 source.n10 source.n9 223.454
R92 source.n12 source.n11 223.454
R93 source.n14 source.n13 223.454
R94 source.n30 source.n29 223.453
R95 source.n28 source.n27 223.453
R96 source.n26 source.n25 223.453
R97 source.n22 source.n21 223.453
R98 source.n20 source.n19 223.453
R99 source.n18 source.n17 223.453
R100 source.n29 source.t2 19.8005
R101 source.n29 source.t3 19.8005
R102 source.n27 source.t13 19.8005
R103 source.n27 source.t12 19.8005
R104 source.n25 source.t9 19.8005
R105 source.n25 source.t14 19.8005
R106 source.n21 source.t23 19.8005
R107 source.n21 source.t21 19.8005
R108 source.n19 source.t29 19.8005
R109 source.n19 source.t19 19.8005
R110 source.n17 source.t25 19.8005
R111 source.n17 source.t28 19.8005
R112 source.n1 source.t20 19.8005
R113 source.n1 source.t24 19.8005
R114 source.n3 source.t31 19.8005
R115 source.n3 source.t26 19.8005
R116 source.n5 source.t18 19.8005
R117 source.n5 source.t16 19.8005
R118 source.n9 source.t15 19.8005
R119 source.n9 source.t8 19.8005
R120 source.n11 source.t0 19.8005
R121 source.n11 source.t4 19.8005
R122 source.n13 source.t1 19.8005
R123 source.n13 source.t6 19.8005
R124 source.n16 source.n15 13.6699
R125 source.n32 source.n0 8.04922
R126 source.n32 source.n31 5.62119
R127 source.n15 source.n14 0.716017
R128 source.n14 source.n12 0.716017
R129 source.n12 source.n10 0.716017
R130 source.n10 source.n8 0.716017
R131 source.n7 source.n6 0.716017
R132 source.n6 source.n4 0.716017
R133 source.n4 source.n2 0.716017
R134 source.n2 source.n0 0.716017
R135 source.n18 source.n16 0.716017
R136 source.n20 source.n18 0.716017
R137 source.n22 source.n20 0.716017
R138 source.n23 source.n22 0.716017
R139 source.n26 source.n24 0.716017
R140 source.n28 source.n26 0.716017
R141 source.n30 source.n28 0.716017
R142 source.n31 source.n30 0.716017
R143 source.n8 source.n7 0.470328
R144 source.n24 source.n23 0.470328
R145 source source.n32 0.188
R146 drain_left.n9 drain_left.n7 240.849
R147 drain_left.n5 drain_left.n3 240.847
R148 drain_left.n2 drain_left.n0 240.847
R149 drain_left.n13 drain_left.n12 240.132
R150 drain_left.n11 drain_left.n10 240.132
R151 drain_left.n9 drain_left.n8 240.132
R152 drain_left.n5 drain_left.n4 240.131
R153 drain_left.n2 drain_left.n1 240.131
R154 drain_left drain_left.n6 23.6846
R155 drain_left.n3 drain_left.t7 19.8005
R156 drain_left.n3 drain_left.t9 19.8005
R157 drain_left.n4 drain_left.t5 19.8005
R158 drain_left.n4 drain_left.t11 19.8005
R159 drain_left.n1 drain_left.t6 19.8005
R160 drain_left.n1 drain_left.t15 19.8005
R161 drain_left.n0 drain_left.t13 19.8005
R162 drain_left.n0 drain_left.t3 19.8005
R163 drain_left.n12 drain_left.t10 19.8005
R164 drain_left.n12 drain_left.t2 19.8005
R165 drain_left.n10 drain_left.t4 19.8005
R166 drain_left.n10 drain_left.t0 19.8005
R167 drain_left.n8 drain_left.t1 19.8005
R168 drain_left.n8 drain_left.t12 19.8005
R169 drain_left.n7 drain_left.t14 19.8005
R170 drain_left.n7 drain_left.t8 19.8005
R171 drain_left drain_left.n13 6.36873
R172 drain_left.n11 drain_left.n9 0.716017
R173 drain_left.n13 drain_left.n11 0.716017
R174 drain_left.n6 drain_left.n5 0.302913
R175 drain_left.n6 drain_left.n2 0.302913
R176 minus.n21 minus.n20 161.3
R177 minus.n19 minus.n0 161.3
R178 minus.n18 minus.n17 161.3
R179 minus.n16 minus.n1 161.3
R180 minus.n15 minus.n14 161.3
R181 minus.n13 minus.n2 161.3
R182 minus.n12 minus.n11 161.3
R183 minus.n10 minus.n3 161.3
R184 minus.n9 minus.n8 161.3
R185 minus.n7 minus.n4 161.3
R186 minus.n43 minus.n42 161.3
R187 minus.n41 minus.n22 161.3
R188 minus.n40 minus.n39 161.3
R189 minus.n38 minus.n23 161.3
R190 minus.n37 minus.n36 161.3
R191 minus.n35 minus.n24 161.3
R192 minus.n34 minus.n33 161.3
R193 minus.n32 minus.n25 161.3
R194 minus.n31 minus.n30 161.3
R195 minus.n29 minus.n26 161.3
R196 minus.n5 minus.t10 147.749
R197 minus.n27 minus.t6 147.749
R198 minus.n6 minus.t1 126.766
R199 minus.n8 minus.t4 126.766
R200 minus.n12 minus.t13 126.766
R201 minus.n13 minus.t2 126.766
R202 minus.n1 minus.t7 126.766
R203 minus.n19 minus.t0 126.766
R204 minus.n20 minus.t9 126.766
R205 minus.n28 minus.t11 126.766
R206 minus.n30 minus.t5 126.766
R207 minus.n34 minus.t8 126.766
R208 minus.n35 minus.t15 126.766
R209 minus.n23 minus.t12 126.766
R210 minus.n41 minus.t14 126.766
R211 minus.n42 minus.t3 126.766
R212 minus.n5 minus.n4 70.4033
R213 minus.n27 minus.n26 70.4033
R214 minus.n13 minus.n12 48.2005
R215 minus.n20 minus.n19 48.2005
R216 minus.n35 minus.n34 48.2005
R217 minus.n42 minus.n41 48.2005
R218 minus.n8 minus.n7 37.246
R219 minus.n18 minus.n1 37.246
R220 minus.n30 minus.n29 37.246
R221 minus.n40 minus.n23 37.246
R222 minus.n8 minus.n3 35.7853
R223 minus.n14 minus.n1 35.7853
R224 minus.n30 minus.n25 35.7853
R225 minus.n36 minus.n23 35.7853
R226 minus.n44 minus.n21 29.2202
R227 minus.n6 minus.n5 20.9576
R228 minus.n28 minus.n27 20.9576
R229 minus.n12 minus.n3 12.4157
R230 minus.n14 minus.n13 12.4157
R231 minus.n34 minus.n25 12.4157
R232 minus.n36 minus.n35 12.4157
R233 minus.n7 minus.n6 10.955
R234 minus.n19 minus.n18 10.955
R235 minus.n29 minus.n28 10.955
R236 minus.n41 minus.n40 10.955
R237 minus.n44 minus.n43 6.56111
R238 minus.n21 minus.n0 0.189894
R239 minus.n17 minus.n0 0.189894
R240 minus.n17 minus.n16 0.189894
R241 minus.n16 minus.n15 0.189894
R242 minus.n15 minus.n2 0.189894
R243 minus.n11 minus.n2 0.189894
R244 minus.n11 minus.n10 0.189894
R245 minus.n10 minus.n9 0.189894
R246 minus.n9 minus.n4 0.189894
R247 minus.n31 minus.n26 0.189894
R248 minus.n32 minus.n31 0.189894
R249 minus.n33 minus.n32 0.189894
R250 minus.n33 minus.n24 0.189894
R251 minus.n37 minus.n24 0.189894
R252 minus.n38 minus.n37 0.189894
R253 minus.n39 minus.n38 0.189894
R254 minus.n39 minus.n22 0.189894
R255 minus.n43 minus.n22 0.189894
R256 minus minus.n44 0.188
R257 drain_right.n9 drain_right.n7 240.849
R258 drain_right.n5 drain_right.n3 240.847
R259 drain_right.n2 drain_right.n0 240.847
R260 drain_right.n9 drain_right.n8 240.132
R261 drain_right.n11 drain_right.n10 240.132
R262 drain_right.n13 drain_right.n12 240.132
R263 drain_right.n5 drain_right.n4 240.131
R264 drain_right.n2 drain_right.n1 240.131
R265 drain_right drain_right.n6 23.1314
R266 drain_right.n3 drain_right.t1 19.8005
R267 drain_right.n3 drain_right.t12 19.8005
R268 drain_right.n4 drain_right.t0 19.8005
R269 drain_right.n4 drain_right.t3 19.8005
R270 drain_right.n1 drain_right.t10 19.8005
R271 drain_right.n1 drain_right.t7 19.8005
R272 drain_right.n0 drain_right.t9 19.8005
R273 drain_right.n0 drain_right.t4 19.8005
R274 drain_right.n7 drain_right.t14 19.8005
R275 drain_right.n7 drain_right.t5 19.8005
R276 drain_right.n8 drain_right.t2 19.8005
R277 drain_right.n8 drain_right.t11 19.8005
R278 drain_right.n10 drain_right.t8 19.8005
R279 drain_right.n10 drain_right.t13 19.8005
R280 drain_right.n12 drain_right.t6 19.8005
R281 drain_right.n12 drain_right.t15 19.8005
R282 drain_right drain_right.n13 6.36873
R283 drain_right.n13 drain_right.n11 0.716017
R284 drain_right.n11 drain_right.n9 0.716017
R285 drain_right.n6 drain_right.n5 0.302913
R286 drain_right.n6 drain_right.n2 0.302913
C0 source drain_left 4.81708f
C1 drain_right plus 0.381348f
C2 minus plus 3.8792f
C3 drain_right minus 1.20611f
C4 plus drain_left 1.42311f
C5 plus source 1.71413f
C6 drain_right drain_left 1.15077f
C7 drain_right source 4.81827f
C8 minus drain_left 0.17967f
C9 minus source 1.70027f
C10 drain_right a_n2210_n1088# 3.92803f
C11 drain_left a_n2210_n1088# 4.21111f
C12 source a_n2210_n1088# 2.632636f
C13 minus a_n2210_n1088# 7.828429f
C14 plus a_n2210_n1088# 8.451294f
C15 drain_right.t9 a_n2210_n1088# 0.017269f
C16 drain_right.t4 a_n2210_n1088# 0.017269f
C17 drain_right.n0 a_n2210_n1088# 0.067882f
C18 drain_right.t10 a_n2210_n1088# 0.017269f
C19 drain_right.t7 a_n2210_n1088# 0.017269f
C20 drain_right.n1 a_n2210_n1088# 0.067102f
C21 drain_right.n2 a_n2210_n1088# 0.487787f
C22 drain_right.t1 a_n2210_n1088# 0.017269f
C23 drain_right.t12 a_n2210_n1088# 0.017269f
C24 drain_right.n3 a_n2210_n1088# 0.067882f
C25 drain_right.t0 a_n2210_n1088# 0.017269f
C26 drain_right.t3 a_n2210_n1088# 0.017269f
C27 drain_right.n4 a_n2210_n1088# 0.067102f
C28 drain_right.n5 a_n2210_n1088# 0.487787f
C29 drain_right.n6 a_n2210_n1088# 0.633748f
C30 drain_right.t14 a_n2210_n1088# 0.017269f
C31 drain_right.t5 a_n2210_n1088# 0.017269f
C32 drain_right.n7 a_n2210_n1088# 0.067882f
C33 drain_right.t2 a_n2210_n1088# 0.017269f
C34 drain_right.t11 a_n2210_n1088# 0.017269f
C35 drain_right.n8 a_n2210_n1088# 0.067102f
C36 drain_right.n9 a_n2210_n1088# 0.5152f
C37 drain_right.t8 a_n2210_n1088# 0.017269f
C38 drain_right.t13 a_n2210_n1088# 0.017269f
C39 drain_right.n10 a_n2210_n1088# 0.067102f
C40 drain_right.n11 a_n2210_n1088# 0.253589f
C41 drain_right.t6 a_n2210_n1088# 0.017269f
C42 drain_right.t15 a_n2210_n1088# 0.017269f
C43 drain_right.n12 a_n2210_n1088# 0.067102f
C44 drain_right.n13 a_n2210_n1088# 0.441338f
C45 minus.n0 a_n2210_n1088# 0.027212f
C46 minus.t7 a_n2210_n1088# 0.046138f
C47 minus.n1 a_n2210_n1088# 0.050843f
C48 minus.n2 a_n2210_n1088# 0.027212f
C49 minus.n3 a_n2210_n1088# 0.006175f
C50 minus.t13 a_n2210_n1088# 0.046138f
C51 minus.n4 a_n2210_n1088# 0.086638f
C52 minus.t1 a_n2210_n1088# 0.046138f
C53 minus.t10 a_n2210_n1088# 0.052958f
C54 minus.n5 a_n2210_n1088# 0.041369f
C55 minus.n6 a_n2210_n1088# 0.04925f
C56 minus.n7 a_n2210_n1088# 0.006175f
C57 minus.t4 a_n2210_n1088# 0.046138f
C58 minus.n8 a_n2210_n1088# 0.050843f
C59 minus.n9 a_n2210_n1088# 0.027212f
C60 minus.n10 a_n2210_n1088# 0.027212f
C61 minus.n11 a_n2210_n1088# 0.027212f
C62 minus.n12 a_n2210_n1088# 0.049417f
C63 minus.t2 a_n2210_n1088# 0.046138f
C64 minus.n13 a_n2210_n1088# 0.049417f
C65 minus.n14 a_n2210_n1088# 0.006175f
C66 minus.n15 a_n2210_n1088# 0.027212f
C67 minus.n16 a_n2210_n1088# 0.027212f
C68 minus.n17 a_n2210_n1088# 0.027212f
C69 minus.n18 a_n2210_n1088# 0.006175f
C70 minus.t0 a_n2210_n1088# 0.046138f
C71 minus.n19 a_n2210_n1088# 0.04925f
C72 minus.t9 a_n2210_n1088# 0.046138f
C73 minus.n20 a_n2210_n1088# 0.047991f
C74 minus.n21 a_n2210_n1088# 0.67815f
C75 minus.n22 a_n2210_n1088# 0.027212f
C76 minus.t12 a_n2210_n1088# 0.046138f
C77 minus.n23 a_n2210_n1088# 0.050843f
C78 minus.n24 a_n2210_n1088# 0.027212f
C79 minus.n25 a_n2210_n1088# 0.006175f
C80 minus.n26 a_n2210_n1088# 0.086638f
C81 minus.t6 a_n2210_n1088# 0.052958f
C82 minus.n27 a_n2210_n1088# 0.041369f
C83 minus.t11 a_n2210_n1088# 0.046138f
C84 minus.n28 a_n2210_n1088# 0.04925f
C85 minus.n29 a_n2210_n1088# 0.006175f
C86 minus.t5 a_n2210_n1088# 0.046138f
C87 minus.n30 a_n2210_n1088# 0.050843f
C88 minus.n31 a_n2210_n1088# 0.027212f
C89 minus.n32 a_n2210_n1088# 0.027212f
C90 minus.n33 a_n2210_n1088# 0.027212f
C91 minus.t8 a_n2210_n1088# 0.046138f
C92 minus.n34 a_n2210_n1088# 0.049417f
C93 minus.t15 a_n2210_n1088# 0.046138f
C94 minus.n35 a_n2210_n1088# 0.049417f
C95 minus.n36 a_n2210_n1088# 0.006175f
C96 minus.n37 a_n2210_n1088# 0.027212f
C97 minus.n38 a_n2210_n1088# 0.027212f
C98 minus.n39 a_n2210_n1088# 0.027212f
C99 minus.n40 a_n2210_n1088# 0.006175f
C100 minus.t14 a_n2210_n1088# 0.046138f
C101 minus.n41 a_n2210_n1088# 0.04925f
C102 minus.t3 a_n2210_n1088# 0.046138f
C103 minus.n42 a_n2210_n1088# 0.047991f
C104 minus.n43 a_n2210_n1088# 0.181811f
C105 minus.n44 a_n2210_n1088# 0.835497f
C106 drain_left.t13 a_n2210_n1088# 0.016967f
C107 drain_left.t3 a_n2210_n1088# 0.016967f
C108 drain_left.n0 a_n2210_n1088# 0.066694f
C109 drain_left.t6 a_n2210_n1088# 0.016967f
C110 drain_left.t15 a_n2210_n1088# 0.016967f
C111 drain_left.n1 a_n2210_n1088# 0.065928f
C112 drain_left.n2 a_n2210_n1088# 0.479251f
C113 drain_left.t7 a_n2210_n1088# 0.016967f
C114 drain_left.t9 a_n2210_n1088# 0.016967f
C115 drain_left.n3 a_n2210_n1088# 0.066694f
C116 drain_left.t5 a_n2210_n1088# 0.016967f
C117 drain_left.t11 a_n2210_n1088# 0.016967f
C118 drain_left.n4 a_n2210_n1088# 0.065928f
C119 drain_left.n5 a_n2210_n1088# 0.479251f
C120 drain_left.n6 a_n2210_n1088# 0.664055f
C121 drain_left.t14 a_n2210_n1088# 0.016967f
C122 drain_left.t8 a_n2210_n1088# 0.016967f
C123 drain_left.n7 a_n2210_n1088# 0.066694f
C124 drain_left.t1 a_n2210_n1088# 0.016967f
C125 drain_left.t12 a_n2210_n1088# 0.016967f
C126 drain_left.n8 a_n2210_n1088# 0.065928f
C127 drain_left.n9 a_n2210_n1088# 0.506185f
C128 drain_left.t4 a_n2210_n1088# 0.016967f
C129 drain_left.t0 a_n2210_n1088# 0.016967f
C130 drain_left.n10 a_n2210_n1088# 0.065928f
C131 drain_left.n11 a_n2210_n1088# 0.249152f
C132 drain_left.t10 a_n2210_n1088# 0.016967f
C133 drain_left.t2 a_n2210_n1088# 0.016967f
C134 drain_left.n12 a_n2210_n1088# 0.065928f
C135 drain_left.n13 a_n2210_n1088# 0.433616f
C136 source.t27 a_n2210_n1088# 0.114274f
C137 source.n0 a_n2210_n1088# 0.516494f
C138 source.t20 a_n2210_n1088# 0.020531f
C139 source.t24 a_n2210_n1088# 0.020531f
C140 source.n1 a_n2210_n1088# 0.066586f
C141 source.n2 a_n2210_n1088# 0.279371f
C142 source.t31 a_n2210_n1088# 0.020531f
C143 source.t26 a_n2210_n1088# 0.020531f
C144 source.n3 a_n2210_n1088# 0.066586f
C145 source.n4 a_n2210_n1088# 0.279371f
C146 source.t18 a_n2210_n1088# 0.020531f
C147 source.t16 a_n2210_n1088# 0.020531f
C148 source.n5 a_n2210_n1088# 0.066586f
C149 source.n6 a_n2210_n1088# 0.279371f
C150 source.t22 a_n2210_n1088# 0.114274f
C151 source.n7 a_n2210_n1088# 0.267109f
C152 source.t10 a_n2210_n1088# 0.114274f
C153 source.n8 a_n2210_n1088# 0.267109f
C154 source.t15 a_n2210_n1088# 0.020531f
C155 source.t8 a_n2210_n1088# 0.020531f
C156 source.n9 a_n2210_n1088# 0.066586f
C157 source.n10 a_n2210_n1088# 0.279371f
C158 source.t0 a_n2210_n1088# 0.020531f
C159 source.t4 a_n2210_n1088# 0.020531f
C160 source.n11 a_n2210_n1088# 0.066586f
C161 source.n12 a_n2210_n1088# 0.279371f
C162 source.t1 a_n2210_n1088# 0.020531f
C163 source.t6 a_n2210_n1088# 0.020531f
C164 source.n13 a_n2210_n1088# 0.066586f
C165 source.n14 a_n2210_n1088# 0.279371f
C166 source.t11 a_n2210_n1088# 0.114274f
C167 source.n15 a_n2210_n1088# 0.72773f
C168 source.t30 a_n2210_n1088# 0.114274f
C169 source.n16 a_n2210_n1088# 0.72773f
C170 source.t25 a_n2210_n1088# 0.020531f
C171 source.t28 a_n2210_n1088# 0.020531f
C172 source.n17 a_n2210_n1088# 0.066586f
C173 source.n18 a_n2210_n1088# 0.279371f
C174 source.t29 a_n2210_n1088# 0.020531f
C175 source.t19 a_n2210_n1088# 0.020531f
C176 source.n19 a_n2210_n1088# 0.066586f
C177 source.n20 a_n2210_n1088# 0.279371f
C178 source.t23 a_n2210_n1088# 0.020531f
C179 source.t21 a_n2210_n1088# 0.020531f
C180 source.n21 a_n2210_n1088# 0.066586f
C181 source.n22 a_n2210_n1088# 0.279371f
C182 source.t17 a_n2210_n1088# 0.114274f
C183 source.n23 a_n2210_n1088# 0.267109f
C184 source.t7 a_n2210_n1088# 0.114274f
C185 source.n24 a_n2210_n1088# 0.267109f
C186 source.t9 a_n2210_n1088# 0.020531f
C187 source.t14 a_n2210_n1088# 0.020531f
C188 source.n25 a_n2210_n1088# 0.066586f
C189 source.n26 a_n2210_n1088# 0.279371f
C190 source.t13 a_n2210_n1088# 0.020531f
C191 source.t12 a_n2210_n1088# 0.020531f
C192 source.n27 a_n2210_n1088# 0.066586f
C193 source.n28 a_n2210_n1088# 0.279371f
C194 source.t2 a_n2210_n1088# 0.020531f
C195 source.t3 a_n2210_n1088# 0.020531f
C196 source.n29 a_n2210_n1088# 0.066586f
C197 source.n30 a_n2210_n1088# 0.279371f
C198 source.t5 a_n2210_n1088# 0.114274f
C199 source.n31 a_n2210_n1088# 0.425244f
C200 source.n32 a_n2210_n1088# 0.532202f
C201 plus.n0 a_n2210_n1088# 0.027601f
C202 plus.t13 a_n2210_n1088# 0.046798f
C203 plus.t5 a_n2210_n1088# 0.046798f
C204 plus.t15 a_n2210_n1088# 0.046798f
C205 plus.n1 a_n2210_n1088# 0.051571f
C206 plus.n2 a_n2210_n1088# 0.027601f
C207 plus.t11 a_n2210_n1088# 0.046798f
C208 plus.t3 a_n2210_n1088# 0.046798f
C209 plus.n3 a_n2210_n1088# 0.027601f
C210 plus.t14 a_n2210_n1088# 0.046798f
C211 plus.n4 a_n2210_n1088# 0.051571f
C212 plus.t1 a_n2210_n1088# 0.053716f
C213 plus.n5 a_n2210_n1088# 0.041961f
C214 plus.t7 a_n2210_n1088# 0.046798f
C215 plus.n6 a_n2210_n1088# 0.049954f
C216 plus.n7 a_n2210_n1088# 0.006263f
C217 plus.n8 a_n2210_n1088# 0.087879f
C218 plus.n9 a_n2210_n1088# 0.027601f
C219 plus.n10 a_n2210_n1088# 0.027601f
C220 plus.n11 a_n2210_n1088# 0.006263f
C221 plus.n12 a_n2210_n1088# 0.050125f
C222 plus.n13 a_n2210_n1088# 0.050125f
C223 plus.n14 a_n2210_n1088# 0.006263f
C224 plus.n15 a_n2210_n1088# 0.027601f
C225 plus.n16 a_n2210_n1088# 0.027601f
C226 plus.n17 a_n2210_n1088# 0.027601f
C227 plus.n18 a_n2210_n1088# 0.006263f
C228 plus.n19 a_n2210_n1088# 0.049954f
C229 plus.n20 a_n2210_n1088# 0.048678f
C230 plus.n21 a_n2210_n1088# 0.193411f
C231 plus.n22 a_n2210_n1088# 0.027601f
C232 plus.t2 a_n2210_n1088# 0.046798f
C233 plus.t12 a_n2210_n1088# 0.046798f
C234 plus.t9 a_n2210_n1088# 0.046798f
C235 plus.n23 a_n2210_n1088# 0.051571f
C236 plus.n24 a_n2210_n1088# 0.027601f
C237 plus.t0 a_n2210_n1088# 0.046798f
C238 plus.n25 a_n2210_n1088# 0.027601f
C239 plus.t10 a_n2210_n1088# 0.046798f
C240 plus.t4 a_n2210_n1088# 0.046798f
C241 plus.n26 a_n2210_n1088# 0.051571f
C242 plus.t6 a_n2210_n1088# 0.053716f
C243 plus.n27 a_n2210_n1088# 0.041961f
C244 plus.t8 a_n2210_n1088# 0.046798f
C245 plus.n28 a_n2210_n1088# 0.049954f
C246 plus.n29 a_n2210_n1088# 0.006263f
C247 plus.n30 a_n2210_n1088# 0.087879f
C248 plus.n31 a_n2210_n1088# 0.027601f
C249 plus.n32 a_n2210_n1088# 0.027601f
C250 plus.n33 a_n2210_n1088# 0.006263f
C251 plus.n34 a_n2210_n1088# 0.050125f
C252 plus.n35 a_n2210_n1088# 0.050125f
C253 plus.n36 a_n2210_n1088# 0.006263f
C254 plus.n37 a_n2210_n1088# 0.027601f
C255 plus.n38 a_n2210_n1088# 0.027601f
C256 plus.n39 a_n2210_n1088# 0.027601f
C257 plus.n40 a_n2210_n1088# 0.006263f
C258 plus.n41 a_n2210_n1088# 0.049954f
C259 plus.n42 a_n2210_n1088# 0.048678f
C260 plus.n43 a_n2210_n1088# 0.664915f
.ends

