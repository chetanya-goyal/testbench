* NGSPICE file created from diffpair635.ext - technology: sky130A

.subckt diffpair635 minus drain_right drain_left source plus
X0 drain_left.t11 plus.t0 source.t17 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X1 source.t7 minus.t0 drain_right.t11 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X2 source.t2 minus.t1 drain_right.t10 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X3 source.t21 plus.t1 drain_left.t10 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X4 a_n2298_n4888# a_n2298_n4888# a_n2298_n4888# a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.8
X5 drain_right.t9 minus.t2 source.t9 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X6 a_n2298_n4888# a_n2298_n4888# a_n2298_n4888# a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X7 drain_right.t8 minus.t3 source.t22 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X8 source.t13 plus.t2 drain_left.t9 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X9 drain_right.t7 minus.t4 source.t8 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X10 source.t0 minus.t5 drain_right.t6 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X11 source.t16 plus.t3 drain_left.t8 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X12 drain_right.t5 minus.t6 source.t23 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X13 drain_right.t4 minus.t7 source.t3 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X14 source.t1 minus.t8 drain_right.t3 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X15 source.t4 minus.t9 drain_right.t2 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X16 drain_right.t1 minus.t10 source.t6 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X17 drain_left.t7 plus.t4 source.t12 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X18 drain_left.t6 plus.t5 source.t15 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X19 source.t11 plus.t6 drain_left.t5 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X20 a_n2298_n4888# a_n2298_n4888# a_n2298_n4888# a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X21 drain_left.t4 plus.t7 source.t20 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X22 drain_left.t3 plus.t8 source.t19 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X23 source.t18 plus.t9 drain_left.t2 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X24 drain_left.t1 plus.t10 source.t14 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X25 source.t5 minus.t11 drain_right.t0 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X26 a_n2298_n4888# a_n2298_n4888# a_n2298_n4888# a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X27 source.t10 plus.t11 drain_left.t0 a_n2298_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
R0 plus.n4 plus.t11 673
R1 plus.n20 plus.t0 673
R2 plus.n14 plus.t4 651.605
R3 plus.n12 plus.t9 651.605
R4 plus.n2 plus.t5 651.605
R5 plus.n7 plus.t6 651.605
R6 plus.n5 plus.t10 651.605
R7 plus.n30 plus.t1 651.605
R8 plus.n28 plus.t7 651.605
R9 plus.n18 plus.t2 651.605
R10 plus.n23 plus.t8 651.605
R11 plus.n21 plus.t3 651.605
R12 plus.n6 plus.n3 161.3
R13 plus.n11 plus.n10 161.3
R14 plus.n12 plus.n1 161.3
R15 plus.n13 plus.n0 161.3
R16 plus.n15 plus.n14 161.3
R17 plus.n22 plus.n19 161.3
R18 plus.n27 plus.n26 161.3
R19 plus.n28 plus.n17 161.3
R20 plus.n29 plus.n16 161.3
R21 plus.n31 plus.n30 161.3
R22 plus.n8 plus.n7 80.6037
R23 plus.n9 plus.n2 80.6037
R24 plus.n24 plus.n23 80.6037
R25 plus.n25 plus.n18 80.6037
R26 plus.n7 plus.n2 48.2005
R27 plus.n23 plus.n18 48.2005
R28 plus.n4 plus.n3 44.853
R29 plus.n20 plus.n19 44.853
R30 plus.n11 plus.n2 41.6278
R31 plus.n7 plus.n6 41.6278
R32 plus.n27 plus.n18 41.6278
R33 plus.n23 plus.n22 41.6278
R34 plus plus.n31 34.9384
R35 plus.n14 plus.n13 25.5611
R36 plus.n30 plus.n29 25.5611
R37 plus.n13 plus.n12 22.6399
R38 plus.n29 plus.n28 22.6399
R39 plus.n5 plus.n4 20.5405
R40 plus.n21 plus.n20 20.5405
R41 plus plus.n15 15.3755
R42 plus.n12 plus.n11 6.57323
R43 plus.n6 plus.n5 6.57323
R44 plus.n28 plus.n27 6.57323
R45 plus.n22 plus.n21 6.57323
R46 plus.n9 plus.n8 0.380177
R47 plus.n25 plus.n24 0.380177
R48 plus.n8 plus.n3 0.285035
R49 plus.n10 plus.n9 0.285035
R50 plus.n26 plus.n25 0.285035
R51 plus.n24 plus.n19 0.285035
R52 plus.n10 plus.n1 0.189894
R53 plus.n1 plus.n0 0.189894
R54 plus.n15 plus.n0 0.189894
R55 plus.n31 plus.n16 0.189894
R56 plus.n17 plus.n16 0.189894
R57 plus.n26 plus.n17 0.189894
R58 source.n0 source.t12 44.1297
R59 source.n5 source.t10 44.1296
R60 source.n6 source.t23 44.1296
R61 source.n11 source.t1 44.1296
R62 source.n23 source.t9 44.1295
R63 source.n18 source.t2 44.1295
R64 source.n17 source.t17 44.1295
R65 source.n12 source.t21 44.1295
R66 source.n2 source.n1 43.1397
R67 source.n4 source.n3 43.1397
R68 source.n8 source.n7 43.1397
R69 source.n10 source.n9 43.1397
R70 source.n22 source.n21 43.1396
R71 source.n20 source.n19 43.1396
R72 source.n16 source.n15 43.1396
R73 source.n14 source.n13 43.1396
R74 source.n12 source.n11 28.3225
R75 source.n24 source.n0 22.5725
R76 source.n24 source.n23 5.7505
R77 source.n21 source.t22 0.9905
R78 source.n21 source.t7 0.9905
R79 source.n19 source.t3 0.9905
R80 source.n19 source.t5 0.9905
R81 source.n15 source.t19 0.9905
R82 source.n15 source.t16 0.9905
R83 source.n13 source.t20 0.9905
R84 source.n13 source.t13 0.9905
R85 source.n1 source.t15 0.9905
R86 source.n1 source.t18 0.9905
R87 source.n3 source.t14 0.9905
R88 source.n3 source.t11 0.9905
R89 source.n7 source.t8 0.9905
R90 source.n7 source.t0 0.9905
R91 source.n9 source.t6 0.9905
R92 source.n9 source.t4 0.9905
R93 source.n11 source.n10 0.974638
R94 source.n10 source.n8 0.974638
R95 source.n8 source.n6 0.974638
R96 source.n5 source.n4 0.974638
R97 source.n4 source.n2 0.974638
R98 source.n2 source.n0 0.974638
R99 source.n14 source.n12 0.974638
R100 source.n16 source.n14 0.974638
R101 source.n17 source.n16 0.974638
R102 source.n20 source.n18 0.974638
R103 source.n22 source.n20 0.974638
R104 source.n23 source.n22 0.974638
R105 source.n6 source.n5 0.470328
R106 source.n18 source.n17 0.470328
R107 source source.n24 0.188
R108 drain_left.n6 drain_left.n4 60.7926
R109 drain_left.n3 drain_left.n2 60.7372
R110 drain_left.n3 drain_left.n0 60.7372
R111 drain_left.n8 drain_left.n7 59.8185
R112 drain_left.n6 drain_left.n5 59.8185
R113 drain_left.n3 drain_left.n1 59.8184
R114 drain_left drain_left.n3 38.2984
R115 drain_left drain_left.n8 6.62735
R116 drain_left.n1 drain_left.t9 0.9905
R117 drain_left.n1 drain_left.t3 0.9905
R118 drain_left.n2 drain_left.t8 0.9905
R119 drain_left.n2 drain_left.t11 0.9905
R120 drain_left.n0 drain_left.t10 0.9905
R121 drain_left.n0 drain_left.t4 0.9905
R122 drain_left.n7 drain_left.t2 0.9905
R123 drain_left.n7 drain_left.t7 0.9905
R124 drain_left.n5 drain_left.t5 0.9905
R125 drain_left.n5 drain_left.t6 0.9905
R126 drain_left.n4 drain_left.t0 0.9905
R127 drain_left.n4 drain_left.t1 0.9905
R128 drain_left.n8 drain_left.n6 0.974638
R129 minus.n4 minus.t6 673
R130 minus.n20 minus.t1 673
R131 minus.n3 minus.t5 651.605
R132 minus.n7 minus.t4 651.605
R133 minus.n8 minus.t9 651.605
R134 minus.n12 minus.t10 651.605
R135 minus.n14 minus.t8 651.605
R136 minus.n19 minus.t7 651.605
R137 minus.n23 minus.t11 651.605
R138 minus.n24 minus.t3 651.605
R139 minus.n28 minus.t0 651.605
R140 minus.n30 minus.t2 651.605
R141 minus.n15 minus.n14 161.3
R142 minus.n13 minus.n0 161.3
R143 minus.n12 minus.n11 161.3
R144 minus.n10 minus.n1 161.3
R145 minus.n6 minus.n5 161.3
R146 minus.n31 minus.n30 161.3
R147 minus.n29 minus.n16 161.3
R148 minus.n28 minus.n27 161.3
R149 minus.n26 minus.n17 161.3
R150 minus.n22 minus.n21 161.3
R151 minus.n9 minus.n8 80.6037
R152 minus.n7 minus.n2 80.6037
R153 minus.n25 minus.n24 80.6037
R154 minus.n23 minus.n18 80.6037
R155 minus.n8 minus.n7 48.2005
R156 minus.n24 minus.n23 48.2005
R157 minus.n5 minus.n4 44.853
R158 minus.n21 minus.n20 44.853
R159 minus.n32 minus.n15 44.0876
R160 minus.n7 minus.n6 41.6278
R161 minus.n8 minus.n1 41.6278
R162 minus.n23 minus.n22 41.6278
R163 minus.n24 minus.n17 41.6278
R164 minus.n14 minus.n13 25.5611
R165 minus.n30 minus.n29 25.5611
R166 minus.n13 minus.n12 22.6399
R167 minus.n29 minus.n28 22.6399
R168 minus.n4 minus.n3 20.5405
R169 minus.n20 minus.n19 20.5405
R170 minus.n32 minus.n31 6.70126
R171 minus.n6 minus.n3 6.57323
R172 minus.n12 minus.n1 6.57323
R173 minus.n22 minus.n19 6.57323
R174 minus.n28 minus.n17 6.57323
R175 minus.n9 minus.n2 0.380177
R176 minus.n25 minus.n18 0.380177
R177 minus.n10 minus.n9 0.285035
R178 minus.n5 minus.n2 0.285035
R179 minus.n21 minus.n18 0.285035
R180 minus.n26 minus.n25 0.285035
R181 minus.n15 minus.n0 0.189894
R182 minus.n11 minus.n0 0.189894
R183 minus.n11 minus.n10 0.189894
R184 minus.n27 minus.n26 0.189894
R185 minus.n27 minus.n16 0.189894
R186 minus.n31 minus.n16 0.189894
R187 minus minus.n32 0.188
R188 drain_right.n6 drain_right.n4 60.7926
R189 drain_right.n3 drain_right.n2 60.7372
R190 drain_right.n3 drain_right.n0 60.7372
R191 drain_right.n6 drain_right.n5 59.8185
R192 drain_right.n8 drain_right.n7 59.8185
R193 drain_right.n3 drain_right.n1 59.8184
R194 drain_right drain_right.n3 37.7451
R195 drain_right drain_right.n8 6.62735
R196 drain_right.n1 drain_right.t0 0.9905
R197 drain_right.n1 drain_right.t8 0.9905
R198 drain_right.n2 drain_right.t11 0.9905
R199 drain_right.n2 drain_right.t9 0.9905
R200 drain_right.n0 drain_right.t10 0.9905
R201 drain_right.n0 drain_right.t4 0.9905
R202 drain_right.n4 drain_right.t6 0.9905
R203 drain_right.n4 drain_right.t5 0.9905
R204 drain_right.n5 drain_right.t2 0.9905
R205 drain_right.n5 drain_right.t7 0.9905
R206 drain_right.n7 drain_right.t3 0.9905
R207 drain_right.n7 drain_right.t1 0.9905
R208 drain_right.n8 drain_right.n6 0.974638
C0 source plus 13.406599f
C1 minus drain_right 13.7571f
C2 drain_left drain_right 1.16185f
C3 minus source 13.3926f
C4 minus plus 7.48702f
C5 source drain_left 22.3051f
C6 drain_left plus 13.9834f
C7 source drain_right 22.3077f
C8 drain_right plus 0.381869f
C9 minus drain_left 0.17224f
C10 drain_right a_n2298_n4888# 7.766969f
C11 drain_left a_n2298_n4888# 8.089781f
C12 source a_n2298_n4888# 13.748971f
C13 minus a_n2298_n4888# 9.615657f
C14 plus a_n2298_n4888# 11.64863f
C15 drain_right.t10 a_n2298_n4888# 0.42049f
C16 drain_right.t4 a_n2298_n4888# 0.42049f
C17 drain_right.n0 a_n2298_n4888# 3.85024f
C18 drain_right.t0 a_n2298_n4888# 0.42049f
C19 drain_right.t8 a_n2298_n4888# 0.42049f
C20 drain_right.n1 a_n2298_n4888# 3.84422f
C21 drain_right.t11 a_n2298_n4888# 0.42049f
C22 drain_right.t9 a_n2298_n4888# 0.42049f
C23 drain_right.n2 a_n2298_n4888# 3.85024f
C24 drain_right.n3 a_n2298_n4888# 3.02011f
C25 drain_right.t6 a_n2298_n4888# 0.42049f
C26 drain_right.t5 a_n2298_n4888# 0.42049f
C27 drain_right.n4 a_n2298_n4888# 3.85066f
C28 drain_right.t2 a_n2298_n4888# 0.42049f
C29 drain_right.t7 a_n2298_n4888# 0.42049f
C30 drain_right.n5 a_n2298_n4888# 3.84421f
C31 drain_right.n6 a_n2298_n4888# 0.787355f
C32 drain_right.t3 a_n2298_n4888# 0.42049f
C33 drain_right.t1 a_n2298_n4888# 0.42049f
C34 drain_right.n7 a_n2298_n4888# 3.84421f
C35 drain_right.n8 a_n2298_n4888# 0.630113f
C36 minus.n0 a_n2298_n4888# 0.039315f
C37 minus.n1 a_n2298_n4888# 0.008921f
C38 minus.t10 a_n2298_n4888# 1.78136f
C39 minus.n2 a_n2298_n4888# 0.065483f
C40 minus.t5 a_n2298_n4888# 1.78136f
C41 minus.n3 a_n2298_n4888# 0.663732f
C42 minus.t6 a_n2298_n4888# 1.80243f
C43 minus.n4 a_n2298_n4888# 0.645676f
C44 minus.n5 a_n2298_n4888# 0.180484f
C45 minus.n6 a_n2298_n4888# 0.008921f
C46 minus.t4 a_n2298_n4888# 1.78136f
C47 minus.n7 a_n2298_n4888# 0.67165f
C48 minus.t9 a_n2298_n4888# 1.78136f
C49 minus.n8 a_n2298_n4888# 0.67165f
C50 minus.n9 a_n2298_n4888# 0.065483f
C51 minus.n10 a_n2298_n4888# 0.05246f
C52 minus.n11 a_n2298_n4888# 0.039315f
C53 minus.n12 a_n2298_n4888# 0.660669f
C54 minus.n13 a_n2298_n4888# 0.008921f
C55 minus.t8 a_n2298_n4888# 1.78136f
C56 minus.n14 a_n2298_n4888# 0.660063f
C57 minus.n15 a_n2298_n4888# 1.87384f
C58 minus.n16 a_n2298_n4888# 0.039315f
C59 minus.n17 a_n2298_n4888# 0.008921f
C60 minus.n18 a_n2298_n4888# 0.065483f
C61 minus.t7 a_n2298_n4888# 1.78136f
C62 minus.n19 a_n2298_n4888# 0.663732f
C63 minus.t1 a_n2298_n4888# 1.80243f
C64 minus.n20 a_n2298_n4888# 0.645676f
C65 minus.n21 a_n2298_n4888# 0.180484f
C66 minus.n22 a_n2298_n4888# 0.008921f
C67 minus.t11 a_n2298_n4888# 1.78136f
C68 minus.n23 a_n2298_n4888# 0.67165f
C69 minus.t3 a_n2298_n4888# 1.78136f
C70 minus.n24 a_n2298_n4888# 0.67165f
C71 minus.n25 a_n2298_n4888# 0.065483f
C72 minus.n26 a_n2298_n4888# 0.05246f
C73 minus.n27 a_n2298_n4888# 0.039315f
C74 minus.t0 a_n2298_n4888# 1.78136f
C75 minus.n28 a_n2298_n4888# 0.660669f
C76 minus.n29 a_n2298_n4888# 0.008921f
C77 minus.t2 a_n2298_n4888# 1.78136f
C78 minus.n30 a_n2298_n4888# 0.660063f
C79 minus.n31 a_n2298_n4888# 0.275497f
C80 minus.n32 a_n2298_n4888# 2.2209f
C81 drain_left.t10 a_n2298_n4888# 0.421605f
C82 drain_left.t4 a_n2298_n4888# 0.421605f
C83 drain_left.n0 a_n2298_n4888# 3.86044f
C84 drain_left.t9 a_n2298_n4888# 0.421605f
C85 drain_left.t3 a_n2298_n4888# 0.421605f
C86 drain_left.n1 a_n2298_n4888# 3.8544f
C87 drain_left.t8 a_n2298_n4888# 0.421605f
C88 drain_left.t11 a_n2298_n4888# 0.421605f
C89 drain_left.n2 a_n2298_n4888# 3.86044f
C90 drain_left.n3 a_n2298_n4888# 3.08329f
C91 drain_left.t0 a_n2298_n4888# 0.421605f
C92 drain_left.t1 a_n2298_n4888# 0.421605f
C93 drain_left.n4 a_n2298_n4888# 3.86086f
C94 drain_left.t5 a_n2298_n4888# 0.421605f
C95 drain_left.t6 a_n2298_n4888# 0.421605f
C96 drain_left.n5 a_n2298_n4888# 3.8544f
C97 drain_left.n6 a_n2298_n4888# 0.789441f
C98 drain_left.t2 a_n2298_n4888# 0.421605f
C99 drain_left.t7 a_n2298_n4888# 0.421605f
C100 drain_left.n7 a_n2298_n4888# 3.8544f
C101 drain_left.n8 a_n2298_n4888# 0.631782f
C102 source.t12 a_n2298_n4888# 3.76303f
C103 source.n0 a_n2298_n4888# 1.64614f
C104 source.t15 a_n2298_n4888# 0.329271f
C105 source.t18 a_n2298_n4888# 0.329271f
C106 source.n1 a_n2298_n4888# 2.94382f
C107 source.n2 a_n2298_n4888# 0.344725f
C108 source.t14 a_n2298_n4888# 0.329271f
C109 source.t11 a_n2298_n4888# 0.329271f
C110 source.n3 a_n2298_n4888# 2.94382f
C111 source.n4 a_n2298_n4888# 0.344725f
C112 source.t10 a_n2298_n4888# 3.76304f
C113 source.n5 a_n2298_n4888# 0.389663f
C114 source.t23 a_n2298_n4888# 3.76304f
C115 source.n6 a_n2298_n4888# 0.389663f
C116 source.t8 a_n2298_n4888# 0.329271f
C117 source.t0 a_n2298_n4888# 0.329271f
C118 source.n7 a_n2298_n4888# 2.94382f
C119 source.n8 a_n2298_n4888# 0.344725f
C120 source.t6 a_n2298_n4888# 0.329271f
C121 source.t4 a_n2298_n4888# 0.329271f
C122 source.n9 a_n2298_n4888# 2.94382f
C123 source.n10 a_n2298_n4888# 0.344725f
C124 source.t1 a_n2298_n4888# 3.76304f
C125 source.n11 a_n2298_n4888# 2.02761f
C126 source.t21 a_n2298_n4888# 3.76302f
C127 source.n12 a_n2298_n4888# 2.02764f
C128 source.t20 a_n2298_n4888# 0.329271f
C129 source.t13 a_n2298_n4888# 0.329271f
C130 source.n13 a_n2298_n4888# 2.94383f
C131 source.n14 a_n2298_n4888# 0.344719f
C132 source.t19 a_n2298_n4888# 0.329271f
C133 source.t16 a_n2298_n4888# 0.329271f
C134 source.n15 a_n2298_n4888# 2.94383f
C135 source.n16 a_n2298_n4888# 0.344719f
C136 source.t17 a_n2298_n4888# 3.76302f
C137 source.n17 a_n2298_n4888# 0.389684f
C138 source.t2 a_n2298_n4888# 3.76302f
C139 source.n18 a_n2298_n4888# 0.389684f
C140 source.t3 a_n2298_n4888# 0.329271f
C141 source.t5 a_n2298_n4888# 0.329271f
C142 source.n19 a_n2298_n4888# 2.94383f
C143 source.n20 a_n2298_n4888# 0.344719f
C144 source.t22 a_n2298_n4888# 0.329271f
C145 source.t7 a_n2298_n4888# 0.329271f
C146 source.n21 a_n2298_n4888# 2.94383f
C147 source.n22 a_n2298_n4888# 0.344719f
C148 source.t9 a_n2298_n4888# 3.76302f
C149 source.n23 a_n2298_n4888# 0.530094f
C150 source.n24 a_n2298_n4888# 1.89384f
C151 plus.n0 a_n2298_n4888# 0.039632f
C152 plus.t4 a_n2298_n4888# 1.79574f
C153 plus.t9 a_n2298_n4888# 1.79574f
C154 plus.n1 a_n2298_n4888# 0.039632f
C155 plus.t5 a_n2298_n4888# 1.79574f
C156 plus.n2 a_n2298_n4888# 0.677073f
C157 plus.n3 a_n2298_n4888# 0.181941f
C158 plus.t6 a_n2298_n4888# 1.79574f
C159 plus.t10 a_n2298_n4888# 1.79574f
C160 plus.t11 a_n2298_n4888# 1.81698f
C161 plus.n4 a_n2298_n4888# 0.650888f
C162 plus.n5 a_n2298_n4888# 0.66909f
C163 plus.n6 a_n2298_n4888# 0.008993f
C164 plus.n7 a_n2298_n4888# 0.677073f
C165 plus.n8 a_n2298_n4888# 0.066012f
C166 plus.n9 a_n2298_n4888# 0.066012f
C167 plus.n10 a_n2298_n4888# 0.052884f
C168 plus.n11 a_n2298_n4888# 0.008993f
C169 plus.n12 a_n2298_n4888# 0.666003f
C170 plus.n13 a_n2298_n4888# 0.008993f
C171 plus.n14 a_n2298_n4888# 0.665392f
C172 plus.n15 a_n2298_n4888# 0.620063f
C173 plus.n16 a_n2298_n4888# 0.039632f
C174 plus.t1 a_n2298_n4888# 1.79574f
C175 plus.n17 a_n2298_n4888# 0.039632f
C176 plus.t7 a_n2298_n4888# 1.79574f
C177 plus.t2 a_n2298_n4888# 1.79574f
C178 plus.n18 a_n2298_n4888# 0.677073f
C179 plus.n19 a_n2298_n4888# 0.181941f
C180 plus.t8 a_n2298_n4888# 1.79574f
C181 plus.t0 a_n2298_n4888# 1.81698f
C182 plus.n20 a_n2298_n4888# 0.650888f
C183 plus.t3 a_n2298_n4888# 1.79574f
C184 plus.n21 a_n2298_n4888# 0.66909f
C185 plus.n22 a_n2298_n4888# 0.008993f
C186 plus.n23 a_n2298_n4888# 0.677073f
C187 plus.n24 a_n2298_n4888# 0.066012f
C188 plus.n25 a_n2298_n4888# 0.066012f
C189 plus.n26 a_n2298_n4888# 0.052884f
C190 plus.n27 a_n2298_n4888# 0.008993f
C191 plus.n28 a_n2298_n4888# 0.666003f
C192 plus.n29 a_n2298_n4888# 0.008993f
C193 plus.n30 a_n2298_n4888# 0.665392f
C194 plus.n31 a_n2298_n4888# 1.50761f
.ends

