* NGSPICE file created from diffpair621.ext - technology: sky130A

.subckt diffpair621 minus drain_right drain_left source plus
X0 drain_left plus source a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X1 source plus drain_left a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X2 a_n1334_n4888# a_n1334_n4888# a_n1334_n4888# a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.7
X3 source minus drain_right a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X4 source plus drain_left a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X5 drain_right minus source a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X6 source minus drain_right a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X7 a_n1334_n4888# a_n1334_n4888# a_n1334_n4888# a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X8 drain_right minus source a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X9 drain_left plus source a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X10 a_n1334_n4888# a_n1334_n4888# a_n1334_n4888# a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X11 a_n1334_n4888# a_n1334_n4888# a_n1334_n4888# a_n1334_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
.ends

