* NGSPICE file created from diffpair424.ext - technology: sky130A

.subckt diffpair424 minus drain_right drain_left source plus
X0 source.t18 plus.t0 drain_left.t8 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X1 source.t17 plus.t1 drain_left.t9 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X2 a_n1412_n3288# a_n1412_n3288# a_n1412_n3288# a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.25
X3 source.t4 minus.t0 drain_right.t9 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X4 source.t0 minus.t1 drain_right.t8 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X5 source.t3 minus.t2 drain_right.t7 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X6 drain_left.t5 plus.t2 source.t16 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X7 drain_left.t6 plus.t3 source.t15 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X8 drain_right.t6 minus.t3 source.t2 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X9 drain_left.t1 plus.t4 source.t14 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X10 drain_left.t2 plus.t5 source.t13 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X11 drain_left.t0 plus.t6 source.t12 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X12 a_n1412_n3288# a_n1412_n3288# a_n1412_n3288# a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X13 drain_right.t5 minus.t4 source.t8 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X14 drain_right.t4 minus.t5 source.t1 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X15 source.t5 minus.t6 drain_right.t3 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X16 source.t11 plus.t7 drain_left.t7 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X17 a_n1412_n3288# a_n1412_n3288# a_n1412_n3288# a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X18 drain_right.t2 minus.t7 source.t7 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X19 drain_right.t1 minus.t8 source.t6 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X20 drain_left.t4 plus.t8 source.t10 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X21 a_n1412_n3288# a_n1412_n3288# a_n1412_n3288# a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X22 drain_right.t0 minus.t9 source.t19 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X23 source.t9 plus.t9 drain_left.t3 a_n1412_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
R0 plus.n2 plus.t3 1342
R1 plus.n8 plus.t5 1342
R2 plus.n12 plus.t8 1342
R3 plus.n18 plus.t2 1342
R4 plus.n1 plus.t1 1282.12
R5 plus.n5 plus.t6 1282.12
R6 plus.n7 plus.t0 1282.12
R7 plus.n11 plus.t7 1282.12
R8 plus.n15 plus.t4 1282.12
R9 plus.n17 plus.t9 1282.12
R10 plus.n3 plus.n2 161.489
R11 plus.n13 plus.n12 161.489
R12 plus.n4 plus.n3 161.3
R13 plus.n6 plus.n0 161.3
R14 plus.n9 plus.n8 161.3
R15 plus.n14 plus.n13 161.3
R16 plus.n16 plus.n10 161.3
R17 plus.n19 plus.n18 161.3
R18 plus.n4 plus.n1 48.2005
R19 plus.n7 plus.n6 48.2005
R20 plus.n17 plus.n16 48.2005
R21 plus.n14 plus.n11 48.2005
R22 plus.n5 plus.n4 36.5157
R23 plus.n6 plus.n5 36.5157
R24 plus.n16 plus.n15 36.5157
R25 plus.n15 plus.n14 36.5157
R26 plus plus.n19 28.3664
R27 plus.n2 plus.n1 24.8308
R28 plus.n8 plus.n7 24.8308
R29 plus.n18 plus.n17 24.8308
R30 plus.n12 plus.n11 24.8308
R31 plus plus.n9 12.1596
R32 plus.n3 plus.n0 0.189894
R33 plus.n9 plus.n0 0.189894
R34 plus.n19 plus.n10 0.189894
R35 plus.n13 plus.n10 0.189894
R36 drain_left.n60 drain_left.n0 289.615
R37 drain_left.n129 drain_left.n69 289.615
R38 drain_left.n20 drain_left.n19 185
R39 drain_left.n25 drain_left.n24 185
R40 drain_left.n27 drain_left.n26 185
R41 drain_left.n16 drain_left.n15 185
R42 drain_left.n33 drain_left.n32 185
R43 drain_left.n35 drain_left.n34 185
R44 drain_left.n12 drain_left.n11 185
R45 drain_left.n42 drain_left.n41 185
R46 drain_left.n43 drain_left.n10 185
R47 drain_left.n45 drain_left.n44 185
R48 drain_left.n8 drain_left.n7 185
R49 drain_left.n51 drain_left.n50 185
R50 drain_left.n53 drain_left.n52 185
R51 drain_left.n4 drain_left.n3 185
R52 drain_left.n59 drain_left.n58 185
R53 drain_left.n61 drain_left.n60 185
R54 drain_left.n130 drain_left.n129 185
R55 drain_left.n128 drain_left.n127 185
R56 drain_left.n73 drain_left.n72 185
R57 drain_left.n122 drain_left.n121 185
R58 drain_left.n120 drain_left.n119 185
R59 drain_left.n77 drain_left.n76 185
R60 drain_left.n114 drain_left.n113 185
R61 drain_left.n112 drain_left.n79 185
R62 drain_left.n111 drain_left.n110 185
R63 drain_left.n82 drain_left.n80 185
R64 drain_left.n105 drain_left.n104 185
R65 drain_left.n103 drain_left.n102 185
R66 drain_left.n86 drain_left.n85 185
R67 drain_left.n97 drain_left.n96 185
R68 drain_left.n95 drain_left.n94 185
R69 drain_left.n90 drain_left.n89 185
R70 drain_left.n21 drain_left.t5 149.524
R71 drain_left.n91 drain_left.t6 149.524
R72 drain_left.n25 drain_left.n19 104.615
R73 drain_left.n26 drain_left.n25 104.615
R74 drain_left.n26 drain_left.n15 104.615
R75 drain_left.n33 drain_left.n15 104.615
R76 drain_left.n34 drain_left.n33 104.615
R77 drain_left.n34 drain_left.n11 104.615
R78 drain_left.n42 drain_left.n11 104.615
R79 drain_left.n43 drain_left.n42 104.615
R80 drain_left.n44 drain_left.n43 104.615
R81 drain_left.n44 drain_left.n7 104.615
R82 drain_left.n51 drain_left.n7 104.615
R83 drain_left.n52 drain_left.n51 104.615
R84 drain_left.n52 drain_left.n3 104.615
R85 drain_left.n59 drain_left.n3 104.615
R86 drain_left.n60 drain_left.n59 104.615
R87 drain_left.n129 drain_left.n128 104.615
R88 drain_left.n128 drain_left.n72 104.615
R89 drain_left.n121 drain_left.n72 104.615
R90 drain_left.n121 drain_left.n120 104.615
R91 drain_left.n120 drain_left.n76 104.615
R92 drain_left.n113 drain_left.n76 104.615
R93 drain_left.n113 drain_left.n112 104.615
R94 drain_left.n112 drain_left.n111 104.615
R95 drain_left.n111 drain_left.n80 104.615
R96 drain_left.n104 drain_left.n80 104.615
R97 drain_left.n104 drain_left.n103 104.615
R98 drain_left.n103 drain_left.n85 104.615
R99 drain_left.n96 drain_left.n85 104.615
R100 drain_left.n96 drain_left.n95 104.615
R101 drain_left.n95 drain_left.n89 104.615
R102 drain_left.n68 drain_left.n67 59.8722
R103 drain_left.n135 drain_left.n134 59.5527
R104 drain_left.n66 drain_left.n65 59.5525
R105 drain_left.n137 drain_left.n136 59.5525
R106 drain_left.t5 drain_left.n19 52.3082
R107 drain_left.t6 drain_left.n89 52.3082
R108 drain_left.n66 drain_left.n64 47.0369
R109 drain_left.n135 drain_left.n133 47.0369
R110 drain_left drain_left.n68 29.4921
R111 drain_left.n45 drain_left.n10 13.1884
R112 drain_left.n114 drain_left.n79 13.1884
R113 drain_left.n41 drain_left.n40 12.8005
R114 drain_left.n46 drain_left.n8 12.8005
R115 drain_left.n115 drain_left.n77 12.8005
R116 drain_left.n110 drain_left.n81 12.8005
R117 drain_left.n39 drain_left.n12 12.0247
R118 drain_left.n50 drain_left.n49 12.0247
R119 drain_left.n119 drain_left.n118 12.0247
R120 drain_left.n109 drain_left.n82 12.0247
R121 drain_left.n36 drain_left.n35 11.249
R122 drain_left.n53 drain_left.n6 11.249
R123 drain_left.n122 drain_left.n75 11.249
R124 drain_left.n106 drain_left.n105 11.249
R125 drain_left.n32 drain_left.n14 10.4732
R126 drain_left.n54 drain_left.n4 10.4732
R127 drain_left.n123 drain_left.n73 10.4732
R128 drain_left.n102 drain_left.n84 10.4732
R129 drain_left.n21 drain_left.n20 10.2747
R130 drain_left.n91 drain_left.n90 10.2747
R131 drain_left.n31 drain_left.n16 9.69747
R132 drain_left.n58 drain_left.n57 9.69747
R133 drain_left.n127 drain_left.n126 9.69747
R134 drain_left.n101 drain_left.n86 9.69747
R135 drain_left.n64 drain_left.n63 9.45567
R136 drain_left.n133 drain_left.n132 9.45567
R137 drain_left.n63 drain_left.n62 9.3005
R138 drain_left.n2 drain_left.n1 9.3005
R139 drain_left.n57 drain_left.n56 9.3005
R140 drain_left.n55 drain_left.n54 9.3005
R141 drain_left.n6 drain_left.n5 9.3005
R142 drain_left.n49 drain_left.n48 9.3005
R143 drain_left.n47 drain_left.n46 9.3005
R144 drain_left.n23 drain_left.n22 9.3005
R145 drain_left.n18 drain_left.n17 9.3005
R146 drain_left.n29 drain_left.n28 9.3005
R147 drain_left.n31 drain_left.n30 9.3005
R148 drain_left.n14 drain_left.n13 9.3005
R149 drain_left.n37 drain_left.n36 9.3005
R150 drain_left.n39 drain_left.n38 9.3005
R151 drain_left.n40 drain_left.n9 9.3005
R152 drain_left.n93 drain_left.n92 9.3005
R153 drain_left.n88 drain_left.n87 9.3005
R154 drain_left.n99 drain_left.n98 9.3005
R155 drain_left.n101 drain_left.n100 9.3005
R156 drain_left.n84 drain_left.n83 9.3005
R157 drain_left.n107 drain_left.n106 9.3005
R158 drain_left.n109 drain_left.n108 9.3005
R159 drain_left.n81 drain_left.n78 9.3005
R160 drain_left.n132 drain_left.n131 9.3005
R161 drain_left.n71 drain_left.n70 9.3005
R162 drain_left.n126 drain_left.n125 9.3005
R163 drain_left.n124 drain_left.n123 9.3005
R164 drain_left.n75 drain_left.n74 9.3005
R165 drain_left.n118 drain_left.n117 9.3005
R166 drain_left.n116 drain_left.n115 9.3005
R167 drain_left.n28 drain_left.n27 8.92171
R168 drain_left.n61 drain_left.n2 8.92171
R169 drain_left.n130 drain_left.n71 8.92171
R170 drain_left.n98 drain_left.n97 8.92171
R171 drain_left.n24 drain_left.n18 8.14595
R172 drain_left.n62 drain_left.n0 8.14595
R173 drain_left.n131 drain_left.n69 8.14595
R174 drain_left.n94 drain_left.n88 8.14595
R175 drain_left.n23 drain_left.n20 7.3702
R176 drain_left.n93 drain_left.n90 7.3702
R177 drain_left drain_left.n137 6.15322
R178 drain_left.n24 drain_left.n23 5.81868
R179 drain_left.n64 drain_left.n0 5.81868
R180 drain_left.n133 drain_left.n69 5.81868
R181 drain_left.n94 drain_left.n93 5.81868
R182 drain_left.n27 drain_left.n18 5.04292
R183 drain_left.n62 drain_left.n61 5.04292
R184 drain_left.n131 drain_left.n130 5.04292
R185 drain_left.n97 drain_left.n88 5.04292
R186 drain_left.n28 drain_left.n16 4.26717
R187 drain_left.n58 drain_left.n2 4.26717
R188 drain_left.n127 drain_left.n71 4.26717
R189 drain_left.n98 drain_left.n86 4.26717
R190 drain_left.n32 drain_left.n31 3.49141
R191 drain_left.n57 drain_left.n4 3.49141
R192 drain_left.n126 drain_left.n73 3.49141
R193 drain_left.n102 drain_left.n101 3.49141
R194 drain_left.n22 drain_left.n21 2.84303
R195 drain_left.n92 drain_left.n91 2.84303
R196 drain_left.n35 drain_left.n14 2.71565
R197 drain_left.n54 drain_left.n53 2.71565
R198 drain_left.n123 drain_left.n122 2.71565
R199 drain_left.n105 drain_left.n84 2.71565
R200 drain_left.n36 drain_left.n12 1.93989
R201 drain_left.n50 drain_left.n6 1.93989
R202 drain_left.n119 drain_left.n75 1.93989
R203 drain_left.n106 drain_left.n82 1.93989
R204 drain_left.n67 drain_left.t7 1.6505
R205 drain_left.n67 drain_left.t4 1.6505
R206 drain_left.n65 drain_left.t3 1.6505
R207 drain_left.n65 drain_left.t1 1.6505
R208 drain_left.n136 drain_left.t8 1.6505
R209 drain_left.n136 drain_left.t2 1.6505
R210 drain_left.n134 drain_left.t9 1.6505
R211 drain_left.n134 drain_left.t0 1.6505
R212 drain_left.n41 drain_left.n39 1.16414
R213 drain_left.n49 drain_left.n8 1.16414
R214 drain_left.n118 drain_left.n77 1.16414
R215 drain_left.n110 drain_left.n109 1.16414
R216 drain_left.n137 drain_left.n135 0.5005
R217 drain_left.n40 drain_left.n10 0.388379
R218 drain_left.n46 drain_left.n45 0.388379
R219 drain_left.n115 drain_left.n114 0.388379
R220 drain_left.n81 drain_left.n79 0.388379
R221 drain_left.n22 drain_left.n17 0.155672
R222 drain_left.n29 drain_left.n17 0.155672
R223 drain_left.n30 drain_left.n29 0.155672
R224 drain_left.n30 drain_left.n13 0.155672
R225 drain_left.n37 drain_left.n13 0.155672
R226 drain_left.n38 drain_left.n37 0.155672
R227 drain_left.n38 drain_left.n9 0.155672
R228 drain_left.n47 drain_left.n9 0.155672
R229 drain_left.n48 drain_left.n47 0.155672
R230 drain_left.n48 drain_left.n5 0.155672
R231 drain_left.n55 drain_left.n5 0.155672
R232 drain_left.n56 drain_left.n55 0.155672
R233 drain_left.n56 drain_left.n1 0.155672
R234 drain_left.n63 drain_left.n1 0.155672
R235 drain_left.n132 drain_left.n70 0.155672
R236 drain_left.n125 drain_left.n70 0.155672
R237 drain_left.n125 drain_left.n124 0.155672
R238 drain_left.n124 drain_left.n74 0.155672
R239 drain_left.n117 drain_left.n74 0.155672
R240 drain_left.n117 drain_left.n116 0.155672
R241 drain_left.n116 drain_left.n78 0.155672
R242 drain_left.n108 drain_left.n78 0.155672
R243 drain_left.n108 drain_left.n107 0.155672
R244 drain_left.n107 drain_left.n83 0.155672
R245 drain_left.n100 drain_left.n83 0.155672
R246 drain_left.n100 drain_left.n99 0.155672
R247 drain_left.n99 drain_left.n87 0.155672
R248 drain_left.n92 drain_left.n87 0.155672
R249 drain_left.n68 drain_left.n66 0.070154
R250 source.n274 source.n214 289.615
R251 source.n204 source.n144 289.615
R252 source.n60 source.n0 289.615
R253 source.n130 source.n70 289.615
R254 source.n234 source.n233 185
R255 source.n239 source.n238 185
R256 source.n241 source.n240 185
R257 source.n230 source.n229 185
R258 source.n247 source.n246 185
R259 source.n249 source.n248 185
R260 source.n226 source.n225 185
R261 source.n256 source.n255 185
R262 source.n257 source.n224 185
R263 source.n259 source.n258 185
R264 source.n222 source.n221 185
R265 source.n265 source.n264 185
R266 source.n267 source.n266 185
R267 source.n218 source.n217 185
R268 source.n273 source.n272 185
R269 source.n275 source.n274 185
R270 source.n164 source.n163 185
R271 source.n169 source.n168 185
R272 source.n171 source.n170 185
R273 source.n160 source.n159 185
R274 source.n177 source.n176 185
R275 source.n179 source.n178 185
R276 source.n156 source.n155 185
R277 source.n186 source.n185 185
R278 source.n187 source.n154 185
R279 source.n189 source.n188 185
R280 source.n152 source.n151 185
R281 source.n195 source.n194 185
R282 source.n197 source.n196 185
R283 source.n148 source.n147 185
R284 source.n203 source.n202 185
R285 source.n205 source.n204 185
R286 source.n61 source.n60 185
R287 source.n59 source.n58 185
R288 source.n4 source.n3 185
R289 source.n53 source.n52 185
R290 source.n51 source.n50 185
R291 source.n8 source.n7 185
R292 source.n45 source.n44 185
R293 source.n43 source.n10 185
R294 source.n42 source.n41 185
R295 source.n13 source.n11 185
R296 source.n36 source.n35 185
R297 source.n34 source.n33 185
R298 source.n17 source.n16 185
R299 source.n28 source.n27 185
R300 source.n26 source.n25 185
R301 source.n21 source.n20 185
R302 source.n131 source.n130 185
R303 source.n129 source.n128 185
R304 source.n74 source.n73 185
R305 source.n123 source.n122 185
R306 source.n121 source.n120 185
R307 source.n78 source.n77 185
R308 source.n115 source.n114 185
R309 source.n113 source.n80 185
R310 source.n112 source.n111 185
R311 source.n83 source.n81 185
R312 source.n106 source.n105 185
R313 source.n104 source.n103 185
R314 source.n87 source.n86 185
R315 source.n98 source.n97 185
R316 source.n96 source.n95 185
R317 source.n91 source.n90 185
R318 source.n235 source.t2 149.524
R319 source.n165 source.t10 149.524
R320 source.n22 source.t13 149.524
R321 source.n92 source.t1 149.524
R322 source.n239 source.n233 104.615
R323 source.n240 source.n239 104.615
R324 source.n240 source.n229 104.615
R325 source.n247 source.n229 104.615
R326 source.n248 source.n247 104.615
R327 source.n248 source.n225 104.615
R328 source.n256 source.n225 104.615
R329 source.n257 source.n256 104.615
R330 source.n258 source.n257 104.615
R331 source.n258 source.n221 104.615
R332 source.n265 source.n221 104.615
R333 source.n266 source.n265 104.615
R334 source.n266 source.n217 104.615
R335 source.n273 source.n217 104.615
R336 source.n274 source.n273 104.615
R337 source.n169 source.n163 104.615
R338 source.n170 source.n169 104.615
R339 source.n170 source.n159 104.615
R340 source.n177 source.n159 104.615
R341 source.n178 source.n177 104.615
R342 source.n178 source.n155 104.615
R343 source.n186 source.n155 104.615
R344 source.n187 source.n186 104.615
R345 source.n188 source.n187 104.615
R346 source.n188 source.n151 104.615
R347 source.n195 source.n151 104.615
R348 source.n196 source.n195 104.615
R349 source.n196 source.n147 104.615
R350 source.n203 source.n147 104.615
R351 source.n204 source.n203 104.615
R352 source.n60 source.n59 104.615
R353 source.n59 source.n3 104.615
R354 source.n52 source.n3 104.615
R355 source.n52 source.n51 104.615
R356 source.n51 source.n7 104.615
R357 source.n44 source.n7 104.615
R358 source.n44 source.n43 104.615
R359 source.n43 source.n42 104.615
R360 source.n42 source.n11 104.615
R361 source.n35 source.n11 104.615
R362 source.n35 source.n34 104.615
R363 source.n34 source.n16 104.615
R364 source.n27 source.n16 104.615
R365 source.n27 source.n26 104.615
R366 source.n26 source.n20 104.615
R367 source.n130 source.n129 104.615
R368 source.n129 source.n73 104.615
R369 source.n122 source.n73 104.615
R370 source.n122 source.n121 104.615
R371 source.n121 source.n77 104.615
R372 source.n114 source.n77 104.615
R373 source.n114 source.n113 104.615
R374 source.n113 source.n112 104.615
R375 source.n112 source.n81 104.615
R376 source.n105 source.n81 104.615
R377 source.n105 source.n104 104.615
R378 source.n104 source.n86 104.615
R379 source.n97 source.n86 104.615
R380 source.n97 source.n96 104.615
R381 source.n96 source.n90 104.615
R382 source.t2 source.n233 52.3082
R383 source.t10 source.n163 52.3082
R384 source.t13 source.n20 52.3082
R385 source.t1 source.n90 52.3082
R386 source.n67 source.n66 42.8739
R387 source.n69 source.n68 42.8739
R388 source.n137 source.n136 42.8739
R389 source.n139 source.n138 42.8739
R390 source.n213 source.n212 42.8737
R391 source.n211 source.n210 42.8737
R392 source.n143 source.n142 42.8737
R393 source.n141 source.n140 42.8737
R394 source.n279 source.n278 29.8581
R395 source.n209 source.n208 29.8581
R396 source.n65 source.n64 29.8581
R397 source.n135 source.n134 29.8581
R398 source.n141 source.n139 22.2877
R399 source.n280 source.n65 16.2748
R400 source.n259 source.n224 13.1884
R401 source.n189 source.n154 13.1884
R402 source.n45 source.n10 13.1884
R403 source.n115 source.n80 13.1884
R404 source.n255 source.n254 12.8005
R405 source.n260 source.n222 12.8005
R406 source.n185 source.n184 12.8005
R407 source.n190 source.n152 12.8005
R408 source.n46 source.n8 12.8005
R409 source.n41 source.n12 12.8005
R410 source.n116 source.n78 12.8005
R411 source.n111 source.n82 12.8005
R412 source.n253 source.n226 12.0247
R413 source.n264 source.n263 12.0247
R414 source.n183 source.n156 12.0247
R415 source.n194 source.n193 12.0247
R416 source.n50 source.n49 12.0247
R417 source.n40 source.n13 12.0247
R418 source.n120 source.n119 12.0247
R419 source.n110 source.n83 12.0247
R420 source.n250 source.n249 11.249
R421 source.n267 source.n220 11.249
R422 source.n180 source.n179 11.249
R423 source.n197 source.n150 11.249
R424 source.n53 source.n6 11.249
R425 source.n37 source.n36 11.249
R426 source.n123 source.n76 11.249
R427 source.n107 source.n106 11.249
R428 source.n246 source.n228 10.4732
R429 source.n268 source.n218 10.4732
R430 source.n176 source.n158 10.4732
R431 source.n198 source.n148 10.4732
R432 source.n54 source.n4 10.4732
R433 source.n33 source.n15 10.4732
R434 source.n124 source.n74 10.4732
R435 source.n103 source.n85 10.4732
R436 source.n235 source.n234 10.2747
R437 source.n165 source.n164 10.2747
R438 source.n22 source.n21 10.2747
R439 source.n92 source.n91 10.2747
R440 source.n245 source.n230 9.69747
R441 source.n272 source.n271 9.69747
R442 source.n175 source.n160 9.69747
R443 source.n202 source.n201 9.69747
R444 source.n58 source.n57 9.69747
R445 source.n32 source.n17 9.69747
R446 source.n128 source.n127 9.69747
R447 source.n102 source.n87 9.69747
R448 source.n278 source.n277 9.45567
R449 source.n208 source.n207 9.45567
R450 source.n64 source.n63 9.45567
R451 source.n134 source.n133 9.45567
R452 source.n277 source.n276 9.3005
R453 source.n216 source.n215 9.3005
R454 source.n271 source.n270 9.3005
R455 source.n269 source.n268 9.3005
R456 source.n220 source.n219 9.3005
R457 source.n263 source.n262 9.3005
R458 source.n261 source.n260 9.3005
R459 source.n237 source.n236 9.3005
R460 source.n232 source.n231 9.3005
R461 source.n243 source.n242 9.3005
R462 source.n245 source.n244 9.3005
R463 source.n228 source.n227 9.3005
R464 source.n251 source.n250 9.3005
R465 source.n253 source.n252 9.3005
R466 source.n254 source.n223 9.3005
R467 source.n207 source.n206 9.3005
R468 source.n146 source.n145 9.3005
R469 source.n201 source.n200 9.3005
R470 source.n199 source.n198 9.3005
R471 source.n150 source.n149 9.3005
R472 source.n193 source.n192 9.3005
R473 source.n191 source.n190 9.3005
R474 source.n167 source.n166 9.3005
R475 source.n162 source.n161 9.3005
R476 source.n173 source.n172 9.3005
R477 source.n175 source.n174 9.3005
R478 source.n158 source.n157 9.3005
R479 source.n181 source.n180 9.3005
R480 source.n183 source.n182 9.3005
R481 source.n184 source.n153 9.3005
R482 source.n24 source.n23 9.3005
R483 source.n19 source.n18 9.3005
R484 source.n30 source.n29 9.3005
R485 source.n32 source.n31 9.3005
R486 source.n15 source.n14 9.3005
R487 source.n38 source.n37 9.3005
R488 source.n40 source.n39 9.3005
R489 source.n12 source.n9 9.3005
R490 source.n63 source.n62 9.3005
R491 source.n2 source.n1 9.3005
R492 source.n57 source.n56 9.3005
R493 source.n55 source.n54 9.3005
R494 source.n6 source.n5 9.3005
R495 source.n49 source.n48 9.3005
R496 source.n47 source.n46 9.3005
R497 source.n94 source.n93 9.3005
R498 source.n89 source.n88 9.3005
R499 source.n100 source.n99 9.3005
R500 source.n102 source.n101 9.3005
R501 source.n85 source.n84 9.3005
R502 source.n108 source.n107 9.3005
R503 source.n110 source.n109 9.3005
R504 source.n82 source.n79 9.3005
R505 source.n133 source.n132 9.3005
R506 source.n72 source.n71 9.3005
R507 source.n127 source.n126 9.3005
R508 source.n125 source.n124 9.3005
R509 source.n76 source.n75 9.3005
R510 source.n119 source.n118 9.3005
R511 source.n117 source.n116 9.3005
R512 source.n242 source.n241 8.92171
R513 source.n275 source.n216 8.92171
R514 source.n172 source.n171 8.92171
R515 source.n205 source.n146 8.92171
R516 source.n61 source.n2 8.92171
R517 source.n29 source.n28 8.92171
R518 source.n131 source.n72 8.92171
R519 source.n99 source.n98 8.92171
R520 source.n238 source.n232 8.14595
R521 source.n276 source.n214 8.14595
R522 source.n168 source.n162 8.14595
R523 source.n206 source.n144 8.14595
R524 source.n62 source.n0 8.14595
R525 source.n25 source.n19 8.14595
R526 source.n132 source.n70 8.14595
R527 source.n95 source.n89 8.14595
R528 source.n237 source.n234 7.3702
R529 source.n167 source.n164 7.3702
R530 source.n24 source.n21 7.3702
R531 source.n94 source.n91 7.3702
R532 source.n238 source.n237 5.81868
R533 source.n278 source.n214 5.81868
R534 source.n168 source.n167 5.81868
R535 source.n208 source.n144 5.81868
R536 source.n64 source.n0 5.81868
R537 source.n25 source.n24 5.81868
R538 source.n134 source.n70 5.81868
R539 source.n95 source.n94 5.81868
R540 source.n280 source.n279 5.51343
R541 source.n241 source.n232 5.04292
R542 source.n276 source.n275 5.04292
R543 source.n171 source.n162 5.04292
R544 source.n206 source.n205 5.04292
R545 source.n62 source.n61 5.04292
R546 source.n28 source.n19 5.04292
R547 source.n132 source.n131 5.04292
R548 source.n98 source.n89 5.04292
R549 source.n242 source.n230 4.26717
R550 source.n272 source.n216 4.26717
R551 source.n172 source.n160 4.26717
R552 source.n202 source.n146 4.26717
R553 source.n58 source.n2 4.26717
R554 source.n29 source.n17 4.26717
R555 source.n128 source.n72 4.26717
R556 source.n99 source.n87 4.26717
R557 source.n246 source.n245 3.49141
R558 source.n271 source.n218 3.49141
R559 source.n176 source.n175 3.49141
R560 source.n201 source.n148 3.49141
R561 source.n57 source.n4 3.49141
R562 source.n33 source.n32 3.49141
R563 source.n127 source.n74 3.49141
R564 source.n103 source.n102 3.49141
R565 source.n236 source.n235 2.84303
R566 source.n166 source.n165 2.84303
R567 source.n23 source.n22 2.84303
R568 source.n93 source.n92 2.84303
R569 source.n249 source.n228 2.71565
R570 source.n268 source.n267 2.71565
R571 source.n179 source.n158 2.71565
R572 source.n198 source.n197 2.71565
R573 source.n54 source.n53 2.71565
R574 source.n36 source.n15 2.71565
R575 source.n124 source.n123 2.71565
R576 source.n106 source.n85 2.71565
R577 source.n250 source.n226 1.93989
R578 source.n264 source.n220 1.93989
R579 source.n180 source.n156 1.93989
R580 source.n194 source.n150 1.93989
R581 source.n50 source.n6 1.93989
R582 source.n37 source.n13 1.93989
R583 source.n120 source.n76 1.93989
R584 source.n107 source.n83 1.93989
R585 source.n212 source.t7 1.6505
R586 source.n212 source.t5 1.6505
R587 source.n210 source.t19 1.6505
R588 source.n210 source.t3 1.6505
R589 source.n142 source.t14 1.6505
R590 source.n142 source.t11 1.6505
R591 source.n140 source.t16 1.6505
R592 source.n140 source.t9 1.6505
R593 source.n66 source.t12 1.6505
R594 source.n66 source.t18 1.6505
R595 source.n68 source.t15 1.6505
R596 source.n68 source.t17 1.6505
R597 source.n136 source.t8 1.6505
R598 source.n136 source.t0 1.6505
R599 source.n138 source.t6 1.6505
R600 source.n138 source.t4 1.6505
R601 source.n255 source.n253 1.16414
R602 source.n263 source.n222 1.16414
R603 source.n185 source.n183 1.16414
R604 source.n193 source.n152 1.16414
R605 source.n49 source.n8 1.16414
R606 source.n41 source.n40 1.16414
R607 source.n119 source.n78 1.16414
R608 source.n111 source.n110 1.16414
R609 source.n135 source.n69 0.720328
R610 source.n211 source.n209 0.720328
R611 source.n139 source.n137 0.5005
R612 source.n137 source.n135 0.5005
R613 source.n69 source.n67 0.5005
R614 source.n67 source.n65 0.5005
R615 source.n143 source.n141 0.5005
R616 source.n209 source.n143 0.5005
R617 source.n213 source.n211 0.5005
R618 source.n279 source.n213 0.5005
R619 source.n254 source.n224 0.388379
R620 source.n260 source.n259 0.388379
R621 source.n184 source.n154 0.388379
R622 source.n190 source.n189 0.388379
R623 source.n46 source.n45 0.388379
R624 source.n12 source.n10 0.388379
R625 source.n116 source.n115 0.388379
R626 source.n82 source.n80 0.388379
R627 source source.n280 0.188
R628 source.n236 source.n231 0.155672
R629 source.n243 source.n231 0.155672
R630 source.n244 source.n243 0.155672
R631 source.n244 source.n227 0.155672
R632 source.n251 source.n227 0.155672
R633 source.n252 source.n251 0.155672
R634 source.n252 source.n223 0.155672
R635 source.n261 source.n223 0.155672
R636 source.n262 source.n261 0.155672
R637 source.n262 source.n219 0.155672
R638 source.n269 source.n219 0.155672
R639 source.n270 source.n269 0.155672
R640 source.n270 source.n215 0.155672
R641 source.n277 source.n215 0.155672
R642 source.n166 source.n161 0.155672
R643 source.n173 source.n161 0.155672
R644 source.n174 source.n173 0.155672
R645 source.n174 source.n157 0.155672
R646 source.n181 source.n157 0.155672
R647 source.n182 source.n181 0.155672
R648 source.n182 source.n153 0.155672
R649 source.n191 source.n153 0.155672
R650 source.n192 source.n191 0.155672
R651 source.n192 source.n149 0.155672
R652 source.n199 source.n149 0.155672
R653 source.n200 source.n199 0.155672
R654 source.n200 source.n145 0.155672
R655 source.n207 source.n145 0.155672
R656 source.n63 source.n1 0.155672
R657 source.n56 source.n1 0.155672
R658 source.n56 source.n55 0.155672
R659 source.n55 source.n5 0.155672
R660 source.n48 source.n5 0.155672
R661 source.n48 source.n47 0.155672
R662 source.n47 source.n9 0.155672
R663 source.n39 source.n9 0.155672
R664 source.n39 source.n38 0.155672
R665 source.n38 source.n14 0.155672
R666 source.n31 source.n14 0.155672
R667 source.n31 source.n30 0.155672
R668 source.n30 source.n18 0.155672
R669 source.n23 source.n18 0.155672
R670 source.n133 source.n71 0.155672
R671 source.n126 source.n71 0.155672
R672 source.n126 source.n125 0.155672
R673 source.n125 source.n75 0.155672
R674 source.n118 source.n75 0.155672
R675 source.n118 source.n117 0.155672
R676 source.n117 source.n79 0.155672
R677 source.n109 source.n79 0.155672
R678 source.n109 source.n108 0.155672
R679 source.n108 source.n84 0.155672
R680 source.n101 source.n84 0.155672
R681 source.n101 source.n100 0.155672
R682 source.n100 source.n88 0.155672
R683 source.n93 source.n88 0.155672
R684 minus.n8 minus.t8 1342
R685 minus.n2 minus.t5 1342
R686 minus.n18 minus.t3 1342
R687 minus.n12 minus.t9 1342
R688 minus.n7 minus.t0 1282.12
R689 minus.n5 minus.t4 1282.12
R690 minus.n1 minus.t1 1282.12
R691 minus.n17 minus.t6 1282.12
R692 minus.n15 minus.t7 1282.12
R693 minus.n11 minus.t2 1282.12
R694 minus.n3 minus.n2 161.489
R695 minus.n13 minus.n12 161.489
R696 minus.n9 minus.n8 161.3
R697 minus.n6 minus.n0 161.3
R698 minus.n4 minus.n3 161.3
R699 minus.n19 minus.n18 161.3
R700 minus.n16 minus.n10 161.3
R701 minus.n14 minus.n13 161.3
R702 minus.n7 minus.n6 48.2005
R703 minus.n4 minus.n1 48.2005
R704 minus.n14 minus.n11 48.2005
R705 minus.n17 minus.n16 48.2005
R706 minus.n6 minus.n5 36.5157
R707 minus.n5 minus.n4 36.5157
R708 minus.n15 minus.n14 36.5157
R709 minus.n16 minus.n15 36.5157
R710 minus.n20 minus.n9 34.4854
R711 minus.n8 minus.n7 24.8308
R712 minus.n2 minus.n1 24.8308
R713 minus.n12 minus.n11 24.8308
R714 minus.n18 minus.n17 24.8308
R715 minus.n20 minus.n19 6.51565
R716 minus.n9 minus.n0 0.189894
R717 minus.n3 minus.n0 0.189894
R718 minus.n13 minus.n10 0.189894
R719 minus.n19 minus.n10 0.189894
R720 minus minus.n20 0.188
R721 drain_right.n60 drain_right.n0 289.615
R722 drain_right.n132 drain_right.n72 289.615
R723 drain_right.n20 drain_right.n19 185
R724 drain_right.n25 drain_right.n24 185
R725 drain_right.n27 drain_right.n26 185
R726 drain_right.n16 drain_right.n15 185
R727 drain_right.n33 drain_right.n32 185
R728 drain_right.n35 drain_right.n34 185
R729 drain_right.n12 drain_right.n11 185
R730 drain_right.n42 drain_right.n41 185
R731 drain_right.n43 drain_right.n10 185
R732 drain_right.n45 drain_right.n44 185
R733 drain_right.n8 drain_right.n7 185
R734 drain_right.n51 drain_right.n50 185
R735 drain_right.n53 drain_right.n52 185
R736 drain_right.n4 drain_right.n3 185
R737 drain_right.n59 drain_right.n58 185
R738 drain_right.n61 drain_right.n60 185
R739 drain_right.n133 drain_right.n132 185
R740 drain_right.n131 drain_right.n130 185
R741 drain_right.n76 drain_right.n75 185
R742 drain_right.n125 drain_right.n124 185
R743 drain_right.n123 drain_right.n122 185
R744 drain_right.n80 drain_right.n79 185
R745 drain_right.n117 drain_right.n116 185
R746 drain_right.n115 drain_right.n82 185
R747 drain_right.n114 drain_right.n113 185
R748 drain_right.n85 drain_right.n83 185
R749 drain_right.n108 drain_right.n107 185
R750 drain_right.n106 drain_right.n105 185
R751 drain_right.n89 drain_right.n88 185
R752 drain_right.n100 drain_right.n99 185
R753 drain_right.n98 drain_right.n97 185
R754 drain_right.n93 drain_right.n92 185
R755 drain_right.n21 drain_right.t0 149.524
R756 drain_right.n94 drain_right.t1 149.524
R757 drain_right.n25 drain_right.n19 104.615
R758 drain_right.n26 drain_right.n25 104.615
R759 drain_right.n26 drain_right.n15 104.615
R760 drain_right.n33 drain_right.n15 104.615
R761 drain_right.n34 drain_right.n33 104.615
R762 drain_right.n34 drain_right.n11 104.615
R763 drain_right.n42 drain_right.n11 104.615
R764 drain_right.n43 drain_right.n42 104.615
R765 drain_right.n44 drain_right.n43 104.615
R766 drain_right.n44 drain_right.n7 104.615
R767 drain_right.n51 drain_right.n7 104.615
R768 drain_right.n52 drain_right.n51 104.615
R769 drain_right.n52 drain_right.n3 104.615
R770 drain_right.n59 drain_right.n3 104.615
R771 drain_right.n60 drain_right.n59 104.615
R772 drain_right.n132 drain_right.n131 104.615
R773 drain_right.n131 drain_right.n75 104.615
R774 drain_right.n124 drain_right.n75 104.615
R775 drain_right.n124 drain_right.n123 104.615
R776 drain_right.n123 drain_right.n79 104.615
R777 drain_right.n116 drain_right.n79 104.615
R778 drain_right.n116 drain_right.n115 104.615
R779 drain_right.n115 drain_right.n114 104.615
R780 drain_right.n114 drain_right.n83 104.615
R781 drain_right.n107 drain_right.n83 104.615
R782 drain_right.n107 drain_right.n106 104.615
R783 drain_right.n106 drain_right.n88 104.615
R784 drain_right.n99 drain_right.n88 104.615
R785 drain_right.n99 drain_right.n98 104.615
R786 drain_right.n98 drain_right.n92 104.615
R787 drain_right.n71 drain_right.n69 60.0525
R788 drain_right.n68 drain_right.n67 59.8722
R789 drain_right.n71 drain_right.n70 59.5527
R790 drain_right.n66 drain_right.n65 59.5525
R791 drain_right.t0 drain_right.n19 52.3082
R792 drain_right.t1 drain_right.n92 52.3082
R793 drain_right.n66 drain_right.n64 47.0369
R794 drain_right.n137 drain_right.n136 46.5369
R795 drain_right drain_right.n68 28.9388
R796 drain_right.n45 drain_right.n10 13.1884
R797 drain_right.n117 drain_right.n82 13.1884
R798 drain_right.n41 drain_right.n40 12.8005
R799 drain_right.n46 drain_right.n8 12.8005
R800 drain_right.n118 drain_right.n80 12.8005
R801 drain_right.n113 drain_right.n84 12.8005
R802 drain_right.n39 drain_right.n12 12.0247
R803 drain_right.n50 drain_right.n49 12.0247
R804 drain_right.n122 drain_right.n121 12.0247
R805 drain_right.n112 drain_right.n85 12.0247
R806 drain_right.n36 drain_right.n35 11.249
R807 drain_right.n53 drain_right.n6 11.249
R808 drain_right.n125 drain_right.n78 11.249
R809 drain_right.n109 drain_right.n108 11.249
R810 drain_right.n32 drain_right.n14 10.4732
R811 drain_right.n54 drain_right.n4 10.4732
R812 drain_right.n126 drain_right.n76 10.4732
R813 drain_right.n105 drain_right.n87 10.4732
R814 drain_right.n21 drain_right.n20 10.2747
R815 drain_right.n94 drain_right.n93 10.2747
R816 drain_right.n31 drain_right.n16 9.69747
R817 drain_right.n58 drain_right.n57 9.69747
R818 drain_right.n130 drain_right.n129 9.69747
R819 drain_right.n104 drain_right.n89 9.69747
R820 drain_right.n64 drain_right.n63 9.45567
R821 drain_right.n136 drain_right.n135 9.45567
R822 drain_right.n63 drain_right.n62 9.3005
R823 drain_right.n2 drain_right.n1 9.3005
R824 drain_right.n57 drain_right.n56 9.3005
R825 drain_right.n55 drain_right.n54 9.3005
R826 drain_right.n6 drain_right.n5 9.3005
R827 drain_right.n49 drain_right.n48 9.3005
R828 drain_right.n47 drain_right.n46 9.3005
R829 drain_right.n23 drain_right.n22 9.3005
R830 drain_right.n18 drain_right.n17 9.3005
R831 drain_right.n29 drain_right.n28 9.3005
R832 drain_right.n31 drain_right.n30 9.3005
R833 drain_right.n14 drain_right.n13 9.3005
R834 drain_right.n37 drain_right.n36 9.3005
R835 drain_right.n39 drain_right.n38 9.3005
R836 drain_right.n40 drain_right.n9 9.3005
R837 drain_right.n96 drain_right.n95 9.3005
R838 drain_right.n91 drain_right.n90 9.3005
R839 drain_right.n102 drain_right.n101 9.3005
R840 drain_right.n104 drain_right.n103 9.3005
R841 drain_right.n87 drain_right.n86 9.3005
R842 drain_right.n110 drain_right.n109 9.3005
R843 drain_right.n112 drain_right.n111 9.3005
R844 drain_right.n84 drain_right.n81 9.3005
R845 drain_right.n135 drain_right.n134 9.3005
R846 drain_right.n74 drain_right.n73 9.3005
R847 drain_right.n129 drain_right.n128 9.3005
R848 drain_right.n127 drain_right.n126 9.3005
R849 drain_right.n78 drain_right.n77 9.3005
R850 drain_right.n121 drain_right.n120 9.3005
R851 drain_right.n119 drain_right.n118 9.3005
R852 drain_right.n28 drain_right.n27 8.92171
R853 drain_right.n61 drain_right.n2 8.92171
R854 drain_right.n133 drain_right.n74 8.92171
R855 drain_right.n101 drain_right.n100 8.92171
R856 drain_right.n24 drain_right.n18 8.14595
R857 drain_right.n62 drain_right.n0 8.14595
R858 drain_right.n134 drain_right.n72 8.14595
R859 drain_right.n97 drain_right.n91 8.14595
R860 drain_right.n23 drain_right.n20 7.3702
R861 drain_right.n96 drain_right.n93 7.3702
R862 drain_right drain_right.n137 5.90322
R863 drain_right.n24 drain_right.n23 5.81868
R864 drain_right.n64 drain_right.n0 5.81868
R865 drain_right.n136 drain_right.n72 5.81868
R866 drain_right.n97 drain_right.n96 5.81868
R867 drain_right.n27 drain_right.n18 5.04292
R868 drain_right.n62 drain_right.n61 5.04292
R869 drain_right.n134 drain_right.n133 5.04292
R870 drain_right.n100 drain_right.n91 5.04292
R871 drain_right.n28 drain_right.n16 4.26717
R872 drain_right.n58 drain_right.n2 4.26717
R873 drain_right.n130 drain_right.n74 4.26717
R874 drain_right.n101 drain_right.n89 4.26717
R875 drain_right.n32 drain_right.n31 3.49141
R876 drain_right.n57 drain_right.n4 3.49141
R877 drain_right.n129 drain_right.n76 3.49141
R878 drain_right.n105 drain_right.n104 3.49141
R879 drain_right.n22 drain_right.n21 2.84303
R880 drain_right.n95 drain_right.n94 2.84303
R881 drain_right.n35 drain_right.n14 2.71565
R882 drain_right.n54 drain_right.n53 2.71565
R883 drain_right.n126 drain_right.n125 2.71565
R884 drain_right.n108 drain_right.n87 2.71565
R885 drain_right.n36 drain_right.n12 1.93989
R886 drain_right.n50 drain_right.n6 1.93989
R887 drain_right.n122 drain_right.n78 1.93989
R888 drain_right.n109 drain_right.n85 1.93989
R889 drain_right.n67 drain_right.t3 1.6505
R890 drain_right.n67 drain_right.t6 1.6505
R891 drain_right.n65 drain_right.t7 1.6505
R892 drain_right.n65 drain_right.t2 1.6505
R893 drain_right.n69 drain_right.t8 1.6505
R894 drain_right.n69 drain_right.t4 1.6505
R895 drain_right.n70 drain_right.t9 1.6505
R896 drain_right.n70 drain_right.t5 1.6505
R897 drain_right.n41 drain_right.n39 1.16414
R898 drain_right.n49 drain_right.n8 1.16414
R899 drain_right.n121 drain_right.n80 1.16414
R900 drain_right.n113 drain_right.n112 1.16414
R901 drain_right.n137 drain_right.n71 0.5005
R902 drain_right.n40 drain_right.n10 0.388379
R903 drain_right.n46 drain_right.n45 0.388379
R904 drain_right.n118 drain_right.n117 0.388379
R905 drain_right.n84 drain_right.n82 0.388379
R906 drain_right.n22 drain_right.n17 0.155672
R907 drain_right.n29 drain_right.n17 0.155672
R908 drain_right.n30 drain_right.n29 0.155672
R909 drain_right.n30 drain_right.n13 0.155672
R910 drain_right.n37 drain_right.n13 0.155672
R911 drain_right.n38 drain_right.n37 0.155672
R912 drain_right.n38 drain_right.n9 0.155672
R913 drain_right.n47 drain_right.n9 0.155672
R914 drain_right.n48 drain_right.n47 0.155672
R915 drain_right.n48 drain_right.n5 0.155672
R916 drain_right.n55 drain_right.n5 0.155672
R917 drain_right.n56 drain_right.n55 0.155672
R918 drain_right.n56 drain_right.n1 0.155672
R919 drain_right.n63 drain_right.n1 0.155672
R920 drain_right.n135 drain_right.n73 0.155672
R921 drain_right.n128 drain_right.n73 0.155672
R922 drain_right.n128 drain_right.n127 0.155672
R923 drain_right.n127 drain_right.n77 0.155672
R924 drain_right.n120 drain_right.n77 0.155672
R925 drain_right.n120 drain_right.n119 0.155672
R926 drain_right.n119 drain_right.n81 0.155672
R927 drain_right.n111 drain_right.n81 0.155672
R928 drain_right.n111 drain_right.n110 0.155672
R929 drain_right.n110 drain_right.n86 0.155672
R930 drain_right.n103 drain_right.n86 0.155672
R931 drain_right.n103 drain_right.n102 0.155672
R932 drain_right.n102 drain_right.n90 0.155672
R933 drain_right.n95 drain_right.n90 0.155672
R934 drain_right.n68 drain_right.n66 0.070154
C0 source plus 3.1322f
C1 drain_left source 22.7654f
C2 minus drain_right 3.54847f
C3 source drain_right 22.753698f
C4 drain_left plus 3.67974f
C5 drain_right plus 0.290194f
C6 drain_left drain_right 0.693946f
C7 minus source 3.11749f
C8 minus plus 4.91006f
C9 minus drain_left 0.171039f
C10 drain_right a_n1412_n3288# 6.96601f
C11 drain_left a_n1412_n3288# 7.210929f
C12 source a_n1412_n3288# 6.033611f
C13 minus a_n1412_n3288# 5.44009f
C14 plus a_n1412_n3288# 7.47672f
C15 drain_right.n0 a_n1412_n3288# 0.041349f
C16 drain_right.n1 a_n1412_n3288# 0.031216f
C17 drain_right.n2 a_n1412_n3288# 0.016774f
C18 drain_right.n3 a_n1412_n3288# 0.039648f
C19 drain_right.n4 a_n1412_n3288# 0.017761f
C20 drain_right.n5 a_n1412_n3288# 0.031216f
C21 drain_right.n6 a_n1412_n3288# 0.016774f
C22 drain_right.n7 a_n1412_n3288# 0.039648f
C23 drain_right.n8 a_n1412_n3288# 0.017761f
C24 drain_right.n9 a_n1412_n3288# 0.031216f
C25 drain_right.n10 a_n1412_n3288# 0.017267f
C26 drain_right.n11 a_n1412_n3288# 0.039648f
C27 drain_right.n12 a_n1412_n3288# 0.017761f
C28 drain_right.n13 a_n1412_n3288# 0.031216f
C29 drain_right.n14 a_n1412_n3288# 0.016774f
C30 drain_right.n15 a_n1412_n3288# 0.039648f
C31 drain_right.n16 a_n1412_n3288# 0.017761f
C32 drain_right.n17 a_n1412_n3288# 0.031216f
C33 drain_right.n18 a_n1412_n3288# 0.016774f
C34 drain_right.n19 a_n1412_n3288# 0.029736f
C35 drain_right.n20 a_n1412_n3288# 0.028028f
C36 drain_right.t0 a_n1412_n3288# 0.066963f
C37 drain_right.n21 a_n1412_n3288# 0.225063f
C38 drain_right.n22 a_n1412_n3288# 1.57479f
C39 drain_right.n23 a_n1412_n3288# 0.016774f
C40 drain_right.n24 a_n1412_n3288# 0.017761f
C41 drain_right.n25 a_n1412_n3288# 0.039648f
C42 drain_right.n26 a_n1412_n3288# 0.039648f
C43 drain_right.n27 a_n1412_n3288# 0.017761f
C44 drain_right.n28 a_n1412_n3288# 0.016774f
C45 drain_right.n29 a_n1412_n3288# 0.031216f
C46 drain_right.n30 a_n1412_n3288# 0.031216f
C47 drain_right.n31 a_n1412_n3288# 0.016774f
C48 drain_right.n32 a_n1412_n3288# 0.017761f
C49 drain_right.n33 a_n1412_n3288# 0.039648f
C50 drain_right.n34 a_n1412_n3288# 0.039648f
C51 drain_right.n35 a_n1412_n3288# 0.017761f
C52 drain_right.n36 a_n1412_n3288# 0.016774f
C53 drain_right.n37 a_n1412_n3288# 0.031216f
C54 drain_right.n38 a_n1412_n3288# 0.031216f
C55 drain_right.n39 a_n1412_n3288# 0.016774f
C56 drain_right.n40 a_n1412_n3288# 0.016774f
C57 drain_right.n41 a_n1412_n3288# 0.017761f
C58 drain_right.n42 a_n1412_n3288# 0.039648f
C59 drain_right.n43 a_n1412_n3288# 0.039648f
C60 drain_right.n44 a_n1412_n3288# 0.039648f
C61 drain_right.n45 a_n1412_n3288# 0.017267f
C62 drain_right.n46 a_n1412_n3288# 0.016774f
C63 drain_right.n47 a_n1412_n3288# 0.031216f
C64 drain_right.n48 a_n1412_n3288# 0.031216f
C65 drain_right.n49 a_n1412_n3288# 0.016774f
C66 drain_right.n50 a_n1412_n3288# 0.017761f
C67 drain_right.n51 a_n1412_n3288# 0.039648f
C68 drain_right.n52 a_n1412_n3288# 0.039648f
C69 drain_right.n53 a_n1412_n3288# 0.017761f
C70 drain_right.n54 a_n1412_n3288# 0.016774f
C71 drain_right.n55 a_n1412_n3288# 0.031216f
C72 drain_right.n56 a_n1412_n3288# 0.031216f
C73 drain_right.n57 a_n1412_n3288# 0.016774f
C74 drain_right.n58 a_n1412_n3288# 0.017761f
C75 drain_right.n59 a_n1412_n3288# 0.039648f
C76 drain_right.n60 a_n1412_n3288# 0.081362f
C77 drain_right.n61 a_n1412_n3288# 0.017761f
C78 drain_right.n62 a_n1412_n3288# 0.016774f
C79 drain_right.n63 a_n1412_n3288# 0.067037f
C80 drain_right.n64 a_n1412_n3288# 0.067644f
C81 drain_right.t7 a_n1412_n3288# 0.296014f
C82 drain_right.t2 a_n1412_n3288# 0.296014f
C83 drain_right.n65 a_n1412_n3288# 2.63406f
C84 drain_right.n66 a_n1412_n3288# 0.436001f
C85 drain_right.t3 a_n1412_n3288# 0.296014f
C86 drain_right.t6 a_n1412_n3288# 0.296014f
C87 drain_right.n67 a_n1412_n3288# 2.63598f
C88 drain_right.n68 a_n1412_n3288# 1.67091f
C89 drain_right.t8 a_n1412_n3288# 0.296014f
C90 drain_right.t4 a_n1412_n3288# 0.296014f
C91 drain_right.n69 a_n1412_n3288# 2.63719f
C92 drain_right.t9 a_n1412_n3288# 0.296014f
C93 drain_right.t5 a_n1412_n3288# 0.296014f
C94 drain_right.n70 a_n1412_n3288# 2.63407f
C95 drain_right.n71 a_n1412_n3288# 0.734572f
C96 drain_right.n72 a_n1412_n3288# 0.041349f
C97 drain_right.n73 a_n1412_n3288# 0.031216f
C98 drain_right.n74 a_n1412_n3288# 0.016774f
C99 drain_right.n75 a_n1412_n3288# 0.039648f
C100 drain_right.n76 a_n1412_n3288# 0.017761f
C101 drain_right.n77 a_n1412_n3288# 0.031216f
C102 drain_right.n78 a_n1412_n3288# 0.016774f
C103 drain_right.n79 a_n1412_n3288# 0.039648f
C104 drain_right.n80 a_n1412_n3288# 0.017761f
C105 drain_right.n81 a_n1412_n3288# 0.031216f
C106 drain_right.n82 a_n1412_n3288# 0.017267f
C107 drain_right.n83 a_n1412_n3288# 0.039648f
C108 drain_right.n84 a_n1412_n3288# 0.016774f
C109 drain_right.n85 a_n1412_n3288# 0.017761f
C110 drain_right.n86 a_n1412_n3288# 0.031216f
C111 drain_right.n87 a_n1412_n3288# 0.016774f
C112 drain_right.n88 a_n1412_n3288# 0.039648f
C113 drain_right.n89 a_n1412_n3288# 0.017761f
C114 drain_right.n90 a_n1412_n3288# 0.031216f
C115 drain_right.n91 a_n1412_n3288# 0.016774f
C116 drain_right.n92 a_n1412_n3288# 0.029736f
C117 drain_right.n93 a_n1412_n3288# 0.028028f
C118 drain_right.t1 a_n1412_n3288# 0.066963f
C119 drain_right.n94 a_n1412_n3288# 0.225063f
C120 drain_right.n95 a_n1412_n3288# 1.57479f
C121 drain_right.n96 a_n1412_n3288# 0.016774f
C122 drain_right.n97 a_n1412_n3288# 0.017761f
C123 drain_right.n98 a_n1412_n3288# 0.039648f
C124 drain_right.n99 a_n1412_n3288# 0.039648f
C125 drain_right.n100 a_n1412_n3288# 0.017761f
C126 drain_right.n101 a_n1412_n3288# 0.016774f
C127 drain_right.n102 a_n1412_n3288# 0.031216f
C128 drain_right.n103 a_n1412_n3288# 0.031216f
C129 drain_right.n104 a_n1412_n3288# 0.016774f
C130 drain_right.n105 a_n1412_n3288# 0.017761f
C131 drain_right.n106 a_n1412_n3288# 0.039648f
C132 drain_right.n107 a_n1412_n3288# 0.039648f
C133 drain_right.n108 a_n1412_n3288# 0.017761f
C134 drain_right.n109 a_n1412_n3288# 0.016774f
C135 drain_right.n110 a_n1412_n3288# 0.031216f
C136 drain_right.n111 a_n1412_n3288# 0.031216f
C137 drain_right.n112 a_n1412_n3288# 0.016774f
C138 drain_right.n113 a_n1412_n3288# 0.017761f
C139 drain_right.n114 a_n1412_n3288# 0.039648f
C140 drain_right.n115 a_n1412_n3288# 0.039648f
C141 drain_right.n116 a_n1412_n3288# 0.039648f
C142 drain_right.n117 a_n1412_n3288# 0.017267f
C143 drain_right.n118 a_n1412_n3288# 0.016774f
C144 drain_right.n119 a_n1412_n3288# 0.031216f
C145 drain_right.n120 a_n1412_n3288# 0.031216f
C146 drain_right.n121 a_n1412_n3288# 0.016774f
C147 drain_right.n122 a_n1412_n3288# 0.017761f
C148 drain_right.n123 a_n1412_n3288# 0.039648f
C149 drain_right.n124 a_n1412_n3288# 0.039648f
C150 drain_right.n125 a_n1412_n3288# 0.017761f
C151 drain_right.n126 a_n1412_n3288# 0.016774f
C152 drain_right.n127 a_n1412_n3288# 0.031216f
C153 drain_right.n128 a_n1412_n3288# 0.031216f
C154 drain_right.n129 a_n1412_n3288# 0.016774f
C155 drain_right.n130 a_n1412_n3288# 0.017761f
C156 drain_right.n131 a_n1412_n3288# 0.039648f
C157 drain_right.n132 a_n1412_n3288# 0.081362f
C158 drain_right.n133 a_n1412_n3288# 0.017761f
C159 drain_right.n134 a_n1412_n3288# 0.016774f
C160 drain_right.n135 a_n1412_n3288# 0.067037f
C161 drain_right.n136 a_n1412_n3288# 0.066501f
C162 drain_right.n137 a_n1412_n3288# 0.364545f
C163 minus.n0 a_n1412_n3288# 0.055019f
C164 minus.t8 a_n1412_n3288# 0.475048f
C165 minus.t0 a_n1412_n3288# 0.466423f
C166 minus.t4 a_n1412_n3288# 0.466423f
C167 minus.t1 a_n1412_n3288# 0.466423f
C168 minus.n1 a_n1412_n3288# 0.187854f
C169 minus.t5 a_n1412_n3288# 0.475048f
C170 minus.n2 a_n1412_n3288# 0.205709f
C171 minus.n3 a_n1412_n3288# 0.129286f
C172 minus.n4 a_n1412_n3288# 0.020965f
C173 minus.n5 a_n1412_n3288# 0.187854f
C174 minus.n6 a_n1412_n3288# 0.020965f
C175 minus.n7 a_n1412_n3288# 0.187854f
C176 minus.n8 a_n1412_n3288# 0.205622f
C177 minus.n9 a_n1412_n3288# 1.8021f
C178 minus.n10 a_n1412_n3288# 0.055019f
C179 minus.t6 a_n1412_n3288# 0.466423f
C180 minus.t7 a_n1412_n3288# 0.466423f
C181 minus.t2 a_n1412_n3288# 0.466423f
C182 minus.n11 a_n1412_n3288# 0.187854f
C183 minus.t9 a_n1412_n3288# 0.475048f
C184 minus.n12 a_n1412_n3288# 0.205709f
C185 minus.n13 a_n1412_n3288# 0.129286f
C186 minus.n14 a_n1412_n3288# 0.020965f
C187 minus.n15 a_n1412_n3288# 0.187854f
C188 minus.n16 a_n1412_n3288# 0.020965f
C189 minus.n17 a_n1412_n3288# 0.187854f
C190 minus.t3 a_n1412_n3288# 0.475048f
C191 minus.n18 a_n1412_n3288# 0.205622f
C192 minus.n19 a_n1412_n3288# 0.361728f
C193 minus.n20 a_n1412_n3288# 2.19905f
C194 source.n0 a_n1412_n3288# 0.042722f
C195 source.n1 a_n1412_n3288# 0.032252f
C196 source.n2 a_n1412_n3288# 0.017331f
C197 source.n3 a_n1412_n3288# 0.040964f
C198 source.n4 a_n1412_n3288# 0.01835f
C199 source.n5 a_n1412_n3288# 0.032252f
C200 source.n6 a_n1412_n3288# 0.017331f
C201 source.n7 a_n1412_n3288# 0.040964f
C202 source.n8 a_n1412_n3288# 0.01835f
C203 source.n9 a_n1412_n3288# 0.032252f
C204 source.n10 a_n1412_n3288# 0.01784f
C205 source.n11 a_n1412_n3288# 0.040964f
C206 source.n12 a_n1412_n3288# 0.017331f
C207 source.n13 a_n1412_n3288# 0.01835f
C208 source.n14 a_n1412_n3288# 0.032252f
C209 source.n15 a_n1412_n3288# 0.017331f
C210 source.n16 a_n1412_n3288# 0.040964f
C211 source.n17 a_n1412_n3288# 0.01835f
C212 source.n18 a_n1412_n3288# 0.032252f
C213 source.n19 a_n1412_n3288# 0.017331f
C214 source.n20 a_n1412_n3288# 0.030723f
C215 source.n21 a_n1412_n3288# 0.028958f
C216 source.t13 a_n1412_n3288# 0.069185f
C217 source.n22 a_n1412_n3288# 0.232533f
C218 source.n23 a_n1412_n3288# 1.62706f
C219 source.n24 a_n1412_n3288# 0.017331f
C220 source.n25 a_n1412_n3288# 0.01835f
C221 source.n26 a_n1412_n3288# 0.040964f
C222 source.n27 a_n1412_n3288# 0.040964f
C223 source.n28 a_n1412_n3288# 0.01835f
C224 source.n29 a_n1412_n3288# 0.017331f
C225 source.n30 a_n1412_n3288# 0.032252f
C226 source.n31 a_n1412_n3288# 0.032252f
C227 source.n32 a_n1412_n3288# 0.017331f
C228 source.n33 a_n1412_n3288# 0.01835f
C229 source.n34 a_n1412_n3288# 0.040964f
C230 source.n35 a_n1412_n3288# 0.040964f
C231 source.n36 a_n1412_n3288# 0.01835f
C232 source.n37 a_n1412_n3288# 0.017331f
C233 source.n38 a_n1412_n3288# 0.032252f
C234 source.n39 a_n1412_n3288# 0.032252f
C235 source.n40 a_n1412_n3288# 0.017331f
C236 source.n41 a_n1412_n3288# 0.01835f
C237 source.n42 a_n1412_n3288# 0.040964f
C238 source.n43 a_n1412_n3288# 0.040964f
C239 source.n44 a_n1412_n3288# 0.040964f
C240 source.n45 a_n1412_n3288# 0.01784f
C241 source.n46 a_n1412_n3288# 0.017331f
C242 source.n47 a_n1412_n3288# 0.032252f
C243 source.n48 a_n1412_n3288# 0.032252f
C244 source.n49 a_n1412_n3288# 0.017331f
C245 source.n50 a_n1412_n3288# 0.01835f
C246 source.n51 a_n1412_n3288# 0.040964f
C247 source.n52 a_n1412_n3288# 0.040964f
C248 source.n53 a_n1412_n3288# 0.01835f
C249 source.n54 a_n1412_n3288# 0.017331f
C250 source.n55 a_n1412_n3288# 0.032252f
C251 source.n56 a_n1412_n3288# 0.032252f
C252 source.n57 a_n1412_n3288# 0.017331f
C253 source.n58 a_n1412_n3288# 0.01835f
C254 source.n59 a_n1412_n3288# 0.040964f
C255 source.n60 a_n1412_n3288# 0.084062f
C256 source.n61 a_n1412_n3288# 0.01835f
C257 source.n62 a_n1412_n3288# 0.017331f
C258 source.n63 a_n1412_n3288# 0.069262f
C259 source.n64 a_n1412_n3288# 0.046393f
C260 source.n65 a_n1412_n3288# 1.29063f
C261 source.t12 a_n1412_n3288# 0.305838f
C262 source.t18 a_n1412_n3288# 0.305838f
C263 source.n66 a_n1412_n3288# 2.61859f
C264 source.n67 a_n1412_n3288# 0.433658f
C265 source.t15 a_n1412_n3288# 0.305838f
C266 source.t17 a_n1412_n3288# 0.305838f
C267 source.n68 a_n1412_n3288# 2.61859f
C268 source.n69 a_n1412_n3288# 0.456504f
C269 source.n70 a_n1412_n3288# 0.042722f
C270 source.n71 a_n1412_n3288# 0.032252f
C271 source.n72 a_n1412_n3288# 0.017331f
C272 source.n73 a_n1412_n3288# 0.040964f
C273 source.n74 a_n1412_n3288# 0.01835f
C274 source.n75 a_n1412_n3288# 0.032252f
C275 source.n76 a_n1412_n3288# 0.017331f
C276 source.n77 a_n1412_n3288# 0.040964f
C277 source.n78 a_n1412_n3288# 0.01835f
C278 source.n79 a_n1412_n3288# 0.032252f
C279 source.n80 a_n1412_n3288# 0.01784f
C280 source.n81 a_n1412_n3288# 0.040964f
C281 source.n82 a_n1412_n3288# 0.017331f
C282 source.n83 a_n1412_n3288# 0.01835f
C283 source.n84 a_n1412_n3288# 0.032252f
C284 source.n85 a_n1412_n3288# 0.017331f
C285 source.n86 a_n1412_n3288# 0.040964f
C286 source.n87 a_n1412_n3288# 0.01835f
C287 source.n88 a_n1412_n3288# 0.032252f
C288 source.n89 a_n1412_n3288# 0.017331f
C289 source.n90 a_n1412_n3288# 0.030723f
C290 source.n91 a_n1412_n3288# 0.028958f
C291 source.t1 a_n1412_n3288# 0.069185f
C292 source.n92 a_n1412_n3288# 0.232533f
C293 source.n93 a_n1412_n3288# 1.62706f
C294 source.n94 a_n1412_n3288# 0.017331f
C295 source.n95 a_n1412_n3288# 0.01835f
C296 source.n96 a_n1412_n3288# 0.040964f
C297 source.n97 a_n1412_n3288# 0.040964f
C298 source.n98 a_n1412_n3288# 0.01835f
C299 source.n99 a_n1412_n3288# 0.017331f
C300 source.n100 a_n1412_n3288# 0.032252f
C301 source.n101 a_n1412_n3288# 0.032252f
C302 source.n102 a_n1412_n3288# 0.017331f
C303 source.n103 a_n1412_n3288# 0.01835f
C304 source.n104 a_n1412_n3288# 0.040964f
C305 source.n105 a_n1412_n3288# 0.040964f
C306 source.n106 a_n1412_n3288# 0.01835f
C307 source.n107 a_n1412_n3288# 0.017331f
C308 source.n108 a_n1412_n3288# 0.032252f
C309 source.n109 a_n1412_n3288# 0.032252f
C310 source.n110 a_n1412_n3288# 0.017331f
C311 source.n111 a_n1412_n3288# 0.01835f
C312 source.n112 a_n1412_n3288# 0.040964f
C313 source.n113 a_n1412_n3288# 0.040964f
C314 source.n114 a_n1412_n3288# 0.040964f
C315 source.n115 a_n1412_n3288# 0.01784f
C316 source.n116 a_n1412_n3288# 0.017331f
C317 source.n117 a_n1412_n3288# 0.032252f
C318 source.n118 a_n1412_n3288# 0.032252f
C319 source.n119 a_n1412_n3288# 0.017331f
C320 source.n120 a_n1412_n3288# 0.01835f
C321 source.n121 a_n1412_n3288# 0.040964f
C322 source.n122 a_n1412_n3288# 0.040964f
C323 source.n123 a_n1412_n3288# 0.01835f
C324 source.n124 a_n1412_n3288# 0.017331f
C325 source.n125 a_n1412_n3288# 0.032252f
C326 source.n126 a_n1412_n3288# 0.032252f
C327 source.n127 a_n1412_n3288# 0.017331f
C328 source.n128 a_n1412_n3288# 0.01835f
C329 source.n129 a_n1412_n3288# 0.040964f
C330 source.n130 a_n1412_n3288# 0.084062f
C331 source.n131 a_n1412_n3288# 0.01835f
C332 source.n132 a_n1412_n3288# 0.017331f
C333 source.n133 a_n1412_n3288# 0.069262f
C334 source.n134 a_n1412_n3288# 0.046393f
C335 source.n135 a_n1412_n3288# 0.151335f
C336 source.t8 a_n1412_n3288# 0.305838f
C337 source.t0 a_n1412_n3288# 0.305838f
C338 source.n136 a_n1412_n3288# 2.61859f
C339 source.n137 a_n1412_n3288# 0.433658f
C340 source.t6 a_n1412_n3288# 0.305838f
C341 source.t4 a_n1412_n3288# 0.305838f
C342 source.n138 a_n1412_n3288# 2.61859f
C343 source.n139 a_n1412_n3288# 2.15329f
C344 source.t16 a_n1412_n3288# 0.305838f
C345 source.t9 a_n1412_n3288# 0.305838f
C346 source.n140 a_n1412_n3288# 2.61857f
C347 source.n141 a_n1412_n3288# 2.1533f
C348 source.t14 a_n1412_n3288# 0.305838f
C349 source.t11 a_n1412_n3288# 0.305838f
C350 source.n142 a_n1412_n3288# 2.61857f
C351 source.n143 a_n1412_n3288# 0.433674f
C352 source.n144 a_n1412_n3288# 0.042722f
C353 source.n145 a_n1412_n3288# 0.032252f
C354 source.n146 a_n1412_n3288# 0.017331f
C355 source.n147 a_n1412_n3288# 0.040964f
C356 source.n148 a_n1412_n3288# 0.01835f
C357 source.n149 a_n1412_n3288# 0.032252f
C358 source.n150 a_n1412_n3288# 0.017331f
C359 source.n151 a_n1412_n3288# 0.040964f
C360 source.n152 a_n1412_n3288# 0.01835f
C361 source.n153 a_n1412_n3288# 0.032252f
C362 source.n154 a_n1412_n3288# 0.01784f
C363 source.n155 a_n1412_n3288# 0.040964f
C364 source.n156 a_n1412_n3288# 0.01835f
C365 source.n157 a_n1412_n3288# 0.032252f
C366 source.n158 a_n1412_n3288# 0.017331f
C367 source.n159 a_n1412_n3288# 0.040964f
C368 source.n160 a_n1412_n3288# 0.01835f
C369 source.n161 a_n1412_n3288# 0.032252f
C370 source.n162 a_n1412_n3288# 0.017331f
C371 source.n163 a_n1412_n3288# 0.030723f
C372 source.n164 a_n1412_n3288# 0.028958f
C373 source.t10 a_n1412_n3288# 0.069185f
C374 source.n165 a_n1412_n3288# 0.232533f
C375 source.n166 a_n1412_n3288# 1.62706f
C376 source.n167 a_n1412_n3288# 0.017331f
C377 source.n168 a_n1412_n3288# 0.01835f
C378 source.n169 a_n1412_n3288# 0.040964f
C379 source.n170 a_n1412_n3288# 0.040964f
C380 source.n171 a_n1412_n3288# 0.01835f
C381 source.n172 a_n1412_n3288# 0.017331f
C382 source.n173 a_n1412_n3288# 0.032252f
C383 source.n174 a_n1412_n3288# 0.032252f
C384 source.n175 a_n1412_n3288# 0.017331f
C385 source.n176 a_n1412_n3288# 0.01835f
C386 source.n177 a_n1412_n3288# 0.040964f
C387 source.n178 a_n1412_n3288# 0.040964f
C388 source.n179 a_n1412_n3288# 0.01835f
C389 source.n180 a_n1412_n3288# 0.017331f
C390 source.n181 a_n1412_n3288# 0.032252f
C391 source.n182 a_n1412_n3288# 0.032252f
C392 source.n183 a_n1412_n3288# 0.017331f
C393 source.n184 a_n1412_n3288# 0.017331f
C394 source.n185 a_n1412_n3288# 0.01835f
C395 source.n186 a_n1412_n3288# 0.040964f
C396 source.n187 a_n1412_n3288# 0.040964f
C397 source.n188 a_n1412_n3288# 0.040964f
C398 source.n189 a_n1412_n3288# 0.01784f
C399 source.n190 a_n1412_n3288# 0.017331f
C400 source.n191 a_n1412_n3288# 0.032252f
C401 source.n192 a_n1412_n3288# 0.032252f
C402 source.n193 a_n1412_n3288# 0.017331f
C403 source.n194 a_n1412_n3288# 0.01835f
C404 source.n195 a_n1412_n3288# 0.040964f
C405 source.n196 a_n1412_n3288# 0.040964f
C406 source.n197 a_n1412_n3288# 0.01835f
C407 source.n198 a_n1412_n3288# 0.017331f
C408 source.n199 a_n1412_n3288# 0.032252f
C409 source.n200 a_n1412_n3288# 0.032252f
C410 source.n201 a_n1412_n3288# 0.017331f
C411 source.n202 a_n1412_n3288# 0.01835f
C412 source.n203 a_n1412_n3288# 0.040964f
C413 source.n204 a_n1412_n3288# 0.084062f
C414 source.n205 a_n1412_n3288# 0.01835f
C415 source.n206 a_n1412_n3288# 0.017331f
C416 source.n207 a_n1412_n3288# 0.069262f
C417 source.n208 a_n1412_n3288# 0.046393f
C418 source.n209 a_n1412_n3288# 0.151335f
C419 source.t19 a_n1412_n3288# 0.305838f
C420 source.t3 a_n1412_n3288# 0.305838f
C421 source.n210 a_n1412_n3288# 2.61857f
C422 source.n211 a_n1412_n3288# 0.45652f
C423 source.t7 a_n1412_n3288# 0.305838f
C424 source.t5 a_n1412_n3288# 0.305838f
C425 source.n212 a_n1412_n3288# 2.61857f
C426 source.n213 a_n1412_n3288# 0.433674f
C427 source.n214 a_n1412_n3288# 0.042722f
C428 source.n215 a_n1412_n3288# 0.032252f
C429 source.n216 a_n1412_n3288# 0.017331f
C430 source.n217 a_n1412_n3288# 0.040964f
C431 source.n218 a_n1412_n3288# 0.01835f
C432 source.n219 a_n1412_n3288# 0.032252f
C433 source.n220 a_n1412_n3288# 0.017331f
C434 source.n221 a_n1412_n3288# 0.040964f
C435 source.n222 a_n1412_n3288# 0.01835f
C436 source.n223 a_n1412_n3288# 0.032252f
C437 source.n224 a_n1412_n3288# 0.01784f
C438 source.n225 a_n1412_n3288# 0.040964f
C439 source.n226 a_n1412_n3288# 0.01835f
C440 source.n227 a_n1412_n3288# 0.032252f
C441 source.n228 a_n1412_n3288# 0.017331f
C442 source.n229 a_n1412_n3288# 0.040964f
C443 source.n230 a_n1412_n3288# 0.01835f
C444 source.n231 a_n1412_n3288# 0.032252f
C445 source.n232 a_n1412_n3288# 0.017331f
C446 source.n233 a_n1412_n3288# 0.030723f
C447 source.n234 a_n1412_n3288# 0.028958f
C448 source.t2 a_n1412_n3288# 0.069185f
C449 source.n235 a_n1412_n3288# 0.232533f
C450 source.n236 a_n1412_n3288# 1.62706f
C451 source.n237 a_n1412_n3288# 0.017331f
C452 source.n238 a_n1412_n3288# 0.01835f
C453 source.n239 a_n1412_n3288# 0.040964f
C454 source.n240 a_n1412_n3288# 0.040964f
C455 source.n241 a_n1412_n3288# 0.01835f
C456 source.n242 a_n1412_n3288# 0.017331f
C457 source.n243 a_n1412_n3288# 0.032252f
C458 source.n244 a_n1412_n3288# 0.032252f
C459 source.n245 a_n1412_n3288# 0.017331f
C460 source.n246 a_n1412_n3288# 0.01835f
C461 source.n247 a_n1412_n3288# 0.040964f
C462 source.n248 a_n1412_n3288# 0.040964f
C463 source.n249 a_n1412_n3288# 0.01835f
C464 source.n250 a_n1412_n3288# 0.017331f
C465 source.n251 a_n1412_n3288# 0.032252f
C466 source.n252 a_n1412_n3288# 0.032252f
C467 source.n253 a_n1412_n3288# 0.017331f
C468 source.n254 a_n1412_n3288# 0.017331f
C469 source.n255 a_n1412_n3288# 0.01835f
C470 source.n256 a_n1412_n3288# 0.040964f
C471 source.n257 a_n1412_n3288# 0.040964f
C472 source.n258 a_n1412_n3288# 0.040964f
C473 source.n259 a_n1412_n3288# 0.01784f
C474 source.n260 a_n1412_n3288# 0.017331f
C475 source.n261 a_n1412_n3288# 0.032252f
C476 source.n262 a_n1412_n3288# 0.032252f
C477 source.n263 a_n1412_n3288# 0.017331f
C478 source.n264 a_n1412_n3288# 0.01835f
C479 source.n265 a_n1412_n3288# 0.040964f
C480 source.n266 a_n1412_n3288# 0.040964f
C481 source.n267 a_n1412_n3288# 0.01835f
C482 source.n268 a_n1412_n3288# 0.017331f
C483 source.n269 a_n1412_n3288# 0.032252f
C484 source.n270 a_n1412_n3288# 0.032252f
C485 source.n271 a_n1412_n3288# 0.017331f
C486 source.n272 a_n1412_n3288# 0.01835f
C487 source.n273 a_n1412_n3288# 0.040964f
C488 source.n274 a_n1412_n3288# 0.084062f
C489 source.n275 a_n1412_n3288# 0.01835f
C490 source.n276 a_n1412_n3288# 0.017331f
C491 source.n277 a_n1412_n3288# 0.069262f
C492 source.n278 a_n1412_n3288# 0.046393f
C493 source.n279 a_n1412_n3288# 0.303831f
C494 source.n280 a_n1412_n3288# 2.02079f
C495 drain_left.n0 a_n1412_n3288# 0.041471f
C496 drain_left.n1 a_n1412_n3288# 0.031308f
C497 drain_left.n2 a_n1412_n3288# 0.016824f
C498 drain_left.n3 a_n1412_n3288# 0.039765f
C499 drain_left.n4 a_n1412_n3288# 0.017813f
C500 drain_left.n5 a_n1412_n3288# 0.031308f
C501 drain_left.n6 a_n1412_n3288# 0.016824f
C502 drain_left.n7 a_n1412_n3288# 0.039765f
C503 drain_left.n8 a_n1412_n3288# 0.017813f
C504 drain_left.n9 a_n1412_n3288# 0.031308f
C505 drain_left.n10 a_n1412_n3288# 0.017318f
C506 drain_left.n11 a_n1412_n3288# 0.039765f
C507 drain_left.n12 a_n1412_n3288# 0.017813f
C508 drain_left.n13 a_n1412_n3288# 0.031308f
C509 drain_left.n14 a_n1412_n3288# 0.016824f
C510 drain_left.n15 a_n1412_n3288# 0.039765f
C511 drain_left.n16 a_n1412_n3288# 0.017813f
C512 drain_left.n17 a_n1412_n3288# 0.031308f
C513 drain_left.n18 a_n1412_n3288# 0.016824f
C514 drain_left.n19 a_n1412_n3288# 0.029824f
C515 drain_left.n20 a_n1412_n3288# 0.028111f
C516 drain_left.t5 a_n1412_n3288# 0.06716f
C517 drain_left.n21 a_n1412_n3288# 0.225727f
C518 drain_left.n22 a_n1412_n3288# 1.57943f
C519 drain_left.n23 a_n1412_n3288# 0.016824f
C520 drain_left.n24 a_n1412_n3288# 0.017813f
C521 drain_left.n25 a_n1412_n3288# 0.039765f
C522 drain_left.n26 a_n1412_n3288# 0.039765f
C523 drain_left.n27 a_n1412_n3288# 0.017813f
C524 drain_left.n28 a_n1412_n3288# 0.016824f
C525 drain_left.n29 a_n1412_n3288# 0.031308f
C526 drain_left.n30 a_n1412_n3288# 0.031308f
C527 drain_left.n31 a_n1412_n3288# 0.016824f
C528 drain_left.n32 a_n1412_n3288# 0.017813f
C529 drain_left.n33 a_n1412_n3288# 0.039765f
C530 drain_left.n34 a_n1412_n3288# 0.039765f
C531 drain_left.n35 a_n1412_n3288# 0.017813f
C532 drain_left.n36 a_n1412_n3288# 0.016824f
C533 drain_left.n37 a_n1412_n3288# 0.031308f
C534 drain_left.n38 a_n1412_n3288# 0.031308f
C535 drain_left.n39 a_n1412_n3288# 0.016824f
C536 drain_left.n40 a_n1412_n3288# 0.016824f
C537 drain_left.n41 a_n1412_n3288# 0.017813f
C538 drain_left.n42 a_n1412_n3288# 0.039765f
C539 drain_left.n43 a_n1412_n3288# 0.039765f
C540 drain_left.n44 a_n1412_n3288# 0.039765f
C541 drain_left.n45 a_n1412_n3288# 0.017318f
C542 drain_left.n46 a_n1412_n3288# 0.016824f
C543 drain_left.n47 a_n1412_n3288# 0.031308f
C544 drain_left.n48 a_n1412_n3288# 0.031308f
C545 drain_left.n49 a_n1412_n3288# 0.016824f
C546 drain_left.n50 a_n1412_n3288# 0.017813f
C547 drain_left.n51 a_n1412_n3288# 0.039765f
C548 drain_left.n52 a_n1412_n3288# 0.039765f
C549 drain_left.n53 a_n1412_n3288# 0.017813f
C550 drain_left.n54 a_n1412_n3288# 0.016824f
C551 drain_left.n55 a_n1412_n3288# 0.031308f
C552 drain_left.n56 a_n1412_n3288# 0.031308f
C553 drain_left.n57 a_n1412_n3288# 0.016824f
C554 drain_left.n58 a_n1412_n3288# 0.017813f
C555 drain_left.n59 a_n1412_n3288# 0.039765f
C556 drain_left.n60 a_n1412_n3288# 0.081602f
C557 drain_left.n61 a_n1412_n3288# 0.017813f
C558 drain_left.n62 a_n1412_n3288# 0.016824f
C559 drain_left.n63 a_n1412_n3288# 0.067234f
C560 drain_left.n64 a_n1412_n3288# 0.067843f
C561 drain_left.t3 a_n1412_n3288# 0.296886f
C562 drain_left.t1 a_n1412_n3288# 0.296886f
C563 drain_left.n65 a_n1412_n3288# 2.64183f
C564 drain_left.n66 a_n1412_n3288# 0.437287f
C565 drain_left.t7 a_n1412_n3288# 0.296886f
C566 drain_left.t4 a_n1412_n3288# 0.296886f
C567 drain_left.n67 a_n1412_n3288# 2.64375f
C568 drain_left.n68 a_n1412_n3288# 1.74129f
C569 drain_left.n69 a_n1412_n3288# 0.041471f
C570 drain_left.n70 a_n1412_n3288# 0.031308f
C571 drain_left.n71 a_n1412_n3288# 0.016824f
C572 drain_left.n72 a_n1412_n3288# 0.039765f
C573 drain_left.n73 a_n1412_n3288# 0.017813f
C574 drain_left.n74 a_n1412_n3288# 0.031308f
C575 drain_left.n75 a_n1412_n3288# 0.016824f
C576 drain_left.n76 a_n1412_n3288# 0.039765f
C577 drain_left.n77 a_n1412_n3288# 0.017813f
C578 drain_left.n78 a_n1412_n3288# 0.031308f
C579 drain_left.n79 a_n1412_n3288# 0.017318f
C580 drain_left.n80 a_n1412_n3288# 0.039765f
C581 drain_left.n81 a_n1412_n3288# 0.016824f
C582 drain_left.n82 a_n1412_n3288# 0.017813f
C583 drain_left.n83 a_n1412_n3288# 0.031308f
C584 drain_left.n84 a_n1412_n3288# 0.016824f
C585 drain_left.n85 a_n1412_n3288# 0.039765f
C586 drain_left.n86 a_n1412_n3288# 0.017813f
C587 drain_left.n87 a_n1412_n3288# 0.031308f
C588 drain_left.n88 a_n1412_n3288# 0.016824f
C589 drain_left.n89 a_n1412_n3288# 0.029824f
C590 drain_left.n90 a_n1412_n3288# 0.028111f
C591 drain_left.t6 a_n1412_n3288# 0.06716f
C592 drain_left.n91 a_n1412_n3288# 0.225727f
C593 drain_left.n92 a_n1412_n3288# 1.57943f
C594 drain_left.n93 a_n1412_n3288# 0.016824f
C595 drain_left.n94 a_n1412_n3288# 0.017813f
C596 drain_left.n95 a_n1412_n3288# 0.039765f
C597 drain_left.n96 a_n1412_n3288# 0.039765f
C598 drain_left.n97 a_n1412_n3288# 0.017813f
C599 drain_left.n98 a_n1412_n3288# 0.016824f
C600 drain_left.n99 a_n1412_n3288# 0.031308f
C601 drain_left.n100 a_n1412_n3288# 0.031308f
C602 drain_left.n101 a_n1412_n3288# 0.016824f
C603 drain_left.n102 a_n1412_n3288# 0.017813f
C604 drain_left.n103 a_n1412_n3288# 0.039765f
C605 drain_left.n104 a_n1412_n3288# 0.039765f
C606 drain_left.n105 a_n1412_n3288# 0.017813f
C607 drain_left.n106 a_n1412_n3288# 0.016824f
C608 drain_left.n107 a_n1412_n3288# 0.031308f
C609 drain_left.n108 a_n1412_n3288# 0.031308f
C610 drain_left.n109 a_n1412_n3288# 0.016824f
C611 drain_left.n110 a_n1412_n3288# 0.017813f
C612 drain_left.n111 a_n1412_n3288# 0.039765f
C613 drain_left.n112 a_n1412_n3288# 0.039765f
C614 drain_left.n113 a_n1412_n3288# 0.039765f
C615 drain_left.n114 a_n1412_n3288# 0.017318f
C616 drain_left.n115 a_n1412_n3288# 0.016824f
C617 drain_left.n116 a_n1412_n3288# 0.031308f
C618 drain_left.n117 a_n1412_n3288# 0.031308f
C619 drain_left.n118 a_n1412_n3288# 0.016824f
C620 drain_left.n119 a_n1412_n3288# 0.017813f
C621 drain_left.n120 a_n1412_n3288# 0.039765f
C622 drain_left.n121 a_n1412_n3288# 0.039765f
C623 drain_left.n122 a_n1412_n3288# 0.017813f
C624 drain_left.n123 a_n1412_n3288# 0.016824f
C625 drain_left.n124 a_n1412_n3288# 0.031308f
C626 drain_left.n125 a_n1412_n3288# 0.031308f
C627 drain_left.n126 a_n1412_n3288# 0.016824f
C628 drain_left.n127 a_n1412_n3288# 0.017813f
C629 drain_left.n128 a_n1412_n3288# 0.039765f
C630 drain_left.n129 a_n1412_n3288# 0.081602f
C631 drain_left.n130 a_n1412_n3288# 0.017813f
C632 drain_left.n131 a_n1412_n3288# 0.016824f
C633 drain_left.n132 a_n1412_n3288# 0.067234f
C634 drain_left.n133 a_n1412_n3288# 0.067843f
C635 drain_left.t9 a_n1412_n3288# 0.296886f
C636 drain_left.t0 a_n1412_n3288# 0.296886f
C637 drain_left.n134 a_n1412_n3288# 2.64184f
C638 drain_left.n135 a_n1412_n3288# 0.470269f
C639 drain_left.t8 a_n1412_n3288# 0.296886f
C640 drain_left.t2 a_n1412_n3288# 0.296886f
C641 drain_left.n136 a_n1412_n3288# 2.64183f
C642 drain_left.n137 a_n1412_n3288# 0.622061f
C643 plus.n0 a_n1412_n3288# 0.056523f
C644 plus.t0 a_n1412_n3288# 0.479171f
C645 plus.t6 a_n1412_n3288# 0.479171f
C646 plus.t1 a_n1412_n3288# 0.479171f
C647 plus.n1 a_n1412_n3288# 0.192988f
C648 plus.t3 a_n1412_n3288# 0.488031f
C649 plus.n2 a_n1412_n3288# 0.211331f
C650 plus.n3 a_n1412_n3288# 0.13282f
C651 plus.n4 a_n1412_n3288# 0.021538f
C652 plus.n5 a_n1412_n3288# 0.192988f
C653 plus.n6 a_n1412_n3288# 0.021538f
C654 plus.n7 a_n1412_n3288# 0.192988f
C655 plus.t5 a_n1412_n3288# 0.488031f
C656 plus.n8 a_n1412_n3288# 0.211242f
C657 plus.n9 a_n1412_n3288# 0.634519f
C658 plus.n10 a_n1412_n3288# 0.056523f
C659 plus.t2 a_n1412_n3288# 0.488031f
C660 plus.t9 a_n1412_n3288# 0.479171f
C661 plus.t4 a_n1412_n3288# 0.479171f
C662 plus.t7 a_n1412_n3288# 0.479171f
C663 plus.n11 a_n1412_n3288# 0.192988f
C664 plus.t8 a_n1412_n3288# 0.488031f
C665 plus.n12 a_n1412_n3288# 0.211331f
C666 plus.n13 a_n1412_n3288# 0.13282f
C667 plus.n14 a_n1412_n3288# 0.021538f
C668 plus.n15 a_n1412_n3288# 0.192988f
C669 plus.n16 a_n1412_n3288# 0.021538f
C670 plus.n17 a_n1412_n3288# 0.192988f
C671 plus.n18 a_n1412_n3288# 0.211242f
C672 plus.n19 a_n1412_n3288# 1.56088f
.ends

