* NGSPICE file created from diffpair316.ext - technology: sky130A

.subckt diffpair316 minus drain_right drain_left source plus
X0 source.t24 plus.t0 drain_left.t0 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X1 source.t5 minus.t0 drain_right.t13 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X2 drain_left.t12 plus.t1 source.t23 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X3 a_n2524_n2088# a_n2524_n2088# a_n2524_n2088# a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.8
X4 a_n2524_n2088# a_n2524_n2088# a_n2524_n2088# a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X5 drain_left.t3 plus.t2 source.t22 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X6 drain_left.t13 plus.t3 source.t21 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X7 drain_right.t12 minus.t1 source.t1 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X8 drain_right.t11 minus.t2 source.t8 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X9 drain_right.t10 minus.t3 source.t10 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X10 drain_left.t7 plus.t4 source.t20 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X11 drain_right.t9 minus.t4 source.t9 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X12 source.t2 minus.t5 drain_right.t8 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X13 drain_right.t7 minus.t6 source.t6 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X14 drain_right.t6 minus.t7 source.t7 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X15 source.t19 plus.t5 drain_left.t8 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X16 drain_right.t5 minus.t8 source.t0 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X17 source.t3 minus.t9 drain_right.t4 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X18 source.t25 minus.t10 drain_right.t3 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X19 a_n2524_n2088# a_n2524_n2088# a_n2524_n2088# a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X20 drain_right.t2 minus.t11 source.t26 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X21 drain_left.t9 plus.t6 source.t18 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.8
X22 source.t17 plus.t7 drain_left.t10 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X23 source.t16 plus.t8 drain_left.t1 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X24 drain_left.t4 plus.t9 source.t15 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X25 a_n2524_n2088# a_n2524_n2088# a_n2524_n2088# a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.8
X26 source.t27 minus.t12 drain_right.t1 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X27 drain_left.t2 plus.t10 source.t14 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X28 source.t13 plus.t11 drain_left.t6 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X29 drain_left.t11 plus.t12 source.t12 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.8
X30 source.t4 minus.t13 drain_right.t0 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
X31 source.t11 plus.t13 drain_left.t5 a_n2524_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.8
R0 plus.n5 plus.t12 253.701
R1 plus.n23 plus.t4 253.701
R2 plus.n16 plus.t6 229.855
R3 plus.n14 plus.t7 229.855
R4 plus.n2 plus.t10 229.855
R5 plus.n9 plus.t8 229.855
R6 plus.n8 plus.t9 229.855
R7 plus.n4 plus.t11 229.855
R8 plus.n34 plus.t1 229.855
R9 plus.n32 plus.t5 229.855
R10 plus.n20 plus.t3 229.855
R11 plus.n27 plus.t13 229.855
R12 plus.n26 plus.t2 229.855
R13 plus.n22 plus.t0 229.855
R14 plus.n7 plus.n6 161.3
R15 plus.n13 plus.n12 161.3
R16 plus.n14 plus.n1 161.3
R17 plus.n15 plus.n0 161.3
R18 plus.n17 plus.n16 161.3
R19 plus.n25 plus.n24 161.3
R20 plus.n31 plus.n30 161.3
R21 plus.n32 plus.n19 161.3
R22 plus.n33 plus.n18 161.3
R23 plus.n35 plus.n34 161.3
R24 plus.n8 plus.n3 80.6037
R25 plus.n10 plus.n9 80.6037
R26 plus.n11 plus.n2 80.6037
R27 plus.n26 plus.n21 80.6037
R28 plus.n28 plus.n27 80.6037
R29 plus.n29 plus.n20 80.6037
R30 plus.n9 plus.n2 48.2005
R31 plus.n9 plus.n8 48.2005
R32 plus.n27 plus.n20 48.2005
R33 plus.n27 plus.n26 48.2005
R34 plus.n24 plus.n23 44.9119
R35 plus.n6 plus.n5 44.9119
R36 plus.n16 plus.n15 35.055
R37 plus.n34 plus.n33 35.055
R38 plus.n13 plus.n2 32.1338
R39 plus.n8 plus.n7 32.1338
R40 plus.n31 plus.n20 32.1338
R41 plus.n26 plus.n25 32.1338
R42 plus plus.n35 30.5161
R43 plus.n23 plus.n22 17.739
R44 plus.n5 plus.n4 17.739
R45 plus.n14 plus.n13 16.0672
R46 plus.n7 plus.n4 16.0672
R47 plus.n32 plus.n31 16.0672
R48 plus.n25 plus.n22 16.0672
R49 plus.n15 plus.n14 13.146
R50 plus.n33 plus.n32 13.146
R51 plus plus.n17 10.0971
R52 plus.n10 plus.n3 0.380177
R53 plus.n11 plus.n10 0.380177
R54 plus.n29 plus.n28 0.380177
R55 plus.n28 plus.n21 0.380177
R56 plus.n6 plus.n3 0.285035
R57 plus.n12 plus.n11 0.285035
R58 plus.n30 plus.n29 0.285035
R59 plus.n24 plus.n21 0.285035
R60 plus.n12 plus.n1 0.189894
R61 plus.n1 plus.n0 0.189894
R62 plus.n17 plus.n0 0.189894
R63 plus.n35 plus.n18 0.189894
R64 plus.n19 plus.n18 0.189894
R65 plus.n30 plus.n19 0.189894
R66 drain_left.n26 drain_left.n0 289.615
R67 drain_left.n63 drain_left.n37 289.615
R68 drain_left.n11 drain_left.n10 185
R69 drain_left.n8 drain_left.n7 185
R70 drain_left.n17 drain_left.n16 185
R71 drain_left.n19 drain_left.n18 185
R72 drain_left.n4 drain_left.n3 185
R73 drain_left.n25 drain_left.n24 185
R74 drain_left.n27 drain_left.n26 185
R75 drain_left.n64 drain_left.n63 185
R76 drain_left.n62 drain_left.n61 185
R77 drain_left.n41 drain_left.n40 185
R78 drain_left.n56 drain_left.n55 185
R79 drain_left.n54 drain_left.n53 185
R80 drain_left.n45 drain_left.n44 185
R81 drain_left.n48 drain_left.n47 185
R82 drain_left.t12 drain_left.n9 147.661
R83 drain_left.t11 drain_left.n46 147.661
R84 drain_left.n10 drain_left.n7 104.615
R85 drain_left.n17 drain_left.n7 104.615
R86 drain_left.n18 drain_left.n17 104.615
R87 drain_left.n18 drain_left.n3 104.615
R88 drain_left.n25 drain_left.n3 104.615
R89 drain_left.n26 drain_left.n25 104.615
R90 drain_left.n63 drain_left.n62 104.615
R91 drain_left.n62 drain_left.n40 104.615
R92 drain_left.n55 drain_left.n40 104.615
R93 drain_left.n55 drain_left.n54 104.615
R94 drain_left.n54 drain_left.n44 104.615
R95 drain_left.n47 drain_left.n44 104.615
R96 drain_left.n35 drain_left.n33 68.1648
R97 drain_left.n71 drain_left.n70 67.1908
R98 drain_left.n69 drain_left.n68 67.1908
R99 drain_left.n73 drain_left.n72 67.1907
R100 drain_left.n35 drain_left.n34 67.1907
R101 drain_left.n32 drain_left.n31 67.1907
R102 drain_left.n10 drain_left.t12 52.3082
R103 drain_left.n47 drain_left.t11 52.3082
R104 drain_left.n32 drain_left.n30 49.8383
R105 drain_left.n69 drain_left.n67 49.8383
R106 drain_left drain_left.n36 28.4229
R107 drain_left.n11 drain_left.n9 15.6674
R108 drain_left.n48 drain_left.n46 15.6674
R109 drain_left.n12 drain_left.n8 12.8005
R110 drain_left.n49 drain_left.n45 12.8005
R111 drain_left.n16 drain_left.n15 12.0247
R112 drain_left.n53 drain_left.n52 12.0247
R113 drain_left.n19 drain_left.n6 11.249
R114 drain_left.n56 drain_left.n43 11.249
R115 drain_left.n20 drain_left.n4 10.4732
R116 drain_left.n57 drain_left.n41 10.4732
R117 drain_left.n24 drain_left.n23 9.69747
R118 drain_left.n61 drain_left.n60 9.69747
R119 drain_left.n30 drain_left.n29 9.45567
R120 drain_left.n67 drain_left.n66 9.45567
R121 drain_left.n29 drain_left.n28 9.3005
R122 drain_left.n2 drain_left.n1 9.3005
R123 drain_left.n23 drain_left.n22 9.3005
R124 drain_left.n21 drain_left.n20 9.3005
R125 drain_left.n6 drain_left.n5 9.3005
R126 drain_left.n15 drain_left.n14 9.3005
R127 drain_left.n13 drain_left.n12 9.3005
R128 drain_left.n66 drain_left.n65 9.3005
R129 drain_left.n39 drain_left.n38 9.3005
R130 drain_left.n60 drain_left.n59 9.3005
R131 drain_left.n58 drain_left.n57 9.3005
R132 drain_left.n43 drain_left.n42 9.3005
R133 drain_left.n52 drain_left.n51 9.3005
R134 drain_left.n50 drain_left.n49 9.3005
R135 drain_left.n27 drain_left.n2 8.92171
R136 drain_left.n64 drain_left.n39 8.92171
R137 drain_left.n28 drain_left.n0 8.14595
R138 drain_left.n65 drain_left.n37 8.14595
R139 drain_left drain_left.n73 6.62735
R140 drain_left.n30 drain_left.n0 5.81868
R141 drain_left.n67 drain_left.n37 5.81868
R142 drain_left.n28 drain_left.n27 5.04292
R143 drain_left.n65 drain_left.n64 5.04292
R144 drain_left.n13 drain_left.n9 4.38594
R145 drain_left.n50 drain_left.n46 4.38594
R146 drain_left.n24 drain_left.n2 4.26717
R147 drain_left.n61 drain_left.n39 4.26717
R148 drain_left.n23 drain_left.n4 3.49141
R149 drain_left.n60 drain_left.n41 3.49141
R150 drain_left.n33 drain_left.t0 3.3005
R151 drain_left.n33 drain_left.t7 3.3005
R152 drain_left.n34 drain_left.t5 3.3005
R153 drain_left.n34 drain_left.t3 3.3005
R154 drain_left.n31 drain_left.t8 3.3005
R155 drain_left.n31 drain_left.t13 3.3005
R156 drain_left.n72 drain_left.t10 3.3005
R157 drain_left.n72 drain_left.t9 3.3005
R158 drain_left.n70 drain_left.t1 3.3005
R159 drain_left.n70 drain_left.t2 3.3005
R160 drain_left.n68 drain_left.t6 3.3005
R161 drain_left.n68 drain_left.t4 3.3005
R162 drain_left.n20 drain_left.n19 2.71565
R163 drain_left.n57 drain_left.n56 2.71565
R164 drain_left.n16 drain_left.n6 1.93989
R165 drain_left.n53 drain_left.n43 1.93989
R166 drain_left.n15 drain_left.n8 1.16414
R167 drain_left.n52 drain_left.n45 1.16414
R168 drain_left.n71 drain_left.n69 0.974638
R169 drain_left.n73 drain_left.n71 0.974638
R170 drain_left.n36 drain_left.n32 0.675757
R171 drain_left.n12 drain_left.n11 0.388379
R172 drain_left.n49 drain_left.n48 0.388379
R173 drain_left.n36 drain_left.n35 0.188688
R174 drain_left.n14 drain_left.n13 0.155672
R175 drain_left.n14 drain_left.n5 0.155672
R176 drain_left.n21 drain_left.n5 0.155672
R177 drain_left.n22 drain_left.n21 0.155672
R178 drain_left.n22 drain_left.n1 0.155672
R179 drain_left.n29 drain_left.n1 0.155672
R180 drain_left.n66 drain_left.n38 0.155672
R181 drain_left.n59 drain_left.n38 0.155672
R182 drain_left.n59 drain_left.n58 0.155672
R183 drain_left.n58 drain_left.n42 0.155672
R184 drain_left.n51 drain_left.n42 0.155672
R185 drain_left.n51 drain_left.n50 0.155672
R186 source.n146 source.n120 289.615
R187 source.n108 source.n82 289.615
R188 source.n26 source.n0 289.615
R189 source.n64 source.n38 289.615
R190 source.n131 source.n130 185
R191 source.n128 source.n127 185
R192 source.n137 source.n136 185
R193 source.n139 source.n138 185
R194 source.n124 source.n123 185
R195 source.n145 source.n144 185
R196 source.n147 source.n146 185
R197 source.n93 source.n92 185
R198 source.n90 source.n89 185
R199 source.n99 source.n98 185
R200 source.n101 source.n100 185
R201 source.n86 source.n85 185
R202 source.n107 source.n106 185
R203 source.n109 source.n108 185
R204 source.n27 source.n26 185
R205 source.n25 source.n24 185
R206 source.n4 source.n3 185
R207 source.n19 source.n18 185
R208 source.n17 source.n16 185
R209 source.n8 source.n7 185
R210 source.n11 source.n10 185
R211 source.n65 source.n64 185
R212 source.n63 source.n62 185
R213 source.n42 source.n41 185
R214 source.n57 source.n56 185
R215 source.n55 source.n54 185
R216 source.n46 source.n45 185
R217 source.n49 source.n48 185
R218 source.t1 source.n129 147.661
R219 source.t20 source.n91 147.661
R220 source.t18 source.n9 147.661
R221 source.t0 source.n47 147.661
R222 source.n130 source.n127 104.615
R223 source.n137 source.n127 104.615
R224 source.n138 source.n137 104.615
R225 source.n138 source.n123 104.615
R226 source.n145 source.n123 104.615
R227 source.n146 source.n145 104.615
R228 source.n92 source.n89 104.615
R229 source.n99 source.n89 104.615
R230 source.n100 source.n99 104.615
R231 source.n100 source.n85 104.615
R232 source.n107 source.n85 104.615
R233 source.n108 source.n107 104.615
R234 source.n26 source.n25 104.615
R235 source.n25 source.n3 104.615
R236 source.n18 source.n3 104.615
R237 source.n18 source.n17 104.615
R238 source.n17 source.n7 104.615
R239 source.n10 source.n7 104.615
R240 source.n64 source.n63 104.615
R241 source.n63 source.n41 104.615
R242 source.n56 source.n41 104.615
R243 source.n56 source.n55 104.615
R244 source.n55 source.n45 104.615
R245 source.n48 source.n45 104.615
R246 source.n130 source.t1 52.3082
R247 source.n92 source.t20 52.3082
R248 source.n10 source.t18 52.3082
R249 source.n48 source.t0 52.3082
R250 source.n33 source.n32 50.512
R251 source.n35 source.n34 50.512
R252 source.n37 source.n36 50.512
R253 source.n71 source.n70 50.512
R254 source.n73 source.n72 50.512
R255 source.n75 source.n74 50.512
R256 source.n119 source.n118 50.5119
R257 source.n117 source.n116 50.5119
R258 source.n115 source.n114 50.5119
R259 source.n81 source.n80 50.5119
R260 source.n79 source.n78 50.5119
R261 source.n77 source.n76 50.5119
R262 source.n151 source.n150 32.1853
R263 source.n113 source.n112 32.1853
R264 source.n31 source.n30 32.1853
R265 source.n69 source.n68 32.1853
R266 source.n77 source.n75 18.6905
R267 source.n131 source.n129 15.6674
R268 source.n93 source.n91 15.6674
R269 source.n11 source.n9 15.6674
R270 source.n49 source.n47 15.6674
R271 source.n132 source.n128 12.8005
R272 source.n94 source.n90 12.8005
R273 source.n12 source.n8 12.8005
R274 source.n50 source.n46 12.8005
R275 source.n136 source.n135 12.0247
R276 source.n98 source.n97 12.0247
R277 source.n16 source.n15 12.0247
R278 source.n54 source.n53 12.0247
R279 source.n152 source.n31 11.9664
R280 source.n139 source.n126 11.249
R281 source.n101 source.n88 11.249
R282 source.n19 source.n6 11.249
R283 source.n57 source.n44 11.249
R284 source.n140 source.n124 10.4732
R285 source.n102 source.n86 10.4732
R286 source.n20 source.n4 10.4732
R287 source.n58 source.n42 10.4732
R288 source.n144 source.n143 9.69747
R289 source.n106 source.n105 9.69747
R290 source.n24 source.n23 9.69747
R291 source.n62 source.n61 9.69747
R292 source.n150 source.n149 9.45567
R293 source.n112 source.n111 9.45567
R294 source.n30 source.n29 9.45567
R295 source.n68 source.n67 9.45567
R296 source.n149 source.n148 9.3005
R297 source.n122 source.n121 9.3005
R298 source.n143 source.n142 9.3005
R299 source.n141 source.n140 9.3005
R300 source.n126 source.n125 9.3005
R301 source.n135 source.n134 9.3005
R302 source.n133 source.n132 9.3005
R303 source.n111 source.n110 9.3005
R304 source.n84 source.n83 9.3005
R305 source.n105 source.n104 9.3005
R306 source.n103 source.n102 9.3005
R307 source.n88 source.n87 9.3005
R308 source.n97 source.n96 9.3005
R309 source.n95 source.n94 9.3005
R310 source.n29 source.n28 9.3005
R311 source.n2 source.n1 9.3005
R312 source.n23 source.n22 9.3005
R313 source.n21 source.n20 9.3005
R314 source.n6 source.n5 9.3005
R315 source.n15 source.n14 9.3005
R316 source.n13 source.n12 9.3005
R317 source.n67 source.n66 9.3005
R318 source.n40 source.n39 9.3005
R319 source.n61 source.n60 9.3005
R320 source.n59 source.n58 9.3005
R321 source.n44 source.n43 9.3005
R322 source.n53 source.n52 9.3005
R323 source.n51 source.n50 9.3005
R324 source.n147 source.n122 8.92171
R325 source.n109 source.n84 8.92171
R326 source.n27 source.n2 8.92171
R327 source.n65 source.n40 8.92171
R328 source.n148 source.n120 8.14595
R329 source.n110 source.n82 8.14595
R330 source.n28 source.n0 8.14595
R331 source.n66 source.n38 8.14595
R332 source.n150 source.n120 5.81868
R333 source.n112 source.n82 5.81868
R334 source.n30 source.n0 5.81868
R335 source.n68 source.n38 5.81868
R336 source.n152 source.n151 5.7505
R337 source.n148 source.n147 5.04292
R338 source.n110 source.n109 5.04292
R339 source.n28 source.n27 5.04292
R340 source.n66 source.n65 5.04292
R341 source.n133 source.n129 4.38594
R342 source.n95 source.n91 4.38594
R343 source.n13 source.n9 4.38594
R344 source.n51 source.n47 4.38594
R345 source.n144 source.n122 4.26717
R346 source.n106 source.n84 4.26717
R347 source.n24 source.n2 4.26717
R348 source.n62 source.n40 4.26717
R349 source.n143 source.n124 3.49141
R350 source.n105 source.n86 3.49141
R351 source.n23 source.n4 3.49141
R352 source.n61 source.n42 3.49141
R353 source.n118 source.t9 3.3005
R354 source.n118 source.t27 3.3005
R355 source.n116 source.t8 3.3005
R356 source.n116 source.t4 3.3005
R357 source.n114 source.t7 3.3005
R358 source.n114 source.t5 3.3005
R359 source.n80 source.t22 3.3005
R360 source.n80 source.t24 3.3005
R361 source.n78 source.t21 3.3005
R362 source.n78 source.t11 3.3005
R363 source.n76 source.t23 3.3005
R364 source.n76 source.t19 3.3005
R365 source.n32 source.t14 3.3005
R366 source.n32 source.t17 3.3005
R367 source.n34 source.t15 3.3005
R368 source.n34 source.t16 3.3005
R369 source.n36 source.t12 3.3005
R370 source.n36 source.t13 3.3005
R371 source.n70 source.t10 3.3005
R372 source.n70 source.t2 3.3005
R373 source.n72 source.t26 3.3005
R374 source.n72 source.t25 3.3005
R375 source.n74 source.t6 3.3005
R376 source.n74 source.t3 3.3005
R377 source.n140 source.n139 2.71565
R378 source.n102 source.n101 2.71565
R379 source.n20 source.n19 2.71565
R380 source.n58 source.n57 2.71565
R381 source.n136 source.n126 1.93989
R382 source.n98 source.n88 1.93989
R383 source.n16 source.n6 1.93989
R384 source.n54 source.n44 1.93989
R385 source.n135 source.n128 1.16414
R386 source.n97 source.n90 1.16414
R387 source.n15 source.n8 1.16414
R388 source.n53 source.n46 1.16414
R389 source.n75 source.n73 0.974638
R390 source.n73 source.n71 0.974638
R391 source.n71 source.n69 0.974638
R392 source.n37 source.n35 0.974638
R393 source.n35 source.n33 0.974638
R394 source.n33 source.n31 0.974638
R395 source.n79 source.n77 0.974638
R396 source.n81 source.n79 0.974638
R397 source.n113 source.n81 0.974638
R398 source.n117 source.n115 0.974638
R399 source.n119 source.n117 0.974638
R400 source.n151 source.n119 0.974638
R401 source.n69 source.n37 0.957397
R402 source.n115 source.n113 0.957397
R403 source.n132 source.n131 0.388379
R404 source.n94 source.n93 0.388379
R405 source.n12 source.n11 0.388379
R406 source.n50 source.n49 0.388379
R407 source source.n152 0.188
R408 source.n134 source.n133 0.155672
R409 source.n134 source.n125 0.155672
R410 source.n141 source.n125 0.155672
R411 source.n142 source.n141 0.155672
R412 source.n142 source.n121 0.155672
R413 source.n149 source.n121 0.155672
R414 source.n96 source.n95 0.155672
R415 source.n96 source.n87 0.155672
R416 source.n103 source.n87 0.155672
R417 source.n104 source.n103 0.155672
R418 source.n104 source.n83 0.155672
R419 source.n111 source.n83 0.155672
R420 source.n29 source.n1 0.155672
R421 source.n22 source.n1 0.155672
R422 source.n22 source.n21 0.155672
R423 source.n21 source.n5 0.155672
R424 source.n14 source.n5 0.155672
R425 source.n14 source.n13 0.155672
R426 source.n67 source.n39 0.155672
R427 source.n60 source.n39 0.155672
R428 source.n60 source.n59 0.155672
R429 source.n59 source.n43 0.155672
R430 source.n52 source.n43 0.155672
R431 source.n52 source.n51 0.155672
R432 minus.n5 minus.t8 253.701
R433 minus.n23 minus.t7 253.701
R434 minus.n4 minus.t5 229.855
R435 minus.n8 minus.t3 229.855
R436 minus.n9 minus.t10 229.855
R437 minus.n10 minus.t11 229.855
R438 minus.n14 minus.t9 229.855
R439 minus.n16 minus.t6 229.855
R440 minus.n22 minus.t0 229.855
R441 minus.n26 minus.t2 229.855
R442 minus.n27 minus.t13 229.855
R443 minus.n28 minus.t4 229.855
R444 minus.n32 minus.t12 229.855
R445 minus.n34 minus.t1 229.855
R446 minus.n17 minus.n16 161.3
R447 minus.n15 minus.n0 161.3
R448 minus.n14 minus.n13 161.3
R449 minus.n12 minus.n1 161.3
R450 minus.n6 minus.n3 161.3
R451 minus.n35 minus.n34 161.3
R452 minus.n33 minus.n18 161.3
R453 minus.n32 minus.n31 161.3
R454 minus.n30 minus.n19 161.3
R455 minus.n24 minus.n21 161.3
R456 minus.n11 minus.n10 80.6037
R457 minus.n9 minus.n2 80.6037
R458 minus.n8 minus.n7 80.6037
R459 minus.n29 minus.n28 80.6037
R460 minus.n27 minus.n20 80.6037
R461 minus.n26 minus.n25 80.6037
R462 minus.n9 minus.n8 48.2005
R463 minus.n10 minus.n9 48.2005
R464 minus.n27 minus.n26 48.2005
R465 minus.n28 minus.n27 48.2005
R466 minus.n6 minus.n5 44.9119
R467 minus.n24 minus.n23 44.9119
R468 minus.n16 minus.n15 35.055
R469 minus.n34 minus.n33 35.055
R470 minus.n36 minus.n17 34.3622
R471 minus.n8 minus.n3 32.1338
R472 minus.n10 minus.n1 32.1338
R473 minus.n26 minus.n21 32.1338
R474 minus.n28 minus.n19 32.1338
R475 minus.n5 minus.n4 17.739
R476 minus.n23 minus.n22 17.739
R477 minus.n4 minus.n3 16.0672
R478 minus.n14 minus.n1 16.0672
R479 minus.n22 minus.n21 16.0672
R480 minus.n32 minus.n19 16.0672
R481 minus.n15 minus.n14 13.146
R482 minus.n33 minus.n32 13.146
R483 minus.n36 minus.n35 6.72588
R484 minus.n11 minus.n2 0.380177
R485 minus.n7 minus.n2 0.380177
R486 minus.n25 minus.n20 0.380177
R487 minus.n29 minus.n20 0.380177
R488 minus.n12 minus.n11 0.285035
R489 minus.n7 minus.n6 0.285035
R490 minus.n25 minus.n24 0.285035
R491 minus.n30 minus.n29 0.285035
R492 minus.n17 minus.n0 0.189894
R493 minus.n13 minus.n0 0.189894
R494 minus.n13 minus.n12 0.189894
R495 minus.n31 minus.n30 0.189894
R496 minus.n31 minus.n18 0.189894
R497 minus.n35 minus.n18 0.189894
R498 minus minus.n36 0.188
R499 drain_right.n26 drain_right.n0 289.615
R500 drain_right.n68 drain_right.n42 289.615
R501 drain_right.n11 drain_right.n10 185
R502 drain_right.n8 drain_right.n7 185
R503 drain_right.n17 drain_right.n16 185
R504 drain_right.n19 drain_right.n18 185
R505 drain_right.n4 drain_right.n3 185
R506 drain_right.n25 drain_right.n24 185
R507 drain_right.n27 drain_right.n26 185
R508 drain_right.n69 drain_right.n68 185
R509 drain_right.n67 drain_right.n66 185
R510 drain_right.n46 drain_right.n45 185
R511 drain_right.n61 drain_right.n60 185
R512 drain_right.n59 drain_right.n58 185
R513 drain_right.n50 drain_right.n49 185
R514 drain_right.n53 drain_right.n52 185
R515 drain_right.t6 drain_right.n9 147.661
R516 drain_right.t7 drain_right.n51 147.661
R517 drain_right.n10 drain_right.n7 104.615
R518 drain_right.n17 drain_right.n7 104.615
R519 drain_right.n18 drain_right.n17 104.615
R520 drain_right.n18 drain_right.n3 104.615
R521 drain_right.n25 drain_right.n3 104.615
R522 drain_right.n26 drain_right.n25 104.615
R523 drain_right.n68 drain_right.n67 104.615
R524 drain_right.n67 drain_right.n45 104.615
R525 drain_right.n60 drain_right.n45 104.615
R526 drain_right.n60 drain_right.n59 104.615
R527 drain_right.n59 drain_right.n49 104.615
R528 drain_right.n52 drain_right.n49 104.615
R529 drain_right.n35 drain_right.n33 68.1648
R530 drain_right.n39 drain_right.n37 68.1648
R531 drain_right.n39 drain_right.n38 67.1908
R532 drain_right.n41 drain_right.n40 67.1908
R533 drain_right.n35 drain_right.n34 67.1907
R534 drain_right.n32 drain_right.n31 67.1907
R535 drain_right.n10 drain_right.t6 52.3082
R536 drain_right.n52 drain_right.t7 52.3082
R537 drain_right.n32 drain_right.n30 49.8383
R538 drain_right.n73 drain_right.n72 48.8641
R539 drain_right drain_right.n36 27.8697
R540 drain_right.n11 drain_right.n9 15.6674
R541 drain_right.n53 drain_right.n51 15.6674
R542 drain_right.n12 drain_right.n8 12.8005
R543 drain_right.n54 drain_right.n50 12.8005
R544 drain_right.n16 drain_right.n15 12.0247
R545 drain_right.n58 drain_right.n57 12.0247
R546 drain_right.n19 drain_right.n6 11.249
R547 drain_right.n61 drain_right.n48 11.249
R548 drain_right.n20 drain_right.n4 10.4732
R549 drain_right.n62 drain_right.n46 10.4732
R550 drain_right.n24 drain_right.n23 9.69747
R551 drain_right.n66 drain_right.n65 9.69747
R552 drain_right.n30 drain_right.n29 9.45567
R553 drain_right.n72 drain_right.n71 9.45567
R554 drain_right.n29 drain_right.n28 9.3005
R555 drain_right.n2 drain_right.n1 9.3005
R556 drain_right.n23 drain_right.n22 9.3005
R557 drain_right.n21 drain_right.n20 9.3005
R558 drain_right.n6 drain_right.n5 9.3005
R559 drain_right.n15 drain_right.n14 9.3005
R560 drain_right.n13 drain_right.n12 9.3005
R561 drain_right.n71 drain_right.n70 9.3005
R562 drain_right.n44 drain_right.n43 9.3005
R563 drain_right.n65 drain_right.n64 9.3005
R564 drain_right.n63 drain_right.n62 9.3005
R565 drain_right.n48 drain_right.n47 9.3005
R566 drain_right.n57 drain_right.n56 9.3005
R567 drain_right.n55 drain_right.n54 9.3005
R568 drain_right.n27 drain_right.n2 8.92171
R569 drain_right.n69 drain_right.n44 8.92171
R570 drain_right.n28 drain_right.n0 8.14595
R571 drain_right.n70 drain_right.n42 8.14595
R572 drain_right drain_right.n73 6.14028
R573 drain_right.n30 drain_right.n0 5.81868
R574 drain_right.n72 drain_right.n42 5.81868
R575 drain_right.n28 drain_right.n27 5.04292
R576 drain_right.n70 drain_right.n69 5.04292
R577 drain_right.n13 drain_right.n9 4.38594
R578 drain_right.n55 drain_right.n51 4.38594
R579 drain_right.n24 drain_right.n2 4.26717
R580 drain_right.n66 drain_right.n44 4.26717
R581 drain_right.n23 drain_right.n4 3.49141
R582 drain_right.n65 drain_right.n46 3.49141
R583 drain_right.n33 drain_right.t1 3.3005
R584 drain_right.n33 drain_right.t12 3.3005
R585 drain_right.n34 drain_right.t0 3.3005
R586 drain_right.n34 drain_right.t9 3.3005
R587 drain_right.n31 drain_right.t13 3.3005
R588 drain_right.n31 drain_right.t11 3.3005
R589 drain_right.n37 drain_right.t8 3.3005
R590 drain_right.n37 drain_right.t5 3.3005
R591 drain_right.n38 drain_right.t3 3.3005
R592 drain_right.n38 drain_right.t10 3.3005
R593 drain_right.n40 drain_right.t4 3.3005
R594 drain_right.n40 drain_right.t2 3.3005
R595 drain_right.n20 drain_right.n19 2.71565
R596 drain_right.n62 drain_right.n61 2.71565
R597 drain_right.n16 drain_right.n6 1.93989
R598 drain_right.n58 drain_right.n48 1.93989
R599 drain_right.n15 drain_right.n8 1.16414
R600 drain_right.n57 drain_right.n50 1.16414
R601 drain_right.n73 drain_right.n41 0.974638
R602 drain_right.n41 drain_right.n39 0.974638
R603 drain_right.n36 drain_right.n32 0.675757
R604 drain_right.n12 drain_right.n11 0.388379
R605 drain_right.n54 drain_right.n53 0.388379
R606 drain_right.n36 drain_right.n35 0.188688
R607 drain_right.n14 drain_right.n13 0.155672
R608 drain_right.n14 drain_right.n5 0.155672
R609 drain_right.n21 drain_right.n5 0.155672
R610 drain_right.n22 drain_right.n21 0.155672
R611 drain_right.n22 drain_right.n1 0.155672
R612 drain_right.n29 drain_right.n1 0.155672
R613 drain_right.n71 drain_right.n43 0.155672
R614 drain_right.n64 drain_right.n43 0.155672
R615 drain_right.n64 drain_right.n63 0.155672
R616 drain_right.n63 drain_right.n47 0.155672
R617 drain_right.n56 drain_right.n47 0.155672
R618 drain_right.n56 drain_right.n55 0.155672
C0 source plus 5.515069f
C1 minus plus 5.17554f
C2 source drain_left 10.461401f
C3 minus drain_left 0.173289f
C4 source drain_right 10.459599f
C5 minus drain_right 5.13693f
C6 source minus 5.50081f
C7 plus drain_left 5.38563f
C8 plus drain_right 0.407427f
C9 drain_right drain_left 1.31523f
C10 drain_right a_n2524_n2088# 6.02339f
C11 drain_left a_n2524_n2088# 6.40957f
C12 source a_n2524_n2088# 4.380037f
C13 minus a_n2524_n2088# 9.516173f
C14 plus a_n2524_n2088# 10.936979f
C15 drain_right.n0 a_n2524_n2088# 0.034468f
C16 drain_right.n1 a_n2524_n2088# 0.024522f
C17 drain_right.n2 a_n2524_n2088# 0.013177f
C18 drain_right.n3 a_n2524_n2088# 0.031146f
C19 drain_right.n4 a_n2524_n2088# 0.013952f
C20 drain_right.n5 a_n2524_n2088# 0.024522f
C21 drain_right.n6 a_n2524_n2088# 0.013177f
C22 drain_right.n7 a_n2524_n2088# 0.031146f
C23 drain_right.n8 a_n2524_n2088# 0.013952f
C24 drain_right.n9 a_n2524_n2088# 0.104939f
C25 drain_right.t6 a_n2524_n2088# 0.050765f
C26 drain_right.n10 a_n2524_n2088# 0.02336f
C27 drain_right.n11 a_n2524_n2088# 0.018398f
C28 drain_right.n12 a_n2524_n2088# 0.013177f
C29 drain_right.n13 a_n2524_n2088# 0.583488f
C30 drain_right.n14 a_n2524_n2088# 0.024522f
C31 drain_right.n15 a_n2524_n2088# 0.013177f
C32 drain_right.n16 a_n2524_n2088# 0.013952f
C33 drain_right.n17 a_n2524_n2088# 0.031146f
C34 drain_right.n18 a_n2524_n2088# 0.031146f
C35 drain_right.n19 a_n2524_n2088# 0.013952f
C36 drain_right.n20 a_n2524_n2088# 0.013177f
C37 drain_right.n21 a_n2524_n2088# 0.024522f
C38 drain_right.n22 a_n2524_n2088# 0.024522f
C39 drain_right.n23 a_n2524_n2088# 0.013177f
C40 drain_right.n24 a_n2524_n2088# 0.013952f
C41 drain_right.n25 a_n2524_n2088# 0.031146f
C42 drain_right.n26 a_n2524_n2088# 0.067426f
C43 drain_right.n27 a_n2524_n2088# 0.013952f
C44 drain_right.n28 a_n2524_n2088# 0.013177f
C45 drain_right.n29 a_n2524_n2088# 0.056682f
C46 drain_right.n30 a_n2524_n2088# 0.057087f
C47 drain_right.t13 a_n2524_n2088# 0.11627f
C48 drain_right.t11 a_n2524_n2088# 0.11627f
C49 drain_right.n31 a_n2524_n2088# 0.969695f
C50 drain_right.n32 a_n2524_n2088# 0.45197f
C51 drain_right.t1 a_n2524_n2088# 0.11627f
C52 drain_right.t12 a_n2524_n2088# 0.11627f
C53 drain_right.n33 a_n2524_n2088# 0.97488f
C54 drain_right.t0 a_n2524_n2088# 0.11627f
C55 drain_right.t9 a_n2524_n2088# 0.11627f
C56 drain_right.n34 a_n2524_n2088# 0.969695f
C57 drain_right.n35 a_n2524_n2088# 0.651568f
C58 drain_right.n36 a_n2524_n2088# 1.02878f
C59 drain_right.t8 a_n2524_n2088# 0.11627f
C60 drain_right.t5 a_n2524_n2088# 0.11627f
C61 drain_right.n37 a_n2524_n2088# 0.97488f
C62 drain_right.t3 a_n2524_n2088# 0.11627f
C63 drain_right.t10 a_n2524_n2088# 0.11627f
C64 drain_right.n38 a_n2524_n2088# 0.969699f
C65 drain_right.n39 a_n2524_n2088# 0.710645f
C66 drain_right.t4 a_n2524_n2088# 0.11627f
C67 drain_right.t2 a_n2524_n2088# 0.11627f
C68 drain_right.n40 a_n2524_n2088# 0.969699f
C69 drain_right.n41 a_n2524_n2088# 0.352975f
C70 drain_right.n42 a_n2524_n2088# 0.034468f
C71 drain_right.n43 a_n2524_n2088# 0.024522f
C72 drain_right.n44 a_n2524_n2088# 0.013177f
C73 drain_right.n45 a_n2524_n2088# 0.031146f
C74 drain_right.n46 a_n2524_n2088# 0.013952f
C75 drain_right.n47 a_n2524_n2088# 0.024522f
C76 drain_right.n48 a_n2524_n2088# 0.013177f
C77 drain_right.n49 a_n2524_n2088# 0.031146f
C78 drain_right.n50 a_n2524_n2088# 0.013952f
C79 drain_right.n51 a_n2524_n2088# 0.104939f
C80 drain_right.t7 a_n2524_n2088# 0.050765f
C81 drain_right.n52 a_n2524_n2088# 0.02336f
C82 drain_right.n53 a_n2524_n2088# 0.018398f
C83 drain_right.n54 a_n2524_n2088# 0.013177f
C84 drain_right.n55 a_n2524_n2088# 0.583488f
C85 drain_right.n56 a_n2524_n2088# 0.024522f
C86 drain_right.n57 a_n2524_n2088# 0.013177f
C87 drain_right.n58 a_n2524_n2088# 0.013952f
C88 drain_right.n59 a_n2524_n2088# 0.031146f
C89 drain_right.n60 a_n2524_n2088# 0.031146f
C90 drain_right.n61 a_n2524_n2088# 0.013952f
C91 drain_right.n62 a_n2524_n2088# 0.013177f
C92 drain_right.n63 a_n2524_n2088# 0.024522f
C93 drain_right.n64 a_n2524_n2088# 0.024522f
C94 drain_right.n65 a_n2524_n2088# 0.013177f
C95 drain_right.n66 a_n2524_n2088# 0.013952f
C96 drain_right.n67 a_n2524_n2088# 0.031146f
C97 drain_right.n68 a_n2524_n2088# 0.067426f
C98 drain_right.n69 a_n2524_n2088# 0.013952f
C99 drain_right.n70 a_n2524_n2088# 0.013177f
C100 drain_right.n71 a_n2524_n2088# 0.056682f
C101 drain_right.n72 a_n2524_n2088# 0.05466f
C102 drain_right.n73 a_n2524_n2088# 0.354704f
C103 minus.n0 a_n2524_n2088# 0.040087f
C104 minus.n1 a_n2524_n2088# 0.009097f
C105 minus.t9 a_n2524_n2088# 0.558115f
C106 minus.n2 a_n2524_n2088# 0.080174f
C107 minus.n3 a_n2524_n2088# 0.009097f
C108 minus.t3 a_n2524_n2088# 0.558115f
C109 minus.t8 a_n2524_n2088# 0.582249f
C110 minus.t5 a_n2524_n2088# 0.558115f
C111 minus.n4 a_n2524_n2088# 0.2592f
C112 minus.n5 a_n2524_n2088# 0.236095f
C113 minus.n6 a_n2524_n2088# 0.187211f
C114 minus.n7 a_n2524_n2088# 0.06677f
C115 minus.n8 a_n2524_n2088# 0.263825f
C116 minus.t10 a_n2524_n2088# 0.558115f
C117 minus.n9 a_n2524_n2088# 0.266544f
C118 minus.t11 a_n2524_n2088# 0.558115f
C119 minus.n10 a_n2524_n2088# 0.263825f
C120 minus.n11 a_n2524_n2088# 0.06677f
C121 minus.n12 a_n2524_n2088# 0.053491f
C122 minus.n13 a_n2524_n2088# 0.040087f
C123 minus.n14 a_n2524_n2088# 0.254234f
C124 minus.n15 a_n2524_n2088# 0.009097f
C125 minus.t6 a_n2524_n2088# 0.558115f
C126 minus.n16 a_n2524_n2088# 0.255223f
C127 minus.n17 a_n2524_n2088# 1.31237f
C128 minus.n18 a_n2524_n2088# 0.040087f
C129 minus.n19 a_n2524_n2088# 0.009097f
C130 minus.n20 a_n2524_n2088# 0.080174f
C131 minus.n21 a_n2524_n2088# 0.009097f
C132 minus.t7 a_n2524_n2088# 0.582249f
C133 minus.t0 a_n2524_n2088# 0.558115f
C134 minus.n22 a_n2524_n2088# 0.2592f
C135 minus.n23 a_n2524_n2088# 0.236095f
C136 minus.n24 a_n2524_n2088# 0.187211f
C137 minus.n25 a_n2524_n2088# 0.06677f
C138 minus.t2 a_n2524_n2088# 0.558115f
C139 minus.n26 a_n2524_n2088# 0.263825f
C140 minus.t13 a_n2524_n2088# 0.558115f
C141 minus.n27 a_n2524_n2088# 0.266544f
C142 minus.t4 a_n2524_n2088# 0.558115f
C143 minus.n28 a_n2524_n2088# 0.263825f
C144 minus.n29 a_n2524_n2088# 0.06677f
C145 minus.n30 a_n2524_n2088# 0.053491f
C146 minus.n31 a_n2524_n2088# 0.040087f
C147 minus.t12 a_n2524_n2088# 0.558115f
C148 minus.n32 a_n2524_n2088# 0.254234f
C149 minus.n33 a_n2524_n2088# 0.009097f
C150 minus.t1 a_n2524_n2088# 0.558115f
C151 minus.n34 a_n2524_n2088# 0.255223f
C152 minus.n35 a_n2524_n2088# 0.283188f
C153 minus.n36 a_n2524_n2088# 1.59459f
C154 source.n0 a_n2524_n2088# 0.039242f
C155 source.n1 a_n2524_n2088# 0.027919f
C156 source.n2 a_n2524_n2088# 0.015002f
C157 source.n3 a_n2524_n2088# 0.03546f
C158 source.n4 a_n2524_n2088# 0.015885f
C159 source.n5 a_n2524_n2088# 0.027919f
C160 source.n6 a_n2524_n2088# 0.015002f
C161 source.n7 a_n2524_n2088# 0.03546f
C162 source.n8 a_n2524_n2088# 0.015885f
C163 source.n9 a_n2524_n2088# 0.119473f
C164 source.t18 a_n2524_n2088# 0.057795f
C165 source.n10 a_n2524_n2088# 0.026595f
C166 source.n11 a_n2524_n2088# 0.020946f
C167 source.n12 a_n2524_n2088# 0.015002f
C168 source.n13 a_n2524_n2088# 0.664299f
C169 source.n14 a_n2524_n2088# 0.027919f
C170 source.n15 a_n2524_n2088# 0.015002f
C171 source.n16 a_n2524_n2088# 0.015885f
C172 source.n17 a_n2524_n2088# 0.03546f
C173 source.n18 a_n2524_n2088# 0.03546f
C174 source.n19 a_n2524_n2088# 0.015885f
C175 source.n20 a_n2524_n2088# 0.015002f
C176 source.n21 a_n2524_n2088# 0.027919f
C177 source.n22 a_n2524_n2088# 0.027919f
C178 source.n23 a_n2524_n2088# 0.015002f
C179 source.n24 a_n2524_n2088# 0.015885f
C180 source.n25 a_n2524_n2088# 0.03546f
C181 source.n26 a_n2524_n2088# 0.076765f
C182 source.n27 a_n2524_n2088# 0.015885f
C183 source.n28 a_n2524_n2088# 0.015002f
C184 source.n29 a_n2524_n2088# 0.064533f
C185 source.n30 a_n2524_n2088# 0.042953f
C186 source.n31 a_n2524_n2088# 0.74258f
C187 source.t14 a_n2524_n2088# 0.132373f
C188 source.t17 a_n2524_n2088# 0.132373f
C189 source.n32 a_n2524_n2088# 1.03093f
C190 source.n33 a_n2524_n2088# 0.436979f
C191 source.t15 a_n2524_n2088# 0.132373f
C192 source.t16 a_n2524_n2088# 0.132373f
C193 source.n34 a_n2524_n2088# 1.03093f
C194 source.n35 a_n2524_n2088# 0.436979f
C195 source.t12 a_n2524_n2088# 0.132373f
C196 source.t13 a_n2524_n2088# 0.132373f
C197 source.n36 a_n2524_n2088# 1.03093f
C198 source.n37 a_n2524_n2088# 0.435428f
C199 source.n38 a_n2524_n2088# 0.039242f
C200 source.n39 a_n2524_n2088# 0.027919f
C201 source.n40 a_n2524_n2088# 0.015002f
C202 source.n41 a_n2524_n2088# 0.03546f
C203 source.n42 a_n2524_n2088# 0.015885f
C204 source.n43 a_n2524_n2088# 0.027919f
C205 source.n44 a_n2524_n2088# 0.015002f
C206 source.n45 a_n2524_n2088# 0.03546f
C207 source.n46 a_n2524_n2088# 0.015885f
C208 source.n47 a_n2524_n2088# 0.119473f
C209 source.t0 a_n2524_n2088# 0.057795f
C210 source.n48 a_n2524_n2088# 0.026595f
C211 source.n49 a_n2524_n2088# 0.020946f
C212 source.n50 a_n2524_n2088# 0.015002f
C213 source.n51 a_n2524_n2088# 0.664299f
C214 source.n52 a_n2524_n2088# 0.027919f
C215 source.n53 a_n2524_n2088# 0.015002f
C216 source.n54 a_n2524_n2088# 0.015885f
C217 source.n55 a_n2524_n2088# 0.03546f
C218 source.n56 a_n2524_n2088# 0.03546f
C219 source.n57 a_n2524_n2088# 0.015885f
C220 source.n58 a_n2524_n2088# 0.015002f
C221 source.n59 a_n2524_n2088# 0.027919f
C222 source.n60 a_n2524_n2088# 0.027919f
C223 source.n61 a_n2524_n2088# 0.015002f
C224 source.n62 a_n2524_n2088# 0.015885f
C225 source.n63 a_n2524_n2088# 0.03546f
C226 source.n64 a_n2524_n2088# 0.076765f
C227 source.n65 a_n2524_n2088# 0.015885f
C228 source.n66 a_n2524_n2088# 0.015002f
C229 source.n67 a_n2524_n2088# 0.064533f
C230 source.n68 a_n2524_n2088# 0.042953f
C231 source.n69 a_n2524_n2088# 0.197561f
C232 source.t10 a_n2524_n2088# 0.132373f
C233 source.t2 a_n2524_n2088# 0.132373f
C234 source.n70 a_n2524_n2088# 1.03093f
C235 source.n71 a_n2524_n2088# 0.436979f
C236 source.t26 a_n2524_n2088# 0.132373f
C237 source.t25 a_n2524_n2088# 0.132373f
C238 source.n72 a_n2524_n2088# 1.03093f
C239 source.n73 a_n2524_n2088# 0.436979f
C240 source.t6 a_n2524_n2088# 0.132373f
C241 source.t3 a_n2524_n2088# 0.132373f
C242 source.n74 a_n2524_n2088# 1.03093f
C243 source.n75 a_n2524_n2088# 1.43872f
C244 source.t23 a_n2524_n2088# 0.132373f
C245 source.t19 a_n2524_n2088# 0.132373f
C246 source.n76 a_n2524_n2088# 1.03093f
C247 source.n77 a_n2524_n2088# 1.43873f
C248 source.t21 a_n2524_n2088# 0.132373f
C249 source.t11 a_n2524_n2088# 0.132373f
C250 source.n78 a_n2524_n2088# 1.03093f
C251 source.n79 a_n2524_n2088# 0.436986f
C252 source.t22 a_n2524_n2088# 0.132373f
C253 source.t24 a_n2524_n2088# 0.132373f
C254 source.n80 a_n2524_n2088# 1.03093f
C255 source.n81 a_n2524_n2088# 0.436986f
C256 source.n82 a_n2524_n2088# 0.039242f
C257 source.n83 a_n2524_n2088# 0.027919f
C258 source.n84 a_n2524_n2088# 0.015002f
C259 source.n85 a_n2524_n2088# 0.03546f
C260 source.n86 a_n2524_n2088# 0.015885f
C261 source.n87 a_n2524_n2088# 0.027919f
C262 source.n88 a_n2524_n2088# 0.015002f
C263 source.n89 a_n2524_n2088# 0.03546f
C264 source.n90 a_n2524_n2088# 0.015885f
C265 source.n91 a_n2524_n2088# 0.119473f
C266 source.t20 a_n2524_n2088# 0.057795f
C267 source.n92 a_n2524_n2088# 0.026595f
C268 source.n93 a_n2524_n2088# 0.020946f
C269 source.n94 a_n2524_n2088# 0.015002f
C270 source.n95 a_n2524_n2088# 0.664299f
C271 source.n96 a_n2524_n2088# 0.027919f
C272 source.n97 a_n2524_n2088# 0.015002f
C273 source.n98 a_n2524_n2088# 0.015885f
C274 source.n99 a_n2524_n2088# 0.03546f
C275 source.n100 a_n2524_n2088# 0.03546f
C276 source.n101 a_n2524_n2088# 0.015885f
C277 source.n102 a_n2524_n2088# 0.015002f
C278 source.n103 a_n2524_n2088# 0.027919f
C279 source.n104 a_n2524_n2088# 0.027919f
C280 source.n105 a_n2524_n2088# 0.015002f
C281 source.n106 a_n2524_n2088# 0.015885f
C282 source.n107 a_n2524_n2088# 0.03546f
C283 source.n108 a_n2524_n2088# 0.076765f
C284 source.n109 a_n2524_n2088# 0.015885f
C285 source.n110 a_n2524_n2088# 0.015002f
C286 source.n111 a_n2524_n2088# 0.064533f
C287 source.n112 a_n2524_n2088# 0.042953f
C288 source.n113 a_n2524_n2088# 0.197561f
C289 source.t7 a_n2524_n2088# 0.132373f
C290 source.t5 a_n2524_n2088# 0.132373f
C291 source.n114 a_n2524_n2088# 1.03093f
C292 source.n115 a_n2524_n2088# 0.435435f
C293 source.t8 a_n2524_n2088# 0.132373f
C294 source.t4 a_n2524_n2088# 0.132373f
C295 source.n116 a_n2524_n2088# 1.03093f
C296 source.n117 a_n2524_n2088# 0.436986f
C297 source.t9 a_n2524_n2088# 0.132373f
C298 source.t27 a_n2524_n2088# 0.132373f
C299 source.n118 a_n2524_n2088# 1.03093f
C300 source.n119 a_n2524_n2088# 0.436986f
C301 source.n120 a_n2524_n2088# 0.039242f
C302 source.n121 a_n2524_n2088# 0.027919f
C303 source.n122 a_n2524_n2088# 0.015002f
C304 source.n123 a_n2524_n2088# 0.03546f
C305 source.n124 a_n2524_n2088# 0.015885f
C306 source.n125 a_n2524_n2088# 0.027919f
C307 source.n126 a_n2524_n2088# 0.015002f
C308 source.n127 a_n2524_n2088# 0.03546f
C309 source.n128 a_n2524_n2088# 0.015885f
C310 source.n129 a_n2524_n2088# 0.119473f
C311 source.t1 a_n2524_n2088# 0.057795f
C312 source.n130 a_n2524_n2088# 0.026595f
C313 source.n131 a_n2524_n2088# 0.020946f
C314 source.n132 a_n2524_n2088# 0.015002f
C315 source.n133 a_n2524_n2088# 0.664299f
C316 source.n134 a_n2524_n2088# 0.027919f
C317 source.n135 a_n2524_n2088# 0.015002f
C318 source.n136 a_n2524_n2088# 0.015885f
C319 source.n137 a_n2524_n2088# 0.03546f
C320 source.n138 a_n2524_n2088# 0.03546f
C321 source.n139 a_n2524_n2088# 0.015885f
C322 source.n140 a_n2524_n2088# 0.015002f
C323 source.n141 a_n2524_n2088# 0.027919f
C324 source.n142 a_n2524_n2088# 0.027919f
C325 source.n143 a_n2524_n2088# 0.015002f
C326 source.n144 a_n2524_n2088# 0.015885f
C327 source.n145 a_n2524_n2088# 0.03546f
C328 source.n146 a_n2524_n2088# 0.076765f
C329 source.n147 a_n2524_n2088# 0.015885f
C330 source.n148 a_n2524_n2088# 0.015002f
C331 source.n149 a_n2524_n2088# 0.064533f
C332 source.n150 a_n2524_n2088# 0.042953f
C333 source.n151 a_n2524_n2088# 0.341903f
C334 source.n152 a_n2524_n2088# 1.16182f
C335 drain_left.n0 a_n2524_n2088# 0.034917f
C336 drain_left.n1 a_n2524_n2088# 0.024841f
C337 drain_left.n2 a_n2524_n2088# 0.013349f
C338 drain_left.n3 a_n2524_n2088# 0.031551f
C339 drain_left.n4 a_n2524_n2088# 0.014134f
C340 drain_left.n5 a_n2524_n2088# 0.024841f
C341 drain_left.n6 a_n2524_n2088# 0.013349f
C342 drain_left.n7 a_n2524_n2088# 0.031551f
C343 drain_left.n8 a_n2524_n2088# 0.014134f
C344 drain_left.n9 a_n2524_n2088# 0.106303f
C345 drain_left.t12 a_n2524_n2088# 0.051424f
C346 drain_left.n10 a_n2524_n2088# 0.023664f
C347 drain_left.n11 a_n2524_n2088# 0.018637f
C348 drain_left.n12 a_n2524_n2088# 0.013349f
C349 drain_left.n13 a_n2524_n2088# 0.591074f
C350 drain_left.n14 a_n2524_n2088# 0.024841f
C351 drain_left.n15 a_n2524_n2088# 0.013349f
C352 drain_left.n16 a_n2524_n2088# 0.014134f
C353 drain_left.n17 a_n2524_n2088# 0.031551f
C354 drain_left.n18 a_n2524_n2088# 0.031551f
C355 drain_left.n19 a_n2524_n2088# 0.014134f
C356 drain_left.n20 a_n2524_n2088# 0.013349f
C357 drain_left.n21 a_n2524_n2088# 0.024841f
C358 drain_left.n22 a_n2524_n2088# 0.024841f
C359 drain_left.n23 a_n2524_n2088# 0.013349f
C360 drain_left.n24 a_n2524_n2088# 0.014134f
C361 drain_left.n25 a_n2524_n2088# 0.031551f
C362 drain_left.n26 a_n2524_n2088# 0.068303f
C363 drain_left.n27 a_n2524_n2088# 0.014134f
C364 drain_left.n28 a_n2524_n2088# 0.013349f
C365 drain_left.n29 a_n2524_n2088# 0.057419f
C366 drain_left.n30 a_n2524_n2088# 0.05783f
C367 drain_left.t8 a_n2524_n2088# 0.117782f
C368 drain_left.t13 a_n2524_n2088# 0.117782f
C369 drain_left.n31 a_n2524_n2088# 0.982302f
C370 drain_left.n32 a_n2524_n2088# 0.457846f
C371 drain_left.t0 a_n2524_n2088# 0.117782f
C372 drain_left.t7 a_n2524_n2088# 0.117782f
C373 drain_left.n33 a_n2524_n2088# 0.987555f
C374 drain_left.t5 a_n2524_n2088# 0.117782f
C375 drain_left.t3 a_n2524_n2088# 0.117782f
C376 drain_left.n34 a_n2524_n2088# 0.982302f
C377 drain_left.n35 a_n2524_n2088# 0.660039f
C378 drain_left.n36 a_n2524_n2088# 1.09206f
C379 drain_left.n37 a_n2524_n2088# 0.034917f
C380 drain_left.n38 a_n2524_n2088# 0.024841f
C381 drain_left.n39 a_n2524_n2088# 0.013349f
C382 drain_left.n40 a_n2524_n2088# 0.031551f
C383 drain_left.n41 a_n2524_n2088# 0.014134f
C384 drain_left.n42 a_n2524_n2088# 0.024841f
C385 drain_left.n43 a_n2524_n2088# 0.013349f
C386 drain_left.n44 a_n2524_n2088# 0.031551f
C387 drain_left.n45 a_n2524_n2088# 0.014134f
C388 drain_left.n46 a_n2524_n2088# 0.106303f
C389 drain_left.t11 a_n2524_n2088# 0.051424f
C390 drain_left.n47 a_n2524_n2088# 0.023664f
C391 drain_left.n48 a_n2524_n2088# 0.018637f
C392 drain_left.n49 a_n2524_n2088# 0.013349f
C393 drain_left.n50 a_n2524_n2088# 0.591074f
C394 drain_left.n51 a_n2524_n2088# 0.024841f
C395 drain_left.n52 a_n2524_n2088# 0.013349f
C396 drain_left.n53 a_n2524_n2088# 0.014134f
C397 drain_left.n54 a_n2524_n2088# 0.031551f
C398 drain_left.n55 a_n2524_n2088# 0.031551f
C399 drain_left.n56 a_n2524_n2088# 0.014134f
C400 drain_left.n57 a_n2524_n2088# 0.013349f
C401 drain_left.n58 a_n2524_n2088# 0.024841f
C402 drain_left.n59 a_n2524_n2088# 0.024841f
C403 drain_left.n60 a_n2524_n2088# 0.013349f
C404 drain_left.n61 a_n2524_n2088# 0.014134f
C405 drain_left.n62 a_n2524_n2088# 0.031551f
C406 drain_left.n63 a_n2524_n2088# 0.068303f
C407 drain_left.n64 a_n2524_n2088# 0.014134f
C408 drain_left.n65 a_n2524_n2088# 0.013349f
C409 drain_left.n66 a_n2524_n2088# 0.057419f
C410 drain_left.n67 a_n2524_n2088# 0.05783f
C411 drain_left.t6 a_n2524_n2088# 0.117782f
C412 drain_left.t4 a_n2524_n2088# 0.117782f
C413 drain_left.n68 a_n2524_n2088# 0.982307f
C414 drain_left.n69 a_n2524_n2088# 0.480913f
C415 drain_left.t1 a_n2524_n2088# 0.117782f
C416 drain_left.t2 a_n2524_n2088# 0.117782f
C417 drain_left.n70 a_n2524_n2088# 0.982307f
C418 drain_left.n71 a_n2524_n2088# 0.357564f
C419 drain_left.t10 a_n2524_n2088# 0.117782f
C420 drain_left.t9 a_n2524_n2088# 0.117782f
C421 drain_left.n72 a_n2524_n2088# 0.982302f
C422 drain_left.n73 a_n2524_n2088# 0.580319f
C423 plus.n0 a_n2524_n2088# 0.041059f
C424 plus.t6 a_n2524_n2088# 0.571645f
C425 plus.t7 a_n2524_n2088# 0.571645f
C426 plus.n1 a_n2524_n2088# 0.041059f
C427 plus.t10 a_n2524_n2088# 0.571645f
C428 plus.n2 a_n2524_n2088# 0.270221f
C429 plus.n3 a_n2524_n2088# 0.068388f
C430 plus.t8 a_n2524_n2088# 0.571645f
C431 plus.t9 a_n2524_n2088# 0.571645f
C432 plus.t11 a_n2524_n2088# 0.571645f
C433 plus.n4 a_n2524_n2088# 0.265483f
C434 plus.t12 a_n2524_n2088# 0.596364f
C435 plus.n5 a_n2524_n2088# 0.241819f
C436 plus.n6 a_n2524_n2088# 0.191749f
C437 plus.n7 a_n2524_n2088# 0.009317f
C438 plus.n8 a_n2524_n2088# 0.270221f
C439 plus.n9 a_n2524_n2088# 0.273005f
C440 plus.n10 a_n2524_n2088# 0.082117f
C441 plus.n11 a_n2524_n2088# 0.068388f
C442 plus.n12 a_n2524_n2088# 0.054787f
C443 plus.n13 a_n2524_n2088# 0.009317f
C444 plus.n14 a_n2524_n2088# 0.260397f
C445 plus.n15 a_n2524_n2088# 0.009317f
C446 plus.n16 a_n2524_n2088# 0.26141f
C447 plus.n17 a_n2524_n2088# 0.374446f
C448 plus.n18 a_n2524_n2088# 0.041059f
C449 plus.t1 a_n2524_n2088# 0.571645f
C450 plus.n19 a_n2524_n2088# 0.041059f
C451 plus.t5 a_n2524_n2088# 0.571645f
C452 plus.t3 a_n2524_n2088# 0.571645f
C453 plus.n20 a_n2524_n2088# 0.270221f
C454 plus.n21 a_n2524_n2088# 0.068388f
C455 plus.t13 a_n2524_n2088# 0.571645f
C456 plus.t2 a_n2524_n2088# 0.571645f
C457 plus.t0 a_n2524_n2088# 0.571645f
C458 plus.n22 a_n2524_n2088# 0.265483f
C459 plus.t4 a_n2524_n2088# 0.596364f
C460 plus.n23 a_n2524_n2088# 0.241819f
C461 plus.n24 a_n2524_n2088# 0.191749f
C462 plus.n25 a_n2524_n2088# 0.009317f
C463 plus.n26 a_n2524_n2088# 0.270221f
C464 plus.n27 a_n2524_n2088# 0.273005f
C465 plus.n28 a_n2524_n2088# 0.082117f
C466 plus.n29 a_n2524_n2088# 0.068388f
C467 plus.n30 a_n2524_n2088# 0.054787f
C468 plus.n31 a_n2524_n2088# 0.009317f
C469 plus.n32 a_n2524_n2088# 0.260397f
C470 plus.n33 a_n2524_n2088# 0.009317f
C471 plus.n34 a_n2524_n2088# 0.26141f
C472 plus.n35 a_n2524_n2088# 1.21763f
.ends

