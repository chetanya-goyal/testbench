* NGSPICE file created from diffpair623.ext - technology: sky130A

.subckt diffpair623 minus drain_right drain_left source plus
X0 drain_left.t7 plus.t0 source.t15 a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X1 a_n1746_n4888# a_n1746_n4888# a_n1746_n4888# a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.7
X2 source.t7 minus.t0 drain_right.t7 a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X3 source.t11 plus.t1 drain_left.t6 a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X4 a_n1746_n4888# a_n1746_n4888# a_n1746_n4888# a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X5 drain_right.t6 minus.t1 source.t3 a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X6 source.t8 plus.t2 drain_left.t5 a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X7 source.t6 minus.t2 drain_right.t5 a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X8 source.t9 plus.t3 drain_left.t4 a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X9 drain_right.t4 minus.t3 source.t5 a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X10 source.t4 minus.t4 drain_right.t3 a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X11 a_n1746_n4888# a_n1746_n4888# a_n1746_n4888# a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X12 drain_right.t2 minus.t5 source.t0 a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X13 drain_left.t3 plus.t4 source.t10 a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X14 source.t12 plus.t5 drain_left.t2 a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X15 drain_right.t1 minus.t6 source.t2 a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X16 drain_left.t1 plus.t6 source.t14 a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X17 a_n1746_n4888# a_n1746_n4888# a_n1746_n4888# a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X18 drain_left.t0 plus.t7 source.t13 a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X19 source.t1 minus.t7 drain_right.t0 a_n1746_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
R0 plus.n3 plus.t3 766.869
R1 plus.n13 plus.t0 766.869
R2 plus.n8 plus.t4 744.691
R3 plus.n6 plus.t2 744.691
R4 plus.n2 plus.t6 744.691
R5 plus.n18 plus.t5 744.691
R6 plus.n16 plus.t7 744.691
R7 plus.n12 plus.t1 744.691
R8 plus.n5 plus.n4 161.3
R9 plus.n6 plus.n1 161.3
R10 plus.n7 plus.n0 161.3
R11 plus.n9 plus.n8 161.3
R12 plus.n15 plus.n14 161.3
R13 plus.n16 plus.n11 161.3
R14 plus.n17 plus.n10 161.3
R15 plus.n19 plus.n18 161.3
R16 plus.n4 plus.n3 44.862
R17 plus.n14 plus.n13 44.862
R18 plus plus.n19 32.7793
R19 plus.n8 plus.n7 28.4823
R20 plus.n18 plus.n17 28.4823
R21 plus.n5 plus.n2 24.1005
R22 plus.n6 plus.n5 24.1005
R23 plus.n16 plus.n15 24.1005
R24 plus.n15 plus.n12 24.1005
R25 plus.n7 plus.n6 19.7187
R26 plus.n17 plus.n16 19.7187
R27 plus.n3 plus.n2 19.7081
R28 plus.n13 plus.n12 19.7081
R29 plus plus.n9 15.3073
R30 plus.n4 plus.n1 0.189894
R31 plus.n1 plus.n0 0.189894
R32 plus.n9 plus.n0 0.189894
R33 plus.n19 plus.n10 0.189894
R34 plus.n11 plus.n10 0.189894
R35 plus.n14 plus.n11 0.189894
R36 source.n0 source.t10 44.1297
R37 source.n3 source.t9 44.1296
R38 source.n4 source.t2 44.1296
R39 source.n7 source.t1 44.1296
R40 source.n15 source.t3 44.1295
R41 source.n12 source.t4 44.1295
R42 source.n11 source.t15 44.1295
R43 source.n8 source.t12 44.1295
R44 source.n2 source.n1 43.1397
R45 source.n6 source.n5 43.1397
R46 source.n14 source.n13 43.1396
R47 source.n10 source.n9 43.1396
R48 source.n8 source.n7 28.2363
R49 source.n16 source.n0 22.5294
R50 source.n16 source.n15 5.7074
R51 source.n13 source.t5 0.9905
R52 source.n13 source.t7 0.9905
R53 source.n9 source.t13 0.9905
R54 source.n9 source.t11 0.9905
R55 source.n1 source.t14 0.9905
R56 source.n1 source.t8 0.9905
R57 source.n5 source.t0 0.9905
R58 source.n5 source.t6 0.9905
R59 source.n7 source.n6 0.888431
R60 source.n6 source.n4 0.888431
R61 source.n3 source.n2 0.888431
R62 source.n2 source.n0 0.888431
R63 source.n10 source.n8 0.888431
R64 source.n11 source.n10 0.888431
R65 source.n14 source.n12 0.888431
R66 source.n15 source.n14 0.888431
R67 source.n4 source.n3 0.470328
R68 source.n12 source.n11 0.470328
R69 source source.n16 0.188
R70 drain_left.n5 drain_left.n3 60.7064
R71 drain_left.n2 drain_left.n1 60.207
R72 drain_left.n2 drain_left.n0 60.207
R73 drain_left.n5 drain_left.n4 59.8185
R74 drain_left drain_left.n2 36.5354
R75 drain_left drain_left.n5 6.54115
R76 drain_left.n1 drain_left.t6 0.9905
R77 drain_left.n1 drain_left.t7 0.9905
R78 drain_left.n0 drain_left.t2 0.9905
R79 drain_left.n0 drain_left.t0 0.9905
R80 drain_left.n4 drain_left.t5 0.9905
R81 drain_left.n4 drain_left.t3 0.9905
R82 drain_left.n3 drain_left.t4 0.9905
R83 drain_left.n3 drain_left.t1 0.9905
R84 minus.n3 minus.t6 766.869
R85 minus.n13 minus.t4 766.869
R86 minus.n2 minus.t2 744.691
R87 minus.n6 minus.t5 744.691
R88 minus.n8 minus.t7 744.691
R89 minus.n12 minus.t3 744.691
R90 minus.n16 minus.t0 744.691
R91 minus.n18 minus.t1 744.691
R92 minus.n9 minus.n8 161.3
R93 minus.n7 minus.n0 161.3
R94 minus.n6 minus.n5 161.3
R95 minus.n4 minus.n1 161.3
R96 minus.n19 minus.n18 161.3
R97 minus.n17 minus.n10 161.3
R98 minus.n16 minus.n15 161.3
R99 minus.n14 minus.n11 161.3
R100 minus.n4 minus.n3 44.862
R101 minus.n14 minus.n13 44.862
R102 minus.n20 minus.n9 41.9285
R103 minus.n8 minus.n7 28.4823
R104 minus.n18 minus.n17 28.4823
R105 minus.n6 minus.n1 24.1005
R106 minus.n2 minus.n1 24.1005
R107 minus.n12 minus.n11 24.1005
R108 minus.n16 minus.n11 24.1005
R109 minus.n7 minus.n6 19.7187
R110 minus.n17 minus.n16 19.7187
R111 minus.n3 minus.n2 19.7081
R112 minus.n13 minus.n12 19.7081
R113 minus.n20 minus.n19 6.63308
R114 minus.n9 minus.n0 0.189894
R115 minus.n5 minus.n0 0.189894
R116 minus.n5 minus.n4 0.189894
R117 minus.n15 minus.n14 0.189894
R118 minus.n15 minus.n10 0.189894
R119 minus.n19 minus.n10 0.189894
R120 minus minus.n20 0.188
R121 drain_right.n5 drain_right.n3 60.7064
R122 drain_right.n2 drain_right.n1 60.207
R123 drain_right.n2 drain_right.n0 60.207
R124 drain_right.n5 drain_right.n4 59.8185
R125 drain_right drain_right.n2 35.9822
R126 drain_right drain_right.n5 6.54115
R127 drain_right.n1 drain_right.t7 0.9905
R128 drain_right.n1 drain_right.t6 0.9905
R129 drain_right.n0 drain_right.t3 0.9905
R130 drain_right.n0 drain_right.t4 0.9905
R131 drain_right.n3 drain_right.t5 0.9905
R132 drain_right.n3 drain_right.t1 0.9905
R133 drain_right.n4 drain_right.t0 0.9905
R134 drain_right.n4 drain_right.t2 0.9905
C0 source minus 8.386049f
C1 drain_left source 17.2665f
C2 drain_right source 17.268301f
C3 drain_left minus 0.171089f
C4 source plus 8.40008f
C5 drain_right minus 8.962191f
C6 drain_left drain_right 0.821811f
C7 plus minus 6.80089f
C8 drain_left plus 9.13103f
C9 drain_right plus 0.322995f
C10 drain_right a_n1746_n4888# 7.1781f
C11 drain_left a_n1746_n4888# 7.42522f
C12 source a_n1746_n4888# 13.486982f
C13 minus a_n1746_n4888# 7.302223f
C14 plus a_n1746_n4888# 9.41912f
C15 drain_right.t3 a_n1746_n4888# 0.432364f
C16 drain_right.t4 a_n1746_n4888# 0.432364f
C17 drain_right.n0 a_n1746_n4888# 3.95506f
C18 drain_right.t7 a_n1746_n4888# 0.432364f
C19 drain_right.t6 a_n1746_n4888# 0.432364f
C20 drain_right.n1 a_n1746_n4888# 3.95506f
C21 drain_right.n2 a_n1746_n4888# 2.52482f
C22 drain_right.t5 a_n1746_n4888# 0.432364f
C23 drain_right.t1 a_n1746_n4888# 0.432364f
C24 drain_right.n3 a_n1746_n4888# 3.95859f
C25 drain_right.t0 a_n1746_n4888# 0.432364f
C26 drain_right.t2 a_n1746_n4888# 0.432364f
C27 drain_right.n4 a_n1746_n4888# 3.95276f
C28 drain_right.n5 a_n1746_n4888# 1.02196f
C29 minus.n0 a_n1746_n4888# 0.043724f
C30 minus.n1 a_n1746_n4888# 0.009922f
C31 minus.t5 a_n1746_n4888# 1.73351f
C32 minus.t6 a_n1746_n4888# 1.75219f
C33 minus.t2 a_n1746_n4888# 1.73351f
C34 minus.n2 a_n1746_n4888# 0.650375f
C35 minus.n3 a_n1746_n4888# 0.631754f
C36 minus.n4 a_n1746_n4888# 0.181825f
C37 minus.n5 a_n1746_n4888# 0.043724f
C38 minus.n6 a_n1746_n4888# 0.646419f
C39 minus.n7 a_n1746_n4888# 0.009922f
C40 minus.t7 a_n1746_n4888# 1.73351f
C41 minus.n8 a_n1746_n4888# 0.643588f
C42 minus.n9 a_n1746_n4888# 1.9354f
C43 minus.n10 a_n1746_n4888# 0.043724f
C44 minus.n11 a_n1746_n4888# 0.009922f
C45 minus.t4 a_n1746_n4888# 1.75219f
C46 minus.t3 a_n1746_n4888# 1.73351f
C47 minus.n12 a_n1746_n4888# 0.650375f
C48 minus.n13 a_n1746_n4888# 0.631754f
C49 minus.n14 a_n1746_n4888# 0.181825f
C50 minus.n15 a_n1746_n4888# 0.043724f
C51 minus.t0 a_n1746_n4888# 1.73351f
C52 minus.n16 a_n1746_n4888# 0.646419f
C53 minus.n17 a_n1746_n4888# 0.009922f
C54 minus.t1 a_n1746_n4888# 1.73351f
C55 minus.n18 a_n1746_n4888# 0.643588f
C56 minus.n19 a_n1746_n4888# 0.299479f
C57 minus.n20 a_n1746_n4888# 2.30848f
C58 drain_left.t2 a_n1746_n4888# 0.432249f
C59 drain_left.t0 a_n1746_n4888# 0.432249f
C60 drain_left.n0 a_n1746_n4888# 3.95401f
C61 drain_left.t6 a_n1746_n4888# 0.432249f
C62 drain_left.t7 a_n1746_n4888# 0.432249f
C63 drain_left.n1 a_n1746_n4888# 3.95401f
C64 drain_left.n2 a_n1746_n4888# 2.58118f
C65 drain_left.t4 a_n1746_n4888# 0.432249f
C66 drain_left.t1 a_n1746_n4888# 0.432249f
C67 drain_left.n3 a_n1746_n4888# 3.95754f
C68 drain_left.t5 a_n1746_n4888# 0.432249f
C69 drain_left.t3 a_n1746_n4888# 0.432249f
C70 drain_left.n4 a_n1746_n4888# 3.95171f
C71 drain_left.n5 a_n1746_n4888# 1.02169f
C72 source.t10 a_n1746_n4888# 3.4853f
C73 source.n0 a_n1746_n4888# 1.5162f
C74 source.t14 a_n1746_n4888# 0.304969f
C75 source.t8 a_n1746_n4888# 0.304969f
C76 source.n1 a_n1746_n4888# 2.72655f
C77 source.n2 a_n1746_n4888# 0.308562f
C78 source.t9 a_n1746_n4888# 3.4853f
C79 source.n3 a_n1746_n4888# 0.355544f
C80 source.t2 a_n1746_n4888# 3.4853f
C81 source.n4 a_n1746_n4888# 0.355544f
C82 source.t0 a_n1746_n4888# 0.304969f
C83 source.t6 a_n1746_n4888# 0.304969f
C84 source.n5 a_n1746_n4888# 2.72655f
C85 source.n6 a_n1746_n4888# 0.308562f
C86 source.t1 a_n1746_n4888# 3.4853f
C87 source.n7 a_n1746_n4888# 1.86725f
C88 source.t12 a_n1746_n4888# 3.48529f
C89 source.n8 a_n1746_n4888# 1.86726f
C90 source.t13 a_n1746_n4888# 0.304969f
C91 source.t11 a_n1746_n4888# 0.304969f
C92 source.n9 a_n1746_n4888# 2.72655f
C93 source.n10 a_n1746_n4888# 0.308557f
C94 source.t15 a_n1746_n4888# 3.48529f
C95 source.n11 a_n1746_n4888# 0.355563f
C96 source.t4 a_n1746_n4888# 3.48529f
C97 source.n12 a_n1746_n4888# 0.355563f
C98 source.t5 a_n1746_n4888# 0.304969f
C99 source.t7 a_n1746_n4888# 0.304969f
C100 source.n13 a_n1746_n4888# 2.72655f
C101 source.n14 a_n1746_n4888# 0.308557f
C102 source.t3 a_n1746_n4888# 3.48529f
C103 source.n15 a_n1746_n4888# 0.481433f
C104 source.n16 a_n1746_n4888# 1.75061f
C105 plus.n0 a_n1746_n4888# 0.044066f
C106 plus.t4 a_n1746_n4888# 1.74705f
C107 plus.t2 a_n1746_n4888# 1.74705f
C108 plus.n1 a_n1746_n4888# 0.044066f
C109 plus.t6 a_n1746_n4888# 1.74705f
C110 plus.n2 a_n1746_n4888# 0.655458f
C111 plus.t3 a_n1746_n4888# 1.76589f
C112 plus.n3 a_n1746_n4888# 0.636691f
C113 plus.n4 a_n1746_n4888# 0.183246f
C114 plus.n5 a_n1746_n4888# 0.009999f
C115 plus.n6 a_n1746_n4888# 0.65147f
C116 plus.n7 a_n1746_n4888# 0.009999f
C117 plus.n8 a_n1746_n4888# 0.648618f
C118 plus.n9 a_n1746_n4888# 0.682563f
C119 plus.n10 a_n1746_n4888# 0.044066f
C120 plus.t5 a_n1746_n4888# 1.74705f
C121 plus.n11 a_n1746_n4888# 0.044066f
C122 plus.t7 a_n1746_n4888# 1.74705f
C123 plus.t1 a_n1746_n4888# 1.74705f
C124 plus.n12 a_n1746_n4888# 0.655458f
C125 plus.t0 a_n1746_n4888# 1.76589f
C126 plus.n13 a_n1746_n4888# 0.636691f
C127 plus.n14 a_n1746_n4888# 0.183246f
C128 plus.n15 a_n1746_n4888# 0.009999f
C129 plus.n16 a_n1746_n4888# 0.65147f
C130 plus.n17 a_n1746_n4888# 0.009999f
C131 plus.n18 a_n1746_n4888# 0.648618f
C132 plus.n19 a_n1746_n4888# 1.54323f
.ends

