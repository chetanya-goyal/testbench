* NGSPICE file created from diffpair275.ext - technology: sky130A

.subckt diffpair275 minus drain_right drain_left source plus
X0 source.t23 minus.t0 drain_right.t10 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X1 source.t22 minus.t1 drain_right.t1 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X2 drain_right.t6 minus.t2 source.t21 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X3 source.t9 plus.t0 drain_left.t11 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X4 a_n1598_n2088# a_n1598_n2088# a_n1598_n2088# a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.3
X5 source.t0 plus.t1 drain_left.t10 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X6 source.t8 plus.t2 drain_left.t9 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X7 source.t11 plus.t3 drain_left.t8 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X8 drain_right.t11 minus.t3 source.t20 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X9 drain_right.t8 minus.t4 source.t19 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X10 a_n1598_n2088# a_n1598_n2088# a_n1598_n2088# a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X11 drain_right.t2 minus.t5 source.t18 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X12 source.t1 plus.t4 drain_left.t7 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X13 drain_left.t6 plus.t5 source.t2 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X14 drain_left.t5 plus.t6 source.t3 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X15 drain_left.t4 plus.t7 source.t7 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X16 source.t17 minus.t6 drain_right.t7 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X17 drain_right.t4 minus.t7 source.t16 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X18 drain_left.t3 plus.t8 source.t10 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.3
X19 source.t15 minus.t8 drain_right.t0 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X20 source.t14 minus.t9 drain_right.t9 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.3
X21 source.t4 plus.t9 drain_left.t2 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X22 drain_right.t5 minus.t10 source.t13 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X23 drain_left.t1 plus.t10 source.t6 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X24 source.t12 minus.t11 drain_right.t3 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
X25 a_n1598_n2088# a_n1598_n2088# a_n1598_n2088# a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X26 a_n1598_n2088# a_n1598_n2088# a_n1598_n2088# a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.3
X27 drain_left.t0 plus.t11 source.t5 a_n1598_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.3
R0 minus.n13 minus.t1 633.904
R1 minus.n2 minus.t7 633.904
R2 minus.n28 minus.t5 633.904
R3 minus.n17 minus.t9 633.904
R4 minus.n12 minus.t10 586.433
R5 minus.n10 minus.t6 586.433
R6 minus.n3 minus.t2 586.433
R7 minus.n4 minus.t11 586.433
R8 minus.n27 minus.t0 586.433
R9 minus.n25 minus.t3 586.433
R10 minus.n19 minus.t8 586.433
R11 minus.n18 minus.t4 586.433
R12 minus.n6 minus.n2 161.489
R13 minus.n21 minus.n17 161.489
R14 minus.n14 minus.n13 161.3
R15 minus.n11 minus.n0 161.3
R16 minus.n9 minus.n8 161.3
R17 minus.n7 minus.n1 161.3
R18 minus.n6 minus.n5 161.3
R19 minus.n29 minus.n28 161.3
R20 minus.n26 minus.n15 161.3
R21 minus.n24 minus.n23 161.3
R22 minus.n22 minus.n16 161.3
R23 minus.n21 minus.n20 161.3
R24 minus.n9 minus.n1 73.0308
R25 minus.n24 minus.n16 73.0308
R26 minus.n11 minus.n10 63.5369
R27 minus.n5 minus.n3 63.5369
R28 minus.n20 minus.n19 63.5369
R29 minus.n26 minus.n25 63.5369
R30 minus.n13 minus.n12 44.549
R31 minus.n4 minus.n2 44.549
R32 minus.n18 minus.n17 44.549
R33 minus.n28 minus.n27 44.549
R34 minus.n30 minus.n14 30.6407
R35 minus.n12 minus.n11 28.4823
R36 minus.n5 minus.n4 28.4823
R37 minus.n20 minus.n18 28.4823
R38 minus.n27 minus.n26 28.4823
R39 minus.n10 minus.n9 9.49444
R40 minus.n3 minus.n1 9.49444
R41 minus.n19 minus.n16 9.49444
R42 minus.n25 minus.n24 9.49444
R43 minus.n30 minus.n29 6.51186
R44 minus.n14 minus.n0 0.189894
R45 minus.n8 minus.n0 0.189894
R46 minus.n8 minus.n7 0.189894
R47 minus.n7 minus.n6 0.189894
R48 minus.n22 minus.n21 0.189894
R49 minus.n23 minus.n22 0.189894
R50 minus.n23 minus.n15 0.189894
R51 minus.n29 minus.n15 0.189894
R52 minus minus.n30 0.188
R53 drain_right.n6 drain_right.n4 67.7338
R54 drain_right.n3 drain_right.n2 67.6784
R55 drain_right.n3 drain_right.n0 67.6784
R56 drain_right.n6 drain_right.n5 67.1908
R57 drain_right.n8 drain_right.n7 67.1908
R58 drain_right.n3 drain_right.n1 67.1907
R59 drain_right drain_right.n3 24.9839
R60 drain_right drain_right.n8 6.19632
R61 drain_right.n1 drain_right.t0 3.3005
R62 drain_right.n1 drain_right.t11 3.3005
R63 drain_right.n2 drain_right.t10 3.3005
R64 drain_right.n2 drain_right.t2 3.3005
R65 drain_right.n0 drain_right.t9 3.3005
R66 drain_right.n0 drain_right.t8 3.3005
R67 drain_right.n4 drain_right.t3 3.3005
R68 drain_right.n4 drain_right.t4 3.3005
R69 drain_right.n5 drain_right.t7 3.3005
R70 drain_right.n5 drain_right.t6 3.3005
R71 drain_right.n7 drain_right.t1 3.3005
R72 drain_right.n7 drain_right.t5 3.3005
R73 drain_right.n8 drain_right.n6 0.543603
R74 source.n266 source.n240 289.615
R75 source.n230 source.n204 289.615
R76 source.n198 source.n172 289.615
R77 source.n162 source.n136 289.615
R78 source.n26 source.n0 289.615
R79 source.n62 source.n36 289.615
R80 source.n94 source.n68 289.615
R81 source.n130 source.n104 289.615
R82 source.n251 source.n250 185
R83 source.n248 source.n247 185
R84 source.n257 source.n256 185
R85 source.n259 source.n258 185
R86 source.n244 source.n243 185
R87 source.n265 source.n264 185
R88 source.n267 source.n266 185
R89 source.n215 source.n214 185
R90 source.n212 source.n211 185
R91 source.n221 source.n220 185
R92 source.n223 source.n222 185
R93 source.n208 source.n207 185
R94 source.n229 source.n228 185
R95 source.n231 source.n230 185
R96 source.n183 source.n182 185
R97 source.n180 source.n179 185
R98 source.n189 source.n188 185
R99 source.n191 source.n190 185
R100 source.n176 source.n175 185
R101 source.n197 source.n196 185
R102 source.n199 source.n198 185
R103 source.n147 source.n146 185
R104 source.n144 source.n143 185
R105 source.n153 source.n152 185
R106 source.n155 source.n154 185
R107 source.n140 source.n139 185
R108 source.n161 source.n160 185
R109 source.n163 source.n162 185
R110 source.n27 source.n26 185
R111 source.n25 source.n24 185
R112 source.n4 source.n3 185
R113 source.n19 source.n18 185
R114 source.n17 source.n16 185
R115 source.n8 source.n7 185
R116 source.n11 source.n10 185
R117 source.n63 source.n62 185
R118 source.n61 source.n60 185
R119 source.n40 source.n39 185
R120 source.n55 source.n54 185
R121 source.n53 source.n52 185
R122 source.n44 source.n43 185
R123 source.n47 source.n46 185
R124 source.n95 source.n94 185
R125 source.n93 source.n92 185
R126 source.n72 source.n71 185
R127 source.n87 source.n86 185
R128 source.n85 source.n84 185
R129 source.n76 source.n75 185
R130 source.n79 source.n78 185
R131 source.n131 source.n130 185
R132 source.n129 source.n128 185
R133 source.n108 source.n107 185
R134 source.n123 source.n122 185
R135 source.n121 source.n120 185
R136 source.n112 source.n111 185
R137 source.n115 source.n114 185
R138 source.t18 source.n249 147.661
R139 source.t14 source.n213 147.661
R140 source.t3 source.n181 147.661
R141 source.t11 source.n145 147.661
R142 source.t10 source.n9 147.661
R143 source.t0 source.n45 147.661
R144 source.t16 source.n77 147.661
R145 source.t22 source.n113 147.661
R146 source.n250 source.n247 104.615
R147 source.n257 source.n247 104.615
R148 source.n258 source.n257 104.615
R149 source.n258 source.n243 104.615
R150 source.n265 source.n243 104.615
R151 source.n266 source.n265 104.615
R152 source.n214 source.n211 104.615
R153 source.n221 source.n211 104.615
R154 source.n222 source.n221 104.615
R155 source.n222 source.n207 104.615
R156 source.n229 source.n207 104.615
R157 source.n230 source.n229 104.615
R158 source.n182 source.n179 104.615
R159 source.n189 source.n179 104.615
R160 source.n190 source.n189 104.615
R161 source.n190 source.n175 104.615
R162 source.n197 source.n175 104.615
R163 source.n198 source.n197 104.615
R164 source.n146 source.n143 104.615
R165 source.n153 source.n143 104.615
R166 source.n154 source.n153 104.615
R167 source.n154 source.n139 104.615
R168 source.n161 source.n139 104.615
R169 source.n162 source.n161 104.615
R170 source.n26 source.n25 104.615
R171 source.n25 source.n3 104.615
R172 source.n18 source.n3 104.615
R173 source.n18 source.n17 104.615
R174 source.n17 source.n7 104.615
R175 source.n10 source.n7 104.615
R176 source.n62 source.n61 104.615
R177 source.n61 source.n39 104.615
R178 source.n54 source.n39 104.615
R179 source.n54 source.n53 104.615
R180 source.n53 source.n43 104.615
R181 source.n46 source.n43 104.615
R182 source.n94 source.n93 104.615
R183 source.n93 source.n71 104.615
R184 source.n86 source.n71 104.615
R185 source.n86 source.n85 104.615
R186 source.n85 source.n75 104.615
R187 source.n78 source.n75 104.615
R188 source.n130 source.n129 104.615
R189 source.n129 source.n107 104.615
R190 source.n122 source.n107 104.615
R191 source.n122 source.n121 104.615
R192 source.n121 source.n111 104.615
R193 source.n114 source.n111 104.615
R194 source.n250 source.t18 52.3082
R195 source.n214 source.t14 52.3082
R196 source.n182 source.t3 52.3082
R197 source.n146 source.t11 52.3082
R198 source.n10 source.t10 52.3082
R199 source.n46 source.t0 52.3082
R200 source.n78 source.t16 52.3082
R201 source.n114 source.t22 52.3082
R202 source.n33 source.n32 50.512
R203 source.n35 source.n34 50.512
R204 source.n101 source.n100 50.512
R205 source.n103 source.n102 50.512
R206 source.n239 source.n238 50.5119
R207 source.n237 source.n236 50.5119
R208 source.n171 source.n170 50.5119
R209 source.n169 source.n168 50.5119
R210 source.n271 source.n270 32.1853
R211 source.n235 source.n234 32.1853
R212 source.n203 source.n202 32.1853
R213 source.n167 source.n166 32.1853
R214 source.n31 source.n30 32.1853
R215 source.n67 source.n66 32.1853
R216 source.n99 source.n98 32.1853
R217 source.n135 source.n134 32.1853
R218 source.n167 source.n135 17.2854
R219 source.n251 source.n249 15.6674
R220 source.n215 source.n213 15.6674
R221 source.n183 source.n181 15.6674
R222 source.n147 source.n145 15.6674
R223 source.n11 source.n9 15.6674
R224 source.n47 source.n45 15.6674
R225 source.n79 source.n77 15.6674
R226 source.n115 source.n113 15.6674
R227 source.n252 source.n248 12.8005
R228 source.n216 source.n212 12.8005
R229 source.n184 source.n180 12.8005
R230 source.n148 source.n144 12.8005
R231 source.n12 source.n8 12.8005
R232 source.n48 source.n44 12.8005
R233 source.n80 source.n76 12.8005
R234 source.n116 source.n112 12.8005
R235 source.n256 source.n255 12.0247
R236 source.n220 source.n219 12.0247
R237 source.n188 source.n187 12.0247
R238 source.n152 source.n151 12.0247
R239 source.n16 source.n15 12.0247
R240 source.n52 source.n51 12.0247
R241 source.n84 source.n83 12.0247
R242 source.n120 source.n119 12.0247
R243 source.n272 source.n31 11.7509
R244 source.n259 source.n246 11.249
R245 source.n223 source.n210 11.249
R246 source.n191 source.n178 11.249
R247 source.n155 source.n142 11.249
R248 source.n19 source.n6 11.249
R249 source.n55 source.n42 11.249
R250 source.n87 source.n74 11.249
R251 source.n123 source.n110 11.249
R252 source.n260 source.n244 10.4732
R253 source.n224 source.n208 10.4732
R254 source.n192 source.n176 10.4732
R255 source.n156 source.n140 10.4732
R256 source.n20 source.n4 10.4732
R257 source.n56 source.n40 10.4732
R258 source.n88 source.n72 10.4732
R259 source.n124 source.n108 10.4732
R260 source.n264 source.n263 9.69747
R261 source.n228 source.n227 9.69747
R262 source.n196 source.n195 9.69747
R263 source.n160 source.n159 9.69747
R264 source.n24 source.n23 9.69747
R265 source.n60 source.n59 9.69747
R266 source.n92 source.n91 9.69747
R267 source.n128 source.n127 9.69747
R268 source.n270 source.n269 9.45567
R269 source.n234 source.n233 9.45567
R270 source.n202 source.n201 9.45567
R271 source.n166 source.n165 9.45567
R272 source.n30 source.n29 9.45567
R273 source.n66 source.n65 9.45567
R274 source.n98 source.n97 9.45567
R275 source.n134 source.n133 9.45567
R276 source.n269 source.n268 9.3005
R277 source.n242 source.n241 9.3005
R278 source.n263 source.n262 9.3005
R279 source.n261 source.n260 9.3005
R280 source.n246 source.n245 9.3005
R281 source.n255 source.n254 9.3005
R282 source.n253 source.n252 9.3005
R283 source.n233 source.n232 9.3005
R284 source.n206 source.n205 9.3005
R285 source.n227 source.n226 9.3005
R286 source.n225 source.n224 9.3005
R287 source.n210 source.n209 9.3005
R288 source.n219 source.n218 9.3005
R289 source.n217 source.n216 9.3005
R290 source.n201 source.n200 9.3005
R291 source.n174 source.n173 9.3005
R292 source.n195 source.n194 9.3005
R293 source.n193 source.n192 9.3005
R294 source.n178 source.n177 9.3005
R295 source.n187 source.n186 9.3005
R296 source.n185 source.n184 9.3005
R297 source.n165 source.n164 9.3005
R298 source.n138 source.n137 9.3005
R299 source.n159 source.n158 9.3005
R300 source.n157 source.n156 9.3005
R301 source.n142 source.n141 9.3005
R302 source.n151 source.n150 9.3005
R303 source.n149 source.n148 9.3005
R304 source.n29 source.n28 9.3005
R305 source.n2 source.n1 9.3005
R306 source.n23 source.n22 9.3005
R307 source.n21 source.n20 9.3005
R308 source.n6 source.n5 9.3005
R309 source.n15 source.n14 9.3005
R310 source.n13 source.n12 9.3005
R311 source.n65 source.n64 9.3005
R312 source.n38 source.n37 9.3005
R313 source.n59 source.n58 9.3005
R314 source.n57 source.n56 9.3005
R315 source.n42 source.n41 9.3005
R316 source.n51 source.n50 9.3005
R317 source.n49 source.n48 9.3005
R318 source.n97 source.n96 9.3005
R319 source.n70 source.n69 9.3005
R320 source.n91 source.n90 9.3005
R321 source.n89 source.n88 9.3005
R322 source.n74 source.n73 9.3005
R323 source.n83 source.n82 9.3005
R324 source.n81 source.n80 9.3005
R325 source.n133 source.n132 9.3005
R326 source.n106 source.n105 9.3005
R327 source.n127 source.n126 9.3005
R328 source.n125 source.n124 9.3005
R329 source.n110 source.n109 9.3005
R330 source.n119 source.n118 9.3005
R331 source.n117 source.n116 9.3005
R332 source.n267 source.n242 8.92171
R333 source.n231 source.n206 8.92171
R334 source.n199 source.n174 8.92171
R335 source.n163 source.n138 8.92171
R336 source.n27 source.n2 8.92171
R337 source.n63 source.n38 8.92171
R338 source.n95 source.n70 8.92171
R339 source.n131 source.n106 8.92171
R340 source.n268 source.n240 8.14595
R341 source.n232 source.n204 8.14595
R342 source.n200 source.n172 8.14595
R343 source.n164 source.n136 8.14595
R344 source.n28 source.n0 8.14595
R345 source.n64 source.n36 8.14595
R346 source.n96 source.n68 8.14595
R347 source.n132 source.n104 8.14595
R348 source.n270 source.n240 5.81868
R349 source.n234 source.n204 5.81868
R350 source.n202 source.n172 5.81868
R351 source.n166 source.n136 5.81868
R352 source.n30 source.n0 5.81868
R353 source.n66 source.n36 5.81868
R354 source.n98 source.n68 5.81868
R355 source.n134 source.n104 5.81868
R356 source.n272 source.n271 5.53498
R357 source.n268 source.n267 5.04292
R358 source.n232 source.n231 5.04292
R359 source.n200 source.n199 5.04292
R360 source.n164 source.n163 5.04292
R361 source.n28 source.n27 5.04292
R362 source.n64 source.n63 5.04292
R363 source.n96 source.n95 5.04292
R364 source.n132 source.n131 5.04292
R365 source.n253 source.n249 4.38594
R366 source.n217 source.n213 4.38594
R367 source.n185 source.n181 4.38594
R368 source.n149 source.n145 4.38594
R369 source.n13 source.n9 4.38594
R370 source.n49 source.n45 4.38594
R371 source.n81 source.n77 4.38594
R372 source.n117 source.n113 4.38594
R373 source.n264 source.n242 4.26717
R374 source.n228 source.n206 4.26717
R375 source.n196 source.n174 4.26717
R376 source.n160 source.n138 4.26717
R377 source.n24 source.n2 4.26717
R378 source.n60 source.n38 4.26717
R379 source.n92 source.n70 4.26717
R380 source.n128 source.n106 4.26717
R381 source.n263 source.n244 3.49141
R382 source.n227 source.n208 3.49141
R383 source.n195 source.n176 3.49141
R384 source.n159 source.n140 3.49141
R385 source.n23 source.n4 3.49141
R386 source.n59 source.n40 3.49141
R387 source.n91 source.n72 3.49141
R388 source.n127 source.n108 3.49141
R389 source.n238 source.t20 3.3005
R390 source.n238 source.t23 3.3005
R391 source.n236 source.t19 3.3005
R392 source.n236 source.t15 3.3005
R393 source.n170 source.t7 3.3005
R394 source.n170 source.t9 3.3005
R395 source.n168 source.t6 3.3005
R396 source.n168 source.t8 3.3005
R397 source.n32 source.t5 3.3005
R398 source.n32 source.t1 3.3005
R399 source.n34 source.t2 3.3005
R400 source.n34 source.t4 3.3005
R401 source.n100 source.t21 3.3005
R402 source.n100 source.t12 3.3005
R403 source.n102 source.t13 3.3005
R404 source.n102 source.t17 3.3005
R405 source.n260 source.n259 2.71565
R406 source.n224 source.n223 2.71565
R407 source.n192 source.n191 2.71565
R408 source.n156 source.n155 2.71565
R409 source.n20 source.n19 2.71565
R410 source.n56 source.n55 2.71565
R411 source.n88 source.n87 2.71565
R412 source.n124 source.n123 2.71565
R413 source.n256 source.n246 1.93989
R414 source.n220 source.n210 1.93989
R415 source.n188 source.n178 1.93989
R416 source.n152 source.n142 1.93989
R417 source.n16 source.n6 1.93989
R418 source.n52 source.n42 1.93989
R419 source.n84 source.n74 1.93989
R420 source.n120 source.n110 1.93989
R421 source.n255 source.n248 1.16414
R422 source.n219 source.n212 1.16414
R423 source.n187 source.n180 1.16414
R424 source.n151 source.n144 1.16414
R425 source.n15 source.n8 1.16414
R426 source.n51 source.n44 1.16414
R427 source.n83 source.n76 1.16414
R428 source.n119 source.n112 1.16414
R429 source.n135 source.n103 0.543603
R430 source.n103 source.n101 0.543603
R431 source.n101 source.n99 0.543603
R432 source.n67 source.n35 0.543603
R433 source.n35 source.n33 0.543603
R434 source.n33 source.n31 0.543603
R435 source.n169 source.n167 0.543603
R436 source.n171 source.n169 0.543603
R437 source.n203 source.n171 0.543603
R438 source.n237 source.n235 0.543603
R439 source.n239 source.n237 0.543603
R440 source.n271 source.n239 0.543603
R441 source.n99 source.n67 0.470328
R442 source.n235 source.n203 0.470328
R443 source.n252 source.n251 0.388379
R444 source.n216 source.n215 0.388379
R445 source.n184 source.n183 0.388379
R446 source.n148 source.n147 0.388379
R447 source.n12 source.n11 0.388379
R448 source.n48 source.n47 0.388379
R449 source.n80 source.n79 0.388379
R450 source.n116 source.n115 0.388379
R451 source source.n272 0.188
R452 source.n254 source.n253 0.155672
R453 source.n254 source.n245 0.155672
R454 source.n261 source.n245 0.155672
R455 source.n262 source.n261 0.155672
R456 source.n262 source.n241 0.155672
R457 source.n269 source.n241 0.155672
R458 source.n218 source.n217 0.155672
R459 source.n218 source.n209 0.155672
R460 source.n225 source.n209 0.155672
R461 source.n226 source.n225 0.155672
R462 source.n226 source.n205 0.155672
R463 source.n233 source.n205 0.155672
R464 source.n186 source.n185 0.155672
R465 source.n186 source.n177 0.155672
R466 source.n193 source.n177 0.155672
R467 source.n194 source.n193 0.155672
R468 source.n194 source.n173 0.155672
R469 source.n201 source.n173 0.155672
R470 source.n150 source.n149 0.155672
R471 source.n150 source.n141 0.155672
R472 source.n157 source.n141 0.155672
R473 source.n158 source.n157 0.155672
R474 source.n158 source.n137 0.155672
R475 source.n165 source.n137 0.155672
R476 source.n29 source.n1 0.155672
R477 source.n22 source.n1 0.155672
R478 source.n22 source.n21 0.155672
R479 source.n21 source.n5 0.155672
R480 source.n14 source.n5 0.155672
R481 source.n14 source.n13 0.155672
R482 source.n65 source.n37 0.155672
R483 source.n58 source.n37 0.155672
R484 source.n58 source.n57 0.155672
R485 source.n57 source.n41 0.155672
R486 source.n50 source.n41 0.155672
R487 source.n50 source.n49 0.155672
R488 source.n97 source.n69 0.155672
R489 source.n90 source.n69 0.155672
R490 source.n90 source.n89 0.155672
R491 source.n89 source.n73 0.155672
R492 source.n82 source.n73 0.155672
R493 source.n82 source.n81 0.155672
R494 source.n133 source.n105 0.155672
R495 source.n126 source.n105 0.155672
R496 source.n126 source.n125 0.155672
R497 source.n125 source.n109 0.155672
R498 source.n118 source.n109 0.155672
R499 source.n118 source.n117 0.155672
R500 plus.n2 plus.t1 633.904
R501 plus.n13 plus.t8 633.904
R502 plus.n17 plus.t6 633.904
R503 plus.n28 plus.t3 633.904
R504 plus.n3 plus.t5 586.433
R505 plus.n4 plus.t9 586.433
R506 plus.n10 plus.t11 586.433
R507 plus.n12 plus.t4 586.433
R508 plus.n19 plus.t0 586.433
R509 plus.n18 plus.t7 586.433
R510 plus.n25 plus.t2 586.433
R511 plus.n27 plus.t10 586.433
R512 plus.n6 plus.n2 161.489
R513 plus.n21 plus.n17 161.489
R514 plus.n6 plus.n5 161.3
R515 plus.n7 plus.n1 161.3
R516 plus.n9 plus.n8 161.3
R517 plus.n11 plus.n0 161.3
R518 plus.n14 plus.n13 161.3
R519 plus.n21 plus.n20 161.3
R520 plus.n22 plus.n16 161.3
R521 plus.n24 plus.n23 161.3
R522 plus.n26 plus.n15 161.3
R523 plus.n29 plus.n28 161.3
R524 plus.n9 plus.n1 73.0308
R525 plus.n24 plus.n16 73.0308
R526 plus.n5 plus.n4 63.5369
R527 plus.n11 plus.n10 63.5369
R528 plus.n26 plus.n25 63.5369
R529 plus.n20 plus.n18 63.5369
R530 plus.n3 plus.n2 44.549
R531 plus.n13 plus.n12 44.549
R532 plus.n28 plus.n27 44.549
R533 plus.n19 plus.n17 44.549
R534 plus.n5 plus.n3 28.4823
R535 plus.n12 plus.n11 28.4823
R536 plus.n27 plus.n26 28.4823
R537 plus.n20 plus.n19 28.4823
R538 plus plus.n29 26.7945
R539 plus plus.n14 9.88308
R540 plus.n4 plus.n1 9.49444
R541 plus.n10 plus.n9 9.49444
R542 plus.n25 plus.n24 9.49444
R543 plus.n18 plus.n16 9.49444
R544 plus.n7 plus.n6 0.189894
R545 plus.n8 plus.n7 0.189894
R546 plus.n8 plus.n0 0.189894
R547 plus.n14 plus.n0 0.189894
R548 plus.n29 plus.n15 0.189894
R549 plus.n23 plus.n15 0.189894
R550 plus.n23 plus.n22 0.189894
R551 plus.n22 plus.n21 0.189894
R552 drain_left.n6 drain_left.n4 67.7339
R553 drain_left.n3 drain_left.n2 67.6784
R554 drain_left.n3 drain_left.n0 67.6784
R555 drain_left.n6 drain_left.n5 67.1908
R556 drain_left.n8 drain_left.n7 67.1907
R557 drain_left.n3 drain_left.n1 67.1907
R558 drain_left drain_left.n3 25.5371
R559 drain_left drain_left.n8 6.19632
R560 drain_left.n1 drain_left.t9 3.3005
R561 drain_left.n1 drain_left.t4 3.3005
R562 drain_left.n2 drain_left.t11 3.3005
R563 drain_left.n2 drain_left.t5 3.3005
R564 drain_left.n0 drain_left.t8 3.3005
R565 drain_left.n0 drain_left.t1 3.3005
R566 drain_left.n7 drain_left.t7 3.3005
R567 drain_left.n7 drain_left.t3 3.3005
R568 drain_left.n5 drain_left.t2 3.3005
R569 drain_left.n5 drain_left.t0 3.3005
R570 drain_left.n4 drain_left.t10 3.3005
R571 drain_left.n4 drain_left.t6 3.3005
R572 drain_left.n8 drain_left.n6 0.543603
C0 drain_right source 12.919701f
C1 drain_left source 12.9199f
C2 drain_right drain_left 0.785787f
C3 minus source 2.46494f
C4 minus drain_right 2.53958f
C5 minus drain_left 0.170859f
C6 plus source 2.47896f
C7 plus drain_right 0.30725f
C8 plus drain_left 2.69304f
C9 plus minus 4.03242f
C10 drain_right a_n1598_n2088# 4.78196f
C11 drain_left a_n1598_n2088# 5.04244f
C12 source a_n1598_n2088# 5.244471f
C13 minus a_n1598_n2088# 5.73127f
C14 plus a_n1598_n2088# 7.30073f
C15 drain_left.t8 a_n1598_n2088# 0.155405f
C16 drain_left.t1 a_n1598_n2088# 0.155405f
C17 drain_left.n0 a_n1598_n2088# 1.29889f
C18 drain_left.t9 a_n1598_n2088# 0.155405f
C19 drain_left.t4 a_n1598_n2088# 0.155405f
C20 drain_left.n1 a_n1598_n2088# 1.29608f
C21 drain_left.t11 a_n1598_n2088# 0.155405f
C22 drain_left.t5 a_n1598_n2088# 0.155405f
C23 drain_left.n2 a_n1598_n2088# 1.29889f
C24 drain_left.n3 a_n1598_n2088# 2.19616f
C25 drain_left.t10 a_n1598_n2088# 0.155405f
C26 drain_left.t6 a_n1598_n2088# 0.155405f
C27 drain_left.n4 a_n1598_n2088# 1.29925f
C28 drain_left.t2 a_n1598_n2088# 0.155405f
C29 drain_left.t0 a_n1598_n2088# 0.155405f
C30 drain_left.n5 a_n1598_n2088# 1.29609f
C31 drain_left.n6 a_n1598_n2088# 0.771515f
C32 drain_left.t7 a_n1598_n2088# 0.155405f
C33 drain_left.t3 a_n1598_n2088# 0.155405f
C34 drain_left.n7 a_n1598_n2088# 1.29608f
C35 drain_left.n8 a_n1598_n2088# 0.65356f
C36 plus.n0 a_n1598_n2088# 0.053851f
C37 plus.t4 a_n1598_n2088# 0.276178f
C38 plus.t11 a_n1598_n2088# 0.276178f
C39 plus.n1 a_n1598_n2088# 0.020022f
C40 plus.t1 a_n1598_n2088# 0.285982f
C41 plus.n2 a_n1598_n2088# 0.143378f
C42 plus.t5 a_n1598_n2088# 0.276178f
C43 plus.n3 a_n1598_n2088# 0.12677f
C44 plus.t9 a_n1598_n2088# 0.276178f
C45 plus.n4 a_n1598_n2088# 0.12677f
C46 plus.n5 a_n1598_n2088# 0.022181f
C47 plus.n6 a_n1598_n2088# 0.122563f
C48 plus.n7 a_n1598_n2088# 0.053851f
C49 plus.n8 a_n1598_n2088# 0.053851f
C50 plus.n9 a_n1598_n2088# 0.020022f
C51 plus.n10 a_n1598_n2088# 0.12677f
C52 plus.n11 a_n1598_n2088# 0.022181f
C53 plus.n12 a_n1598_n2088# 0.12677f
C54 plus.t8 a_n1598_n2088# 0.285982f
C55 plus.n13 a_n1598_n2088# 0.143297f
C56 plus.n14 a_n1598_n2088# 0.463019f
C57 plus.n15 a_n1598_n2088# 0.053851f
C58 plus.t3 a_n1598_n2088# 0.285982f
C59 plus.t10 a_n1598_n2088# 0.276178f
C60 plus.t2 a_n1598_n2088# 0.276178f
C61 plus.n16 a_n1598_n2088# 0.020022f
C62 plus.t6 a_n1598_n2088# 0.285982f
C63 plus.n17 a_n1598_n2088# 0.143378f
C64 plus.t7 a_n1598_n2088# 0.276178f
C65 plus.n18 a_n1598_n2088# 0.12677f
C66 plus.t0 a_n1598_n2088# 0.276178f
C67 plus.n19 a_n1598_n2088# 0.12677f
C68 plus.n20 a_n1598_n2088# 0.022181f
C69 plus.n21 a_n1598_n2088# 0.122563f
C70 plus.n22 a_n1598_n2088# 0.053851f
C71 plus.n23 a_n1598_n2088# 0.053851f
C72 plus.n24 a_n1598_n2088# 0.020022f
C73 plus.n25 a_n1598_n2088# 0.12677f
C74 plus.n26 a_n1598_n2088# 0.022181f
C75 plus.n27 a_n1598_n2088# 0.12677f
C76 plus.n28 a_n1598_n2088# 0.143297f
C77 plus.n29 a_n1598_n2088# 1.31274f
C78 source.n0 a_n1598_n2088# 0.039054f
C79 source.n1 a_n1598_n2088# 0.027785f
C80 source.n2 a_n1598_n2088# 0.01493f
C81 source.n3 a_n1598_n2088# 0.035289f
C82 source.n4 a_n1598_n2088# 0.015808f
C83 source.n5 a_n1598_n2088# 0.027785f
C84 source.n6 a_n1598_n2088# 0.01493f
C85 source.n7 a_n1598_n2088# 0.035289f
C86 source.n8 a_n1598_n2088# 0.015808f
C87 source.n9 a_n1598_n2088# 0.118898f
C88 source.t10 a_n1598_n2088# 0.057517f
C89 source.n10 a_n1598_n2088# 0.026467f
C90 source.n11 a_n1598_n2088# 0.020845f
C91 source.n12 a_n1598_n2088# 0.01493f
C92 source.n13 a_n1598_n2088# 0.661105f
C93 source.n14 a_n1598_n2088# 0.027785f
C94 source.n15 a_n1598_n2088# 0.01493f
C95 source.n16 a_n1598_n2088# 0.015808f
C96 source.n17 a_n1598_n2088# 0.035289f
C97 source.n18 a_n1598_n2088# 0.035289f
C98 source.n19 a_n1598_n2088# 0.015808f
C99 source.n20 a_n1598_n2088# 0.01493f
C100 source.n21 a_n1598_n2088# 0.027785f
C101 source.n22 a_n1598_n2088# 0.027785f
C102 source.n23 a_n1598_n2088# 0.01493f
C103 source.n24 a_n1598_n2088# 0.015808f
C104 source.n25 a_n1598_n2088# 0.035289f
C105 source.n26 a_n1598_n2088# 0.076396f
C106 source.n27 a_n1598_n2088# 0.015808f
C107 source.n28 a_n1598_n2088# 0.01493f
C108 source.n29 a_n1598_n2088# 0.064222f
C109 source.n30 a_n1598_n2088# 0.042746f
C110 source.n31 a_n1598_n2088# 0.672995f
C111 source.t5 a_n1598_n2088# 0.131737f
C112 source.t1 a_n1598_n2088# 0.131737f
C113 source.n32 a_n1598_n2088# 1.02598f
C114 source.n33 a_n1598_n2088# 0.357698f
C115 source.t2 a_n1598_n2088# 0.131737f
C116 source.t4 a_n1598_n2088# 0.131737f
C117 source.n34 a_n1598_n2088# 1.02598f
C118 source.n35 a_n1598_n2088# 0.357698f
C119 source.n36 a_n1598_n2088# 0.039054f
C120 source.n37 a_n1598_n2088# 0.027785f
C121 source.n38 a_n1598_n2088# 0.01493f
C122 source.n39 a_n1598_n2088# 0.035289f
C123 source.n40 a_n1598_n2088# 0.015808f
C124 source.n41 a_n1598_n2088# 0.027785f
C125 source.n42 a_n1598_n2088# 0.01493f
C126 source.n43 a_n1598_n2088# 0.035289f
C127 source.n44 a_n1598_n2088# 0.015808f
C128 source.n45 a_n1598_n2088# 0.118898f
C129 source.t0 a_n1598_n2088# 0.057517f
C130 source.n46 a_n1598_n2088# 0.026467f
C131 source.n47 a_n1598_n2088# 0.020845f
C132 source.n48 a_n1598_n2088# 0.01493f
C133 source.n49 a_n1598_n2088# 0.661105f
C134 source.n50 a_n1598_n2088# 0.027785f
C135 source.n51 a_n1598_n2088# 0.01493f
C136 source.n52 a_n1598_n2088# 0.015808f
C137 source.n53 a_n1598_n2088# 0.035289f
C138 source.n54 a_n1598_n2088# 0.035289f
C139 source.n55 a_n1598_n2088# 0.015808f
C140 source.n56 a_n1598_n2088# 0.01493f
C141 source.n57 a_n1598_n2088# 0.027785f
C142 source.n58 a_n1598_n2088# 0.027785f
C143 source.n59 a_n1598_n2088# 0.01493f
C144 source.n60 a_n1598_n2088# 0.015808f
C145 source.n61 a_n1598_n2088# 0.035289f
C146 source.n62 a_n1598_n2088# 0.076396f
C147 source.n63 a_n1598_n2088# 0.015808f
C148 source.n64 a_n1598_n2088# 0.01493f
C149 source.n65 a_n1598_n2088# 0.064222f
C150 source.n66 a_n1598_n2088# 0.042746f
C151 source.n67 a_n1598_n2088# 0.114415f
C152 source.n68 a_n1598_n2088# 0.039054f
C153 source.n69 a_n1598_n2088# 0.027785f
C154 source.n70 a_n1598_n2088# 0.01493f
C155 source.n71 a_n1598_n2088# 0.035289f
C156 source.n72 a_n1598_n2088# 0.015808f
C157 source.n73 a_n1598_n2088# 0.027785f
C158 source.n74 a_n1598_n2088# 0.01493f
C159 source.n75 a_n1598_n2088# 0.035289f
C160 source.n76 a_n1598_n2088# 0.015808f
C161 source.n77 a_n1598_n2088# 0.118898f
C162 source.t16 a_n1598_n2088# 0.057517f
C163 source.n78 a_n1598_n2088# 0.026467f
C164 source.n79 a_n1598_n2088# 0.020845f
C165 source.n80 a_n1598_n2088# 0.01493f
C166 source.n81 a_n1598_n2088# 0.661105f
C167 source.n82 a_n1598_n2088# 0.027785f
C168 source.n83 a_n1598_n2088# 0.01493f
C169 source.n84 a_n1598_n2088# 0.015808f
C170 source.n85 a_n1598_n2088# 0.035289f
C171 source.n86 a_n1598_n2088# 0.035289f
C172 source.n87 a_n1598_n2088# 0.015808f
C173 source.n88 a_n1598_n2088# 0.01493f
C174 source.n89 a_n1598_n2088# 0.027785f
C175 source.n90 a_n1598_n2088# 0.027785f
C176 source.n91 a_n1598_n2088# 0.01493f
C177 source.n92 a_n1598_n2088# 0.015808f
C178 source.n93 a_n1598_n2088# 0.035289f
C179 source.n94 a_n1598_n2088# 0.076396f
C180 source.n95 a_n1598_n2088# 0.015808f
C181 source.n96 a_n1598_n2088# 0.01493f
C182 source.n97 a_n1598_n2088# 0.064222f
C183 source.n98 a_n1598_n2088# 0.042746f
C184 source.n99 a_n1598_n2088# 0.114415f
C185 source.t21 a_n1598_n2088# 0.131737f
C186 source.t12 a_n1598_n2088# 0.131737f
C187 source.n100 a_n1598_n2088# 1.02598f
C188 source.n101 a_n1598_n2088# 0.357698f
C189 source.t13 a_n1598_n2088# 0.131737f
C190 source.t17 a_n1598_n2088# 0.131737f
C191 source.n102 a_n1598_n2088# 1.02598f
C192 source.n103 a_n1598_n2088# 0.357698f
C193 source.n104 a_n1598_n2088# 0.039054f
C194 source.n105 a_n1598_n2088# 0.027785f
C195 source.n106 a_n1598_n2088# 0.01493f
C196 source.n107 a_n1598_n2088# 0.035289f
C197 source.n108 a_n1598_n2088# 0.015808f
C198 source.n109 a_n1598_n2088# 0.027785f
C199 source.n110 a_n1598_n2088# 0.01493f
C200 source.n111 a_n1598_n2088# 0.035289f
C201 source.n112 a_n1598_n2088# 0.015808f
C202 source.n113 a_n1598_n2088# 0.118898f
C203 source.t22 a_n1598_n2088# 0.057517f
C204 source.n114 a_n1598_n2088# 0.026467f
C205 source.n115 a_n1598_n2088# 0.020845f
C206 source.n116 a_n1598_n2088# 0.01493f
C207 source.n117 a_n1598_n2088# 0.661105f
C208 source.n118 a_n1598_n2088# 0.027785f
C209 source.n119 a_n1598_n2088# 0.01493f
C210 source.n120 a_n1598_n2088# 0.015808f
C211 source.n121 a_n1598_n2088# 0.035289f
C212 source.n122 a_n1598_n2088# 0.035289f
C213 source.n123 a_n1598_n2088# 0.015808f
C214 source.n124 a_n1598_n2088# 0.01493f
C215 source.n125 a_n1598_n2088# 0.027785f
C216 source.n126 a_n1598_n2088# 0.027785f
C217 source.n127 a_n1598_n2088# 0.01493f
C218 source.n128 a_n1598_n2088# 0.015808f
C219 source.n129 a_n1598_n2088# 0.035289f
C220 source.n130 a_n1598_n2088# 0.076396f
C221 source.n131 a_n1598_n2088# 0.015808f
C222 source.n132 a_n1598_n2088# 0.01493f
C223 source.n133 a_n1598_n2088# 0.064222f
C224 source.n134 a_n1598_n2088# 0.042746f
C225 source.n135 a_n1598_n2088# 1.03069f
C226 source.n136 a_n1598_n2088# 0.039054f
C227 source.n137 a_n1598_n2088# 0.027785f
C228 source.n138 a_n1598_n2088# 0.01493f
C229 source.n139 a_n1598_n2088# 0.035289f
C230 source.n140 a_n1598_n2088# 0.015808f
C231 source.n141 a_n1598_n2088# 0.027785f
C232 source.n142 a_n1598_n2088# 0.01493f
C233 source.n143 a_n1598_n2088# 0.035289f
C234 source.n144 a_n1598_n2088# 0.015808f
C235 source.n145 a_n1598_n2088# 0.118898f
C236 source.t11 a_n1598_n2088# 0.057517f
C237 source.n146 a_n1598_n2088# 0.026467f
C238 source.n147 a_n1598_n2088# 0.020845f
C239 source.n148 a_n1598_n2088# 0.01493f
C240 source.n149 a_n1598_n2088# 0.661105f
C241 source.n150 a_n1598_n2088# 0.027785f
C242 source.n151 a_n1598_n2088# 0.01493f
C243 source.n152 a_n1598_n2088# 0.015808f
C244 source.n153 a_n1598_n2088# 0.035289f
C245 source.n154 a_n1598_n2088# 0.035289f
C246 source.n155 a_n1598_n2088# 0.015808f
C247 source.n156 a_n1598_n2088# 0.01493f
C248 source.n157 a_n1598_n2088# 0.027785f
C249 source.n158 a_n1598_n2088# 0.027785f
C250 source.n159 a_n1598_n2088# 0.01493f
C251 source.n160 a_n1598_n2088# 0.015808f
C252 source.n161 a_n1598_n2088# 0.035289f
C253 source.n162 a_n1598_n2088# 0.076396f
C254 source.n163 a_n1598_n2088# 0.015808f
C255 source.n164 a_n1598_n2088# 0.01493f
C256 source.n165 a_n1598_n2088# 0.064222f
C257 source.n166 a_n1598_n2088# 0.042746f
C258 source.n167 a_n1598_n2088# 1.03069f
C259 source.t6 a_n1598_n2088# 0.131737f
C260 source.t8 a_n1598_n2088# 0.131737f
C261 source.n168 a_n1598_n2088# 1.02597f
C262 source.n169 a_n1598_n2088# 0.357706f
C263 source.t7 a_n1598_n2088# 0.131737f
C264 source.t9 a_n1598_n2088# 0.131737f
C265 source.n170 a_n1598_n2088# 1.02597f
C266 source.n171 a_n1598_n2088# 0.357706f
C267 source.n172 a_n1598_n2088# 0.039054f
C268 source.n173 a_n1598_n2088# 0.027785f
C269 source.n174 a_n1598_n2088# 0.01493f
C270 source.n175 a_n1598_n2088# 0.035289f
C271 source.n176 a_n1598_n2088# 0.015808f
C272 source.n177 a_n1598_n2088# 0.027785f
C273 source.n178 a_n1598_n2088# 0.01493f
C274 source.n179 a_n1598_n2088# 0.035289f
C275 source.n180 a_n1598_n2088# 0.015808f
C276 source.n181 a_n1598_n2088# 0.118898f
C277 source.t3 a_n1598_n2088# 0.057517f
C278 source.n182 a_n1598_n2088# 0.026467f
C279 source.n183 a_n1598_n2088# 0.020845f
C280 source.n184 a_n1598_n2088# 0.01493f
C281 source.n185 a_n1598_n2088# 0.661105f
C282 source.n186 a_n1598_n2088# 0.027785f
C283 source.n187 a_n1598_n2088# 0.01493f
C284 source.n188 a_n1598_n2088# 0.015808f
C285 source.n189 a_n1598_n2088# 0.035289f
C286 source.n190 a_n1598_n2088# 0.035289f
C287 source.n191 a_n1598_n2088# 0.015808f
C288 source.n192 a_n1598_n2088# 0.01493f
C289 source.n193 a_n1598_n2088# 0.027785f
C290 source.n194 a_n1598_n2088# 0.027785f
C291 source.n195 a_n1598_n2088# 0.01493f
C292 source.n196 a_n1598_n2088# 0.015808f
C293 source.n197 a_n1598_n2088# 0.035289f
C294 source.n198 a_n1598_n2088# 0.076396f
C295 source.n199 a_n1598_n2088# 0.015808f
C296 source.n200 a_n1598_n2088# 0.01493f
C297 source.n201 a_n1598_n2088# 0.064222f
C298 source.n202 a_n1598_n2088# 0.042746f
C299 source.n203 a_n1598_n2088# 0.114415f
C300 source.n204 a_n1598_n2088# 0.039054f
C301 source.n205 a_n1598_n2088# 0.027785f
C302 source.n206 a_n1598_n2088# 0.01493f
C303 source.n207 a_n1598_n2088# 0.035289f
C304 source.n208 a_n1598_n2088# 0.015808f
C305 source.n209 a_n1598_n2088# 0.027785f
C306 source.n210 a_n1598_n2088# 0.01493f
C307 source.n211 a_n1598_n2088# 0.035289f
C308 source.n212 a_n1598_n2088# 0.015808f
C309 source.n213 a_n1598_n2088# 0.118898f
C310 source.t14 a_n1598_n2088# 0.057517f
C311 source.n214 a_n1598_n2088# 0.026467f
C312 source.n215 a_n1598_n2088# 0.020845f
C313 source.n216 a_n1598_n2088# 0.01493f
C314 source.n217 a_n1598_n2088# 0.661105f
C315 source.n218 a_n1598_n2088# 0.027785f
C316 source.n219 a_n1598_n2088# 0.01493f
C317 source.n220 a_n1598_n2088# 0.015808f
C318 source.n221 a_n1598_n2088# 0.035289f
C319 source.n222 a_n1598_n2088# 0.035289f
C320 source.n223 a_n1598_n2088# 0.015808f
C321 source.n224 a_n1598_n2088# 0.01493f
C322 source.n225 a_n1598_n2088# 0.027785f
C323 source.n226 a_n1598_n2088# 0.027785f
C324 source.n227 a_n1598_n2088# 0.01493f
C325 source.n228 a_n1598_n2088# 0.015808f
C326 source.n229 a_n1598_n2088# 0.035289f
C327 source.n230 a_n1598_n2088# 0.076396f
C328 source.n231 a_n1598_n2088# 0.015808f
C329 source.n232 a_n1598_n2088# 0.01493f
C330 source.n233 a_n1598_n2088# 0.064222f
C331 source.n234 a_n1598_n2088# 0.042746f
C332 source.n235 a_n1598_n2088# 0.114415f
C333 source.t19 a_n1598_n2088# 0.131737f
C334 source.t15 a_n1598_n2088# 0.131737f
C335 source.n236 a_n1598_n2088# 1.02597f
C336 source.n237 a_n1598_n2088# 0.357706f
C337 source.t20 a_n1598_n2088# 0.131737f
C338 source.t23 a_n1598_n2088# 0.131737f
C339 source.n238 a_n1598_n2088# 1.02597f
C340 source.n239 a_n1598_n2088# 0.357706f
C341 source.n240 a_n1598_n2088# 0.039054f
C342 source.n241 a_n1598_n2088# 0.027785f
C343 source.n242 a_n1598_n2088# 0.01493f
C344 source.n243 a_n1598_n2088# 0.035289f
C345 source.n244 a_n1598_n2088# 0.015808f
C346 source.n245 a_n1598_n2088# 0.027785f
C347 source.n246 a_n1598_n2088# 0.01493f
C348 source.n247 a_n1598_n2088# 0.035289f
C349 source.n248 a_n1598_n2088# 0.015808f
C350 source.n249 a_n1598_n2088# 0.118898f
C351 source.t18 a_n1598_n2088# 0.057517f
C352 source.n250 a_n1598_n2088# 0.026467f
C353 source.n251 a_n1598_n2088# 0.020845f
C354 source.n252 a_n1598_n2088# 0.01493f
C355 source.n253 a_n1598_n2088# 0.661105f
C356 source.n254 a_n1598_n2088# 0.027785f
C357 source.n255 a_n1598_n2088# 0.01493f
C358 source.n256 a_n1598_n2088# 0.015808f
C359 source.n257 a_n1598_n2088# 0.035289f
C360 source.n258 a_n1598_n2088# 0.035289f
C361 source.n259 a_n1598_n2088# 0.015808f
C362 source.n260 a_n1598_n2088# 0.01493f
C363 source.n261 a_n1598_n2088# 0.027785f
C364 source.n262 a_n1598_n2088# 0.027785f
C365 source.n263 a_n1598_n2088# 0.01493f
C366 source.n264 a_n1598_n2088# 0.015808f
C367 source.n265 a_n1598_n2088# 0.035289f
C368 source.n266 a_n1598_n2088# 0.076396f
C369 source.n267 a_n1598_n2088# 0.015808f
C370 source.n268 a_n1598_n2088# 0.01493f
C371 source.n269 a_n1598_n2088# 0.064222f
C372 source.n270 a_n1598_n2088# 0.042746f
C373 source.n271 a_n1598_n2088# 0.271259f
C374 source.n272 a_n1598_n2088# 1.13689f
C375 drain_right.t9 a_n1598_n2088# 0.154684f
C376 drain_right.t8 a_n1598_n2088# 0.154684f
C377 drain_right.n0 a_n1598_n2088# 1.29286f
C378 drain_right.t0 a_n1598_n2088# 0.154684f
C379 drain_right.t11 a_n1598_n2088# 0.154684f
C380 drain_right.n1 a_n1598_n2088# 1.29007f
C381 drain_right.t10 a_n1598_n2088# 0.154684f
C382 drain_right.t2 a_n1598_n2088# 0.154684f
C383 drain_right.n2 a_n1598_n2088# 1.29286f
C384 drain_right.n3 a_n1598_n2088# 2.11948f
C385 drain_right.t3 a_n1598_n2088# 0.154684f
C386 drain_right.t4 a_n1598_n2088# 0.154684f
C387 drain_right.n4 a_n1598_n2088# 1.29321f
C388 drain_right.t7 a_n1598_n2088# 0.154684f
C389 drain_right.t6 a_n1598_n2088# 0.154684f
C390 drain_right.n5 a_n1598_n2088# 1.29007f
C391 drain_right.n6 a_n1598_n2088# 0.767942f
C392 drain_right.t1 a_n1598_n2088# 0.154684f
C393 drain_right.t5 a_n1598_n2088# 0.154684f
C394 drain_right.n7 a_n1598_n2088# 1.29007f
C395 drain_right.n8 a_n1598_n2088# 0.650522f
C396 minus.n0 a_n1598_n2088# 0.052064f
C397 minus.t1 a_n1598_n2088# 0.276492f
C398 minus.t10 a_n1598_n2088# 0.267014f
C399 minus.t6 a_n1598_n2088# 0.267014f
C400 minus.n1 a_n1598_n2088# 0.019358f
C401 minus.t7 a_n1598_n2088# 0.276492f
C402 minus.n2 a_n1598_n2088# 0.13862f
C403 minus.t2 a_n1598_n2088# 0.267014f
C404 minus.n3 a_n1598_n2088# 0.122564f
C405 minus.t11 a_n1598_n2088# 0.267014f
C406 minus.n4 a_n1598_n2088# 0.122564f
C407 minus.n5 a_n1598_n2088# 0.021444f
C408 minus.n6 a_n1598_n2088# 0.118496f
C409 minus.n7 a_n1598_n2088# 0.052064f
C410 minus.n8 a_n1598_n2088# 0.052064f
C411 minus.n9 a_n1598_n2088# 0.019358f
C412 minus.n10 a_n1598_n2088# 0.122564f
C413 minus.n11 a_n1598_n2088# 0.021444f
C414 minus.n12 a_n1598_n2088# 0.122564f
C415 minus.n13 a_n1598_n2088# 0.138542f
C416 minus.n14 a_n1598_n2088# 1.40447f
C417 minus.n15 a_n1598_n2088# 0.052064f
C418 minus.t0 a_n1598_n2088# 0.267014f
C419 minus.t3 a_n1598_n2088# 0.267014f
C420 minus.n16 a_n1598_n2088# 0.019358f
C421 minus.t9 a_n1598_n2088# 0.276492f
C422 minus.n17 a_n1598_n2088# 0.13862f
C423 minus.t4 a_n1598_n2088# 0.267014f
C424 minus.n18 a_n1598_n2088# 0.122564f
C425 minus.t8 a_n1598_n2088# 0.267014f
C426 minus.n19 a_n1598_n2088# 0.122564f
C427 minus.n20 a_n1598_n2088# 0.021444f
C428 minus.n21 a_n1598_n2088# 0.118496f
C429 minus.n22 a_n1598_n2088# 0.052064f
C430 minus.n23 a_n1598_n2088# 0.052064f
C431 minus.n24 a_n1598_n2088# 0.019358f
C432 minus.n25 a_n1598_n2088# 0.122564f
C433 minus.n26 a_n1598_n2088# 0.021444f
C434 minus.n27 a_n1598_n2088# 0.122564f
C435 minus.t5 a_n1598_n2088# 0.276492f
C436 minus.n28 a_n1598_n2088# 0.138542f
C437 minus.n29 a_n1598_n2088# 0.341839f
C438 minus.n30 a_n1598_n2088# 1.73f
.ends

