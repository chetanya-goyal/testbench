* NGSPICE file created from diffpair308.ext - technology: sky130A

.subckt diffpair308 minus drain_right drain_left source plus
X0 source.t39 plus.t0 drain_left.t10 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X1 source.t38 plus.t1 drain_left.t5 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X2 source.t37 plus.t2 drain_left.t8 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X3 source.t5 minus.t0 drain_right.t19 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X4 drain_left.t3 plus.t3 source.t36 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X5 a_n2982_n2088# a_n2982_n2088# a_n2982_n2088# a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.7
X6 drain_left.t11 plus.t4 source.t35 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X7 source.t34 plus.t5 drain_left.t6 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X8 source.t33 plus.t6 drain_left.t16 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X9 a_n2982_n2088# a_n2982_n2088# a_n2982_n2088# a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X10 source.t1 minus.t1 drain_right.t18 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X11 drain_right.t17 minus.t2 source.t2 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X12 drain_left.t17 plus.t7 source.t32 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X13 source.t31 plus.t8 drain_left.t9 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X14 drain_right.t16 minus.t3 source.t7 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X15 drain_left.t0 plus.t9 source.t30 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X16 drain_right.t15 minus.t4 source.t13 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X17 drain_right.t14 minus.t5 source.t8 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X18 drain_right.t13 minus.t6 source.t18 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X19 source.t19 minus.t7 drain_right.t12 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X20 source.t29 plus.t10 drain_left.t14 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X21 drain_left.t1 plus.t11 source.t28 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X22 drain_left.t4 plus.t12 source.t27 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X23 drain_right.t11 minus.t8 source.t9 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X24 source.t15 minus.t9 drain_right.t10 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X25 source.t26 plus.t13 drain_left.t18 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X26 drain_left.t15 plus.t14 source.t25 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X27 drain_right.t9 minus.t10 source.t17 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X28 drain_left.t19 plus.t15 source.t24 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X29 drain_right.t8 minus.t11 source.t6 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X30 source.t16 minus.t12 drain_right.t7 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X31 drain_left.t12 plus.t16 source.t23 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X32 source.t22 plus.t17 drain_left.t13 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X33 drain_left.t7 plus.t18 source.t21 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X34 a_n2982_n2088# a_n2982_n2088# a_n2982_n2088# a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X35 source.t10 minus.t13 drain_right.t6 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X36 source.t14 minus.t14 drain_right.t5 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X37 drain_right.t4 minus.t15 source.t12 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X38 source.t3 minus.t16 drain_right.t3 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X39 a_n2982_n2088# a_n2982_n2088# a_n2982_n2088# a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X40 drain_right.t2 minus.t17 source.t4 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X41 source.t0 minus.t18 drain_right.t1 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X42 source.t11 minus.t19 drain_right.t0 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X43 source.t20 plus.t19 drain_left.t2 a_n2982_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
R0 plus.n9 plus.t6 288.084
R1 plus.n43 plus.t12 288.084
R2 plus.n32 plus.t4 262.69
R3 plus.n30 plus.t19 262.69
R4 plus.n2 plus.t11 262.69
R5 plus.n24 plus.t0 262.69
R6 plus.n4 plus.t15 262.69
R7 plus.n18 plus.t5 262.69
R8 plus.n6 plus.t14 262.69
R9 plus.n12 plus.t2 262.69
R10 plus.n8 plus.t16 262.69
R11 plus.n66 plus.t8 262.69
R12 plus.n64 plus.t7 262.69
R13 plus.n36 plus.t10 262.69
R14 plus.n58 plus.t18 262.69
R15 plus.n38 plus.t17 262.69
R16 plus.n52 plus.t3 262.69
R17 plus.n40 plus.t1 262.69
R18 plus.n46 plus.t9 262.69
R19 plus.n42 plus.t13 262.69
R20 plus.n11 plus.n10 161.3
R21 plus.n12 plus.n7 161.3
R22 plus.n14 plus.n13 161.3
R23 plus.n15 plus.n6 161.3
R24 plus.n17 plus.n16 161.3
R25 plus.n18 plus.n5 161.3
R26 plus.n20 plus.n19 161.3
R27 plus.n21 plus.n4 161.3
R28 plus.n23 plus.n22 161.3
R29 plus.n24 plus.n3 161.3
R30 plus.n26 plus.n25 161.3
R31 plus.n27 plus.n2 161.3
R32 plus.n29 plus.n28 161.3
R33 plus.n30 plus.n1 161.3
R34 plus.n31 plus.n0 161.3
R35 plus.n33 plus.n32 161.3
R36 plus.n45 plus.n44 161.3
R37 plus.n46 plus.n41 161.3
R38 plus.n48 plus.n47 161.3
R39 plus.n49 plus.n40 161.3
R40 plus.n51 plus.n50 161.3
R41 plus.n52 plus.n39 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n55 plus.n38 161.3
R44 plus.n57 plus.n56 161.3
R45 plus.n58 plus.n37 161.3
R46 plus.n60 plus.n59 161.3
R47 plus.n61 plus.n36 161.3
R48 plus.n63 plus.n62 161.3
R49 plus.n64 plus.n35 161.3
R50 plus.n65 plus.n34 161.3
R51 plus.n67 plus.n66 161.3
R52 plus.n10 plus.n9 45.0031
R53 plus.n44 plus.n43 45.0031
R54 plus.n32 plus.n31 41.6278
R55 plus.n66 plus.n65 41.6278
R56 plus.n30 plus.n29 37.246
R57 plus.n11 plus.n8 37.246
R58 plus.n64 plus.n63 37.246
R59 plus.n45 plus.n42 37.246
R60 plus.n25 plus.n2 32.8641
R61 plus.n13 plus.n12 32.8641
R62 plus.n59 plus.n36 32.8641
R63 plus.n47 plus.n46 32.8641
R64 plus plus.n67 32.1922
R65 plus.n24 plus.n23 28.4823
R66 plus.n17 plus.n6 28.4823
R67 plus.n58 plus.n57 28.4823
R68 plus.n51 plus.n40 28.4823
R69 plus.n19 plus.n18 24.1005
R70 plus.n19 plus.n4 24.1005
R71 plus.n53 plus.n38 24.1005
R72 plus.n53 plus.n52 24.1005
R73 plus.n23 plus.n4 19.7187
R74 plus.n18 plus.n17 19.7187
R75 plus.n57 plus.n38 19.7187
R76 plus.n52 plus.n51 19.7187
R77 plus.n9 plus.n8 15.6319
R78 plus.n43 plus.n42 15.6319
R79 plus.n25 plus.n24 15.3369
R80 plus.n13 plus.n6 15.3369
R81 plus.n59 plus.n58 15.3369
R82 plus.n47 plus.n40 15.3369
R83 plus.n29 plus.n2 10.955
R84 plus.n12 plus.n11 10.955
R85 plus.n63 plus.n36 10.955
R86 plus.n46 plus.n45 10.955
R87 plus plus.n33 10.0384
R88 plus.n31 plus.n30 6.57323
R89 plus.n65 plus.n64 6.57323
R90 plus.n10 plus.n7 0.189894
R91 plus.n14 plus.n7 0.189894
R92 plus.n15 plus.n14 0.189894
R93 plus.n16 plus.n15 0.189894
R94 plus.n16 plus.n5 0.189894
R95 plus.n20 plus.n5 0.189894
R96 plus.n21 plus.n20 0.189894
R97 plus.n22 plus.n21 0.189894
R98 plus.n22 plus.n3 0.189894
R99 plus.n26 plus.n3 0.189894
R100 plus.n27 plus.n26 0.189894
R101 plus.n28 plus.n27 0.189894
R102 plus.n28 plus.n1 0.189894
R103 plus.n1 plus.n0 0.189894
R104 plus.n33 plus.n0 0.189894
R105 plus.n67 plus.n34 0.189894
R106 plus.n35 plus.n34 0.189894
R107 plus.n62 plus.n35 0.189894
R108 plus.n62 plus.n61 0.189894
R109 plus.n61 plus.n60 0.189894
R110 plus.n60 plus.n37 0.189894
R111 plus.n56 plus.n37 0.189894
R112 plus.n56 plus.n55 0.189894
R113 plus.n55 plus.n54 0.189894
R114 plus.n54 plus.n39 0.189894
R115 plus.n50 plus.n39 0.189894
R116 plus.n50 plus.n49 0.189894
R117 plus.n49 plus.n48 0.189894
R118 plus.n48 plus.n41 0.189894
R119 plus.n44 plus.n41 0.189894
R120 drain_left.n10 drain_left.n8 68.0787
R121 drain_left.n6 drain_left.n4 68.0786
R122 drain_left.n2 drain_left.n0 68.0786
R123 drain_left.n14 drain_left.n13 67.1908
R124 drain_left.n12 drain_left.n11 67.1908
R125 drain_left.n10 drain_left.n9 67.1908
R126 drain_left.n16 drain_left.n15 67.1907
R127 drain_left.n7 drain_left.n3 67.1907
R128 drain_left.n6 drain_left.n5 67.1907
R129 drain_left.n2 drain_left.n1 67.1907
R130 drain_left drain_left.n7 29.9251
R131 drain_left drain_left.n16 6.54115
R132 drain_left.n3 drain_left.t13 3.3005
R133 drain_left.n3 drain_left.t3 3.3005
R134 drain_left.n4 drain_left.t18 3.3005
R135 drain_left.n4 drain_left.t4 3.3005
R136 drain_left.n5 drain_left.t5 3.3005
R137 drain_left.n5 drain_left.t0 3.3005
R138 drain_left.n1 drain_left.t14 3.3005
R139 drain_left.n1 drain_left.t7 3.3005
R140 drain_left.n0 drain_left.t9 3.3005
R141 drain_left.n0 drain_left.t17 3.3005
R142 drain_left.n15 drain_left.t2 3.3005
R143 drain_left.n15 drain_left.t11 3.3005
R144 drain_left.n13 drain_left.t10 3.3005
R145 drain_left.n13 drain_left.t1 3.3005
R146 drain_left.n11 drain_left.t6 3.3005
R147 drain_left.n11 drain_left.t19 3.3005
R148 drain_left.n9 drain_left.t8 3.3005
R149 drain_left.n9 drain_left.t15 3.3005
R150 drain_left.n8 drain_left.t16 3.3005
R151 drain_left.n8 drain_left.t12 3.3005
R152 drain_left.n12 drain_left.n10 0.888431
R153 drain_left.n14 drain_left.n12 0.888431
R154 drain_left.n16 drain_left.n14 0.888431
R155 drain_left.n7 drain_left.n6 0.833085
R156 drain_left.n7 drain_left.n2 0.833085
R157 source.n282 source.n256 289.615
R158 source.n242 source.n216 289.615
R159 source.n210 source.n184 289.615
R160 source.n170 source.n144 289.615
R161 source.n26 source.n0 289.615
R162 source.n66 source.n40 289.615
R163 source.n98 source.n72 289.615
R164 source.n138 source.n112 289.615
R165 source.n267 source.n266 185
R166 source.n264 source.n263 185
R167 source.n273 source.n272 185
R168 source.n275 source.n274 185
R169 source.n260 source.n259 185
R170 source.n281 source.n280 185
R171 source.n283 source.n282 185
R172 source.n227 source.n226 185
R173 source.n224 source.n223 185
R174 source.n233 source.n232 185
R175 source.n235 source.n234 185
R176 source.n220 source.n219 185
R177 source.n241 source.n240 185
R178 source.n243 source.n242 185
R179 source.n195 source.n194 185
R180 source.n192 source.n191 185
R181 source.n201 source.n200 185
R182 source.n203 source.n202 185
R183 source.n188 source.n187 185
R184 source.n209 source.n208 185
R185 source.n211 source.n210 185
R186 source.n155 source.n154 185
R187 source.n152 source.n151 185
R188 source.n161 source.n160 185
R189 source.n163 source.n162 185
R190 source.n148 source.n147 185
R191 source.n169 source.n168 185
R192 source.n171 source.n170 185
R193 source.n27 source.n26 185
R194 source.n25 source.n24 185
R195 source.n4 source.n3 185
R196 source.n19 source.n18 185
R197 source.n17 source.n16 185
R198 source.n8 source.n7 185
R199 source.n11 source.n10 185
R200 source.n67 source.n66 185
R201 source.n65 source.n64 185
R202 source.n44 source.n43 185
R203 source.n59 source.n58 185
R204 source.n57 source.n56 185
R205 source.n48 source.n47 185
R206 source.n51 source.n50 185
R207 source.n99 source.n98 185
R208 source.n97 source.n96 185
R209 source.n76 source.n75 185
R210 source.n91 source.n90 185
R211 source.n89 source.n88 185
R212 source.n80 source.n79 185
R213 source.n83 source.n82 185
R214 source.n139 source.n138 185
R215 source.n137 source.n136 185
R216 source.n116 source.n115 185
R217 source.n131 source.n130 185
R218 source.n129 source.n128 185
R219 source.n120 source.n119 185
R220 source.n123 source.n122 185
R221 source.t4 source.n265 147.661
R222 source.t10 source.n225 147.661
R223 source.t27 source.n193 147.661
R224 source.t31 source.n153 147.661
R225 source.t35 source.n9 147.661
R226 source.t33 source.n49 147.661
R227 source.t6 source.n81 147.661
R228 source.t14 source.n121 147.661
R229 source.n266 source.n263 104.615
R230 source.n273 source.n263 104.615
R231 source.n274 source.n273 104.615
R232 source.n274 source.n259 104.615
R233 source.n281 source.n259 104.615
R234 source.n282 source.n281 104.615
R235 source.n226 source.n223 104.615
R236 source.n233 source.n223 104.615
R237 source.n234 source.n233 104.615
R238 source.n234 source.n219 104.615
R239 source.n241 source.n219 104.615
R240 source.n242 source.n241 104.615
R241 source.n194 source.n191 104.615
R242 source.n201 source.n191 104.615
R243 source.n202 source.n201 104.615
R244 source.n202 source.n187 104.615
R245 source.n209 source.n187 104.615
R246 source.n210 source.n209 104.615
R247 source.n154 source.n151 104.615
R248 source.n161 source.n151 104.615
R249 source.n162 source.n161 104.615
R250 source.n162 source.n147 104.615
R251 source.n169 source.n147 104.615
R252 source.n170 source.n169 104.615
R253 source.n26 source.n25 104.615
R254 source.n25 source.n3 104.615
R255 source.n18 source.n3 104.615
R256 source.n18 source.n17 104.615
R257 source.n17 source.n7 104.615
R258 source.n10 source.n7 104.615
R259 source.n66 source.n65 104.615
R260 source.n65 source.n43 104.615
R261 source.n58 source.n43 104.615
R262 source.n58 source.n57 104.615
R263 source.n57 source.n47 104.615
R264 source.n50 source.n47 104.615
R265 source.n98 source.n97 104.615
R266 source.n97 source.n75 104.615
R267 source.n90 source.n75 104.615
R268 source.n90 source.n89 104.615
R269 source.n89 source.n79 104.615
R270 source.n82 source.n79 104.615
R271 source.n138 source.n137 104.615
R272 source.n137 source.n115 104.615
R273 source.n130 source.n115 104.615
R274 source.n130 source.n129 104.615
R275 source.n129 source.n119 104.615
R276 source.n122 source.n119 104.615
R277 source.n266 source.t4 52.3082
R278 source.n226 source.t10 52.3082
R279 source.n194 source.t27 52.3082
R280 source.n154 source.t31 52.3082
R281 source.n10 source.t35 52.3082
R282 source.n50 source.t33 52.3082
R283 source.n82 source.t6 52.3082
R284 source.n122 source.t14 52.3082
R285 source.n33 source.n32 50.512
R286 source.n35 source.n34 50.512
R287 source.n37 source.n36 50.512
R288 source.n39 source.n38 50.512
R289 source.n105 source.n104 50.512
R290 source.n107 source.n106 50.512
R291 source.n109 source.n108 50.512
R292 source.n111 source.n110 50.512
R293 source.n255 source.n254 50.5119
R294 source.n253 source.n252 50.5119
R295 source.n251 source.n250 50.5119
R296 source.n249 source.n248 50.5119
R297 source.n183 source.n182 50.5119
R298 source.n181 source.n180 50.5119
R299 source.n179 source.n178 50.5119
R300 source.n177 source.n176 50.5119
R301 source.n287 source.n286 32.1853
R302 source.n247 source.n246 32.1853
R303 source.n215 source.n214 32.1853
R304 source.n175 source.n174 32.1853
R305 source.n31 source.n30 32.1853
R306 source.n71 source.n70 32.1853
R307 source.n103 source.n102 32.1853
R308 source.n143 source.n142 32.1853
R309 source.n175 source.n143 17.6302
R310 source.n267 source.n265 15.6674
R311 source.n227 source.n225 15.6674
R312 source.n195 source.n193 15.6674
R313 source.n155 source.n153 15.6674
R314 source.n11 source.n9 15.6674
R315 source.n51 source.n49 15.6674
R316 source.n83 source.n81 15.6674
R317 source.n123 source.n121 15.6674
R318 source.n268 source.n264 12.8005
R319 source.n228 source.n224 12.8005
R320 source.n196 source.n192 12.8005
R321 source.n156 source.n152 12.8005
R322 source.n12 source.n8 12.8005
R323 source.n52 source.n48 12.8005
R324 source.n84 source.n80 12.8005
R325 source.n124 source.n120 12.8005
R326 source.n272 source.n271 12.0247
R327 source.n232 source.n231 12.0247
R328 source.n200 source.n199 12.0247
R329 source.n160 source.n159 12.0247
R330 source.n16 source.n15 12.0247
R331 source.n56 source.n55 12.0247
R332 source.n88 source.n87 12.0247
R333 source.n128 source.n127 12.0247
R334 source.n288 source.n31 11.9233
R335 source.n275 source.n262 11.249
R336 source.n235 source.n222 11.249
R337 source.n203 source.n190 11.249
R338 source.n163 source.n150 11.249
R339 source.n19 source.n6 11.249
R340 source.n59 source.n46 11.249
R341 source.n91 source.n78 11.249
R342 source.n131 source.n118 11.249
R343 source.n276 source.n260 10.4732
R344 source.n236 source.n220 10.4732
R345 source.n204 source.n188 10.4732
R346 source.n164 source.n148 10.4732
R347 source.n20 source.n4 10.4732
R348 source.n60 source.n44 10.4732
R349 source.n92 source.n76 10.4732
R350 source.n132 source.n116 10.4732
R351 source.n280 source.n279 9.69747
R352 source.n240 source.n239 9.69747
R353 source.n208 source.n207 9.69747
R354 source.n168 source.n167 9.69747
R355 source.n24 source.n23 9.69747
R356 source.n64 source.n63 9.69747
R357 source.n96 source.n95 9.69747
R358 source.n136 source.n135 9.69747
R359 source.n286 source.n285 9.45567
R360 source.n246 source.n245 9.45567
R361 source.n214 source.n213 9.45567
R362 source.n174 source.n173 9.45567
R363 source.n30 source.n29 9.45567
R364 source.n70 source.n69 9.45567
R365 source.n102 source.n101 9.45567
R366 source.n142 source.n141 9.45567
R367 source.n285 source.n284 9.3005
R368 source.n258 source.n257 9.3005
R369 source.n279 source.n278 9.3005
R370 source.n277 source.n276 9.3005
R371 source.n262 source.n261 9.3005
R372 source.n271 source.n270 9.3005
R373 source.n269 source.n268 9.3005
R374 source.n245 source.n244 9.3005
R375 source.n218 source.n217 9.3005
R376 source.n239 source.n238 9.3005
R377 source.n237 source.n236 9.3005
R378 source.n222 source.n221 9.3005
R379 source.n231 source.n230 9.3005
R380 source.n229 source.n228 9.3005
R381 source.n213 source.n212 9.3005
R382 source.n186 source.n185 9.3005
R383 source.n207 source.n206 9.3005
R384 source.n205 source.n204 9.3005
R385 source.n190 source.n189 9.3005
R386 source.n199 source.n198 9.3005
R387 source.n197 source.n196 9.3005
R388 source.n173 source.n172 9.3005
R389 source.n146 source.n145 9.3005
R390 source.n167 source.n166 9.3005
R391 source.n165 source.n164 9.3005
R392 source.n150 source.n149 9.3005
R393 source.n159 source.n158 9.3005
R394 source.n157 source.n156 9.3005
R395 source.n29 source.n28 9.3005
R396 source.n2 source.n1 9.3005
R397 source.n23 source.n22 9.3005
R398 source.n21 source.n20 9.3005
R399 source.n6 source.n5 9.3005
R400 source.n15 source.n14 9.3005
R401 source.n13 source.n12 9.3005
R402 source.n69 source.n68 9.3005
R403 source.n42 source.n41 9.3005
R404 source.n63 source.n62 9.3005
R405 source.n61 source.n60 9.3005
R406 source.n46 source.n45 9.3005
R407 source.n55 source.n54 9.3005
R408 source.n53 source.n52 9.3005
R409 source.n101 source.n100 9.3005
R410 source.n74 source.n73 9.3005
R411 source.n95 source.n94 9.3005
R412 source.n93 source.n92 9.3005
R413 source.n78 source.n77 9.3005
R414 source.n87 source.n86 9.3005
R415 source.n85 source.n84 9.3005
R416 source.n141 source.n140 9.3005
R417 source.n114 source.n113 9.3005
R418 source.n135 source.n134 9.3005
R419 source.n133 source.n132 9.3005
R420 source.n118 source.n117 9.3005
R421 source.n127 source.n126 9.3005
R422 source.n125 source.n124 9.3005
R423 source.n283 source.n258 8.92171
R424 source.n243 source.n218 8.92171
R425 source.n211 source.n186 8.92171
R426 source.n171 source.n146 8.92171
R427 source.n27 source.n2 8.92171
R428 source.n67 source.n42 8.92171
R429 source.n99 source.n74 8.92171
R430 source.n139 source.n114 8.92171
R431 source.n284 source.n256 8.14595
R432 source.n244 source.n216 8.14595
R433 source.n212 source.n184 8.14595
R434 source.n172 source.n144 8.14595
R435 source.n28 source.n0 8.14595
R436 source.n68 source.n40 8.14595
R437 source.n100 source.n72 8.14595
R438 source.n140 source.n112 8.14595
R439 source.n286 source.n256 5.81868
R440 source.n246 source.n216 5.81868
R441 source.n214 source.n184 5.81868
R442 source.n174 source.n144 5.81868
R443 source.n30 source.n0 5.81868
R444 source.n70 source.n40 5.81868
R445 source.n102 source.n72 5.81868
R446 source.n142 source.n112 5.81868
R447 source.n288 source.n287 5.7074
R448 source.n284 source.n283 5.04292
R449 source.n244 source.n243 5.04292
R450 source.n212 source.n211 5.04292
R451 source.n172 source.n171 5.04292
R452 source.n28 source.n27 5.04292
R453 source.n68 source.n67 5.04292
R454 source.n100 source.n99 5.04292
R455 source.n140 source.n139 5.04292
R456 source.n269 source.n265 4.38594
R457 source.n229 source.n225 4.38594
R458 source.n197 source.n193 4.38594
R459 source.n157 source.n153 4.38594
R460 source.n13 source.n9 4.38594
R461 source.n53 source.n49 4.38594
R462 source.n85 source.n81 4.38594
R463 source.n125 source.n121 4.38594
R464 source.n280 source.n258 4.26717
R465 source.n240 source.n218 4.26717
R466 source.n208 source.n186 4.26717
R467 source.n168 source.n146 4.26717
R468 source.n24 source.n2 4.26717
R469 source.n64 source.n42 4.26717
R470 source.n96 source.n74 4.26717
R471 source.n136 source.n114 4.26717
R472 source.n279 source.n260 3.49141
R473 source.n239 source.n220 3.49141
R474 source.n207 source.n188 3.49141
R475 source.n167 source.n148 3.49141
R476 source.n23 source.n4 3.49141
R477 source.n63 source.n44 3.49141
R478 source.n95 source.n76 3.49141
R479 source.n135 source.n116 3.49141
R480 source.n254 source.t2 3.3005
R481 source.n254 source.t1 3.3005
R482 source.n252 source.t8 3.3005
R483 source.n252 source.t19 3.3005
R484 source.n250 source.t17 3.3005
R485 source.n250 source.t16 3.3005
R486 source.n248 source.t12 3.3005
R487 source.n248 source.t15 3.3005
R488 source.n182 source.t30 3.3005
R489 source.n182 source.t26 3.3005
R490 source.n180 source.t36 3.3005
R491 source.n180 source.t38 3.3005
R492 source.n178 source.t21 3.3005
R493 source.n178 source.t22 3.3005
R494 source.n176 source.t32 3.3005
R495 source.n176 source.t29 3.3005
R496 source.n32 source.t28 3.3005
R497 source.n32 source.t20 3.3005
R498 source.n34 source.t24 3.3005
R499 source.n34 source.t39 3.3005
R500 source.n36 source.t25 3.3005
R501 source.n36 source.t34 3.3005
R502 source.n38 source.t23 3.3005
R503 source.n38 source.t37 3.3005
R504 source.n104 source.t9 3.3005
R505 source.n104 source.t5 3.3005
R506 source.n106 source.t18 3.3005
R507 source.n106 source.t0 3.3005
R508 source.n108 source.t13 3.3005
R509 source.n108 source.t11 3.3005
R510 source.n110 source.t7 3.3005
R511 source.n110 source.t3 3.3005
R512 source.n276 source.n275 2.71565
R513 source.n236 source.n235 2.71565
R514 source.n204 source.n203 2.71565
R515 source.n164 source.n163 2.71565
R516 source.n20 source.n19 2.71565
R517 source.n60 source.n59 2.71565
R518 source.n92 source.n91 2.71565
R519 source.n132 source.n131 2.71565
R520 source.n272 source.n262 1.93989
R521 source.n232 source.n222 1.93989
R522 source.n200 source.n190 1.93989
R523 source.n160 source.n150 1.93989
R524 source.n16 source.n6 1.93989
R525 source.n56 source.n46 1.93989
R526 source.n88 source.n78 1.93989
R527 source.n128 source.n118 1.93989
R528 source.n271 source.n264 1.16414
R529 source.n231 source.n224 1.16414
R530 source.n199 source.n192 1.16414
R531 source.n159 source.n152 1.16414
R532 source.n15 source.n8 1.16414
R533 source.n55 source.n48 1.16414
R534 source.n87 source.n80 1.16414
R535 source.n127 source.n120 1.16414
R536 source.n143 source.n111 0.888431
R537 source.n111 source.n109 0.888431
R538 source.n109 source.n107 0.888431
R539 source.n107 source.n105 0.888431
R540 source.n105 source.n103 0.888431
R541 source.n71 source.n39 0.888431
R542 source.n39 source.n37 0.888431
R543 source.n37 source.n35 0.888431
R544 source.n35 source.n33 0.888431
R545 source.n33 source.n31 0.888431
R546 source.n177 source.n175 0.888431
R547 source.n179 source.n177 0.888431
R548 source.n181 source.n179 0.888431
R549 source.n183 source.n181 0.888431
R550 source.n215 source.n183 0.888431
R551 source.n249 source.n247 0.888431
R552 source.n251 source.n249 0.888431
R553 source.n253 source.n251 0.888431
R554 source.n255 source.n253 0.888431
R555 source.n287 source.n255 0.888431
R556 source.n103 source.n71 0.470328
R557 source.n247 source.n215 0.470328
R558 source.n268 source.n267 0.388379
R559 source.n228 source.n227 0.388379
R560 source.n196 source.n195 0.388379
R561 source.n156 source.n155 0.388379
R562 source.n12 source.n11 0.388379
R563 source.n52 source.n51 0.388379
R564 source.n84 source.n83 0.388379
R565 source.n124 source.n123 0.388379
R566 source source.n288 0.188
R567 source.n270 source.n269 0.155672
R568 source.n270 source.n261 0.155672
R569 source.n277 source.n261 0.155672
R570 source.n278 source.n277 0.155672
R571 source.n278 source.n257 0.155672
R572 source.n285 source.n257 0.155672
R573 source.n230 source.n229 0.155672
R574 source.n230 source.n221 0.155672
R575 source.n237 source.n221 0.155672
R576 source.n238 source.n237 0.155672
R577 source.n238 source.n217 0.155672
R578 source.n245 source.n217 0.155672
R579 source.n198 source.n197 0.155672
R580 source.n198 source.n189 0.155672
R581 source.n205 source.n189 0.155672
R582 source.n206 source.n205 0.155672
R583 source.n206 source.n185 0.155672
R584 source.n213 source.n185 0.155672
R585 source.n158 source.n157 0.155672
R586 source.n158 source.n149 0.155672
R587 source.n165 source.n149 0.155672
R588 source.n166 source.n165 0.155672
R589 source.n166 source.n145 0.155672
R590 source.n173 source.n145 0.155672
R591 source.n29 source.n1 0.155672
R592 source.n22 source.n1 0.155672
R593 source.n22 source.n21 0.155672
R594 source.n21 source.n5 0.155672
R595 source.n14 source.n5 0.155672
R596 source.n14 source.n13 0.155672
R597 source.n69 source.n41 0.155672
R598 source.n62 source.n41 0.155672
R599 source.n62 source.n61 0.155672
R600 source.n61 source.n45 0.155672
R601 source.n54 source.n45 0.155672
R602 source.n54 source.n53 0.155672
R603 source.n101 source.n73 0.155672
R604 source.n94 source.n73 0.155672
R605 source.n94 source.n93 0.155672
R606 source.n93 source.n77 0.155672
R607 source.n86 source.n77 0.155672
R608 source.n86 source.n85 0.155672
R609 source.n141 source.n113 0.155672
R610 source.n134 source.n113 0.155672
R611 source.n134 source.n133 0.155672
R612 source.n133 source.n117 0.155672
R613 source.n126 source.n117 0.155672
R614 source.n126 source.n125 0.155672
R615 minus.n9 minus.t11 288.084
R616 minus.n43 minus.t13 288.084
R617 minus.n8 minus.t0 262.69
R618 minus.n12 minus.t8 262.69
R619 minus.n14 minus.t18 262.69
R620 minus.n18 minus.t6 262.69
R621 minus.n20 minus.t19 262.69
R622 minus.n24 minus.t4 262.69
R623 minus.n26 minus.t16 262.69
R624 minus.n30 minus.t3 262.69
R625 minus.n32 minus.t14 262.69
R626 minus.n42 minus.t15 262.69
R627 minus.n46 minus.t9 262.69
R628 minus.n48 minus.t10 262.69
R629 minus.n52 minus.t12 262.69
R630 minus.n54 minus.t5 262.69
R631 minus.n58 minus.t7 262.69
R632 minus.n60 minus.t2 262.69
R633 minus.n64 minus.t1 262.69
R634 minus.n66 minus.t17 262.69
R635 minus.n33 minus.n32 161.3
R636 minus.n31 minus.n0 161.3
R637 minus.n30 minus.n29 161.3
R638 minus.n28 minus.n1 161.3
R639 minus.n27 minus.n26 161.3
R640 minus.n25 minus.n2 161.3
R641 minus.n24 minus.n23 161.3
R642 minus.n22 minus.n3 161.3
R643 minus.n21 minus.n20 161.3
R644 minus.n19 minus.n4 161.3
R645 minus.n18 minus.n17 161.3
R646 minus.n16 minus.n5 161.3
R647 minus.n15 minus.n14 161.3
R648 minus.n13 minus.n6 161.3
R649 minus.n12 minus.n11 161.3
R650 minus.n10 minus.n7 161.3
R651 minus.n67 minus.n66 161.3
R652 minus.n65 minus.n34 161.3
R653 minus.n64 minus.n63 161.3
R654 minus.n62 minus.n35 161.3
R655 minus.n61 minus.n60 161.3
R656 minus.n59 minus.n36 161.3
R657 minus.n58 minus.n57 161.3
R658 minus.n56 minus.n37 161.3
R659 minus.n55 minus.n54 161.3
R660 minus.n53 minus.n38 161.3
R661 minus.n52 minus.n51 161.3
R662 minus.n50 minus.n39 161.3
R663 minus.n49 minus.n48 161.3
R664 minus.n47 minus.n40 161.3
R665 minus.n46 minus.n45 161.3
R666 minus.n44 minus.n41 161.3
R667 minus.n10 minus.n9 45.0031
R668 minus.n44 minus.n43 45.0031
R669 minus.n32 minus.n31 41.6278
R670 minus.n66 minus.n65 41.6278
R671 minus.n8 minus.n7 37.246
R672 minus.n30 minus.n1 37.246
R673 minus.n42 minus.n41 37.246
R674 minus.n64 minus.n35 37.246
R675 minus.n68 minus.n33 36.0384
R676 minus.n13 minus.n12 32.8641
R677 minus.n26 minus.n25 32.8641
R678 minus.n47 minus.n46 32.8641
R679 minus.n60 minus.n59 32.8641
R680 minus.n14 minus.n5 28.4823
R681 minus.n24 minus.n3 28.4823
R682 minus.n48 minus.n39 28.4823
R683 minus.n58 minus.n37 28.4823
R684 minus.n20 minus.n19 24.1005
R685 minus.n19 minus.n18 24.1005
R686 minus.n53 minus.n52 24.1005
R687 minus.n54 minus.n53 24.1005
R688 minus.n18 minus.n5 19.7187
R689 minus.n20 minus.n3 19.7187
R690 minus.n52 minus.n39 19.7187
R691 minus.n54 minus.n37 19.7187
R692 minus.n9 minus.n8 15.6319
R693 minus.n43 minus.n42 15.6319
R694 minus.n14 minus.n13 15.3369
R695 minus.n25 minus.n24 15.3369
R696 minus.n48 minus.n47 15.3369
R697 minus.n59 minus.n58 15.3369
R698 minus.n12 minus.n7 10.955
R699 minus.n26 minus.n1 10.955
R700 minus.n46 minus.n41 10.955
R701 minus.n60 minus.n35 10.955
R702 minus.n68 minus.n67 6.66717
R703 minus.n31 minus.n30 6.57323
R704 minus.n65 minus.n64 6.57323
R705 minus.n33 minus.n0 0.189894
R706 minus.n29 minus.n0 0.189894
R707 minus.n29 minus.n28 0.189894
R708 minus.n28 minus.n27 0.189894
R709 minus.n27 minus.n2 0.189894
R710 minus.n23 minus.n2 0.189894
R711 minus.n23 minus.n22 0.189894
R712 minus.n22 minus.n21 0.189894
R713 minus.n21 minus.n4 0.189894
R714 minus.n17 minus.n4 0.189894
R715 minus.n17 minus.n16 0.189894
R716 minus.n16 minus.n15 0.189894
R717 minus.n15 minus.n6 0.189894
R718 minus.n11 minus.n6 0.189894
R719 minus.n11 minus.n10 0.189894
R720 minus.n45 minus.n44 0.189894
R721 minus.n45 minus.n40 0.189894
R722 minus.n49 minus.n40 0.189894
R723 minus.n50 minus.n49 0.189894
R724 minus.n51 minus.n50 0.189894
R725 minus.n51 minus.n38 0.189894
R726 minus.n55 minus.n38 0.189894
R727 minus.n56 minus.n55 0.189894
R728 minus.n57 minus.n56 0.189894
R729 minus.n57 minus.n36 0.189894
R730 minus.n61 minus.n36 0.189894
R731 minus.n62 minus.n61 0.189894
R732 minus.n63 minus.n62 0.189894
R733 minus.n63 minus.n34 0.189894
R734 minus.n67 minus.n34 0.189894
R735 minus minus.n68 0.188
R736 drain_right.n10 drain_right.n8 68.0786
R737 drain_right.n6 drain_right.n4 68.0786
R738 drain_right.n2 drain_right.n0 68.0786
R739 drain_right.n10 drain_right.n9 67.1908
R740 drain_right.n12 drain_right.n11 67.1908
R741 drain_right.n14 drain_right.n13 67.1908
R742 drain_right.n16 drain_right.n15 67.1908
R743 drain_right.n7 drain_right.n3 67.1907
R744 drain_right.n6 drain_right.n5 67.1907
R745 drain_right.n2 drain_right.n1 67.1907
R746 drain_right drain_right.n7 29.3718
R747 drain_right drain_right.n16 6.54115
R748 drain_right.n3 drain_right.t7 3.3005
R749 drain_right.n3 drain_right.t14 3.3005
R750 drain_right.n4 drain_right.t18 3.3005
R751 drain_right.n4 drain_right.t2 3.3005
R752 drain_right.n5 drain_right.t12 3.3005
R753 drain_right.n5 drain_right.t17 3.3005
R754 drain_right.n1 drain_right.t10 3.3005
R755 drain_right.n1 drain_right.t9 3.3005
R756 drain_right.n0 drain_right.t6 3.3005
R757 drain_right.n0 drain_right.t4 3.3005
R758 drain_right.n8 drain_right.t19 3.3005
R759 drain_right.n8 drain_right.t8 3.3005
R760 drain_right.n9 drain_right.t1 3.3005
R761 drain_right.n9 drain_right.t11 3.3005
R762 drain_right.n11 drain_right.t0 3.3005
R763 drain_right.n11 drain_right.t13 3.3005
R764 drain_right.n13 drain_right.t3 3.3005
R765 drain_right.n13 drain_right.t15 3.3005
R766 drain_right.n15 drain_right.t5 3.3005
R767 drain_right.n15 drain_right.t16 3.3005
R768 drain_right.n16 drain_right.n14 0.888431
R769 drain_right.n14 drain_right.n12 0.888431
R770 drain_right.n12 drain_right.n10 0.888431
R771 drain_right.n7 drain_right.n6 0.833085
R772 drain_right.n7 drain_right.n2 0.833085
C0 source drain_right 14.088799f
C1 plus drain_right 0.454687f
C2 minus drain_right 6.64334f
C3 drain_right drain_left 1.59885f
C4 source plus 7.16192f
C5 source minus 7.1479f
C6 source drain_left 14.0865f
C7 minus plus 5.75442f
C8 plus drain_left 6.94088f
C9 minus drain_left 0.173554f
C10 drain_right a_n2982_n2088# 6.19181f
C11 drain_left a_n2982_n2088# 6.61692f
C12 source a_n2982_n2088# 5.811326f
C13 minus a_n2982_n2088# 11.466448f
C14 plus a_n2982_n2088# 13.01572f
C15 drain_right.t6 a_n2982_n2088# 0.128092f
C16 drain_right.t4 a_n2982_n2088# 0.128092f
C17 drain_right.n0 a_n2982_n2088# 1.0733f
C18 drain_right.t10 a_n2982_n2088# 0.128092f
C19 drain_right.t9 a_n2982_n2088# 0.128092f
C20 drain_right.n1 a_n2982_n2088# 1.06829f
C21 drain_right.n2 a_n2982_n2088# 0.749516f
C22 drain_right.t7 a_n2982_n2088# 0.128092f
C23 drain_right.t14 a_n2982_n2088# 0.128092f
C24 drain_right.n3 a_n2982_n2088# 1.06829f
C25 drain_right.t18 a_n2982_n2088# 0.128092f
C26 drain_right.t2 a_n2982_n2088# 0.128092f
C27 drain_right.n4 a_n2982_n2088# 1.0733f
C28 drain_right.t12 a_n2982_n2088# 0.128092f
C29 drain_right.t17 a_n2982_n2088# 0.128092f
C30 drain_right.n5 a_n2982_n2088# 1.06829f
C31 drain_right.n6 a_n2982_n2088# 0.749516f
C32 drain_right.n7 a_n2982_n2088# 1.55396f
C33 drain_right.t19 a_n2982_n2088# 0.128092f
C34 drain_right.t8 a_n2982_n2088# 0.128092f
C35 drain_right.n8 a_n2982_n2088# 1.0733f
C36 drain_right.t1 a_n2982_n2088# 0.128092f
C37 drain_right.t11 a_n2982_n2088# 0.128092f
C38 drain_right.n9 a_n2982_n2088# 1.06829f
C39 drain_right.n10 a_n2982_n2088# 0.753576f
C40 drain_right.t0 a_n2982_n2088# 0.128092f
C41 drain_right.t13 a_n2982_n2088# 0.128092f
C42 drain_right.n11 a_n2982_n2088# 1.06829f
C43 drain_right.n12 a_n2982_n2088# 0.373854f
C44 drain_right.t3 a_n2982_n2088# 0.128092f
C45 drain_right.t15 a_n2982_n2088# 0.128092f
C46 drain_right.n13 a_n2982_n2088# 1.06829f
C47 drain_right.n14 a_n2982_n2088# 0.373854f
C48 drain_right.t5 a_n2982_n2088# 0.128092f
C49 drain_right.t16 a_n2982_n2088# 0.128092f
C50 drain_right.n15 a_n2982_n2088# 1.06829f
C51 drain_right.n16 a_n2982_n2088# 0.61281f
C52 minus.n0 a_n2982_n2088# 0.040426f
C53 minus.n1 a_n2982_n2088# 0.009173f
C54 minus.t3 a_n2982_n2088# 0.492482f
C55 minus.n2 a_n2982_n2088# 0.040426f
C56 minus.n3 a_n2982_n2088# 0.009173f
C57 minus.t4 a_n2982_n2088# 0.492482f
C58 minus.n4 a_n2982_n2088# 0.040426f
C59 minus.n5 a_n2982_n2088# 0.009173f
C60 minus.t6 a_n2982_n2088# 0.492482f
C61 minus.n6 a_n2982_n2088# 0.040426f
C62 minus.n7 a_n2982_n2088# 0.009173f
C63 minus.t8 a_n2982_n2088# 0.492482f
C64 minus.t11 a_n2982_n2088# 0.512578f
C65 minus.t0 a_n2982_n2088# 0.492482f
C66 minus.n8 a_n2982_n2088# 0.234333f
C67 minus.n9 a_n2982_n2088# 0.210377f
C68 minus.n10 a_n2982_n2088# 0.172554f
C69 minus.n11 a_n2982_n2088# 0.040426f
C70 minus.n12 a_n2982_n2088# 0.227571f
C71 minus.n13 a_n2982_n2088# 0.009173f
C72 minus.t18 a_n2982_n2088# 0.492482f
C73 minus.n14 a_n2982_n2088# 0.227571f
C74 minus.n15 a_n2982_n2088# 0.040426f
C75 minus.n16 a_n2982_n2088# 0.040426f
C76 minus.n17 a_n2982_n2088# 0.040426f
C77 minus.n18 a_n2982_n2088# 0.227571f
C78 minus.n19 a_n2982_n2088# 0.009173f
C79 minus.t19 a_n2982_n2088# 0.492482f
C80 minus.n20 a_n2982_n2088# 0.227571f
C81 minus.n21 a_n2982_n2088# 0.040426f
C82 minus.n22 a_n2982_n2088# 0.040426f
C83 minus.n23 a_n2982_n2088# 0.040426f
C84 minus.n24 a_n2982_n2088# 0.227571f
C85 minus.n25 a_n2982_n2088# 0.009173f
C86 minus.t16 a_n2982_n2088# 0.492482f
C87 minus.n26 a_n2982_n2088# 0.227571f
C88 minus.n27 a_n2982_n2088# 0.040426f
C89 minus.n28 a_n2982_n2088# 0.040426f
C90 minus.n29 a_n2982_n2088# 0.040426f
C91 minus.n30 a_n2982_n2088# 0.227571f
C92 minus.n31 a_n2982_n2088# 0.009173f
C93 minus.t14 a_n2982_n2088# 0.492482f
C94 minus.n32 a_n2982_n2088# 0.227197f
C95 minus.n33 a_n2982_n2088# 1.42434f
C96 minus.n34 a_n2982_n2088# 0.040426f
C97 minus.n35 a_n2982_n2088# 0.009173f
C98 minus.n36 a_n2982_n2088# 0.040426f
C99 minus.n37 a_n2982_n2088# 0.009173f
C100 minus.n38 a_n2982_n2088# 0.040426f
C101 minus.n39 a_n2982_n2088# 0.009173f
C102 minus.n40 a_n2982_n2088# 0.040426f
C103 minus.n41 a_n2982_n2088# 0.009173f
C104 minus.t13 a_n2982_n2088# 0.512578f
C105 minus.t15 a_n2982_n2088# 0.492482f
C106 minus.n42 a_n2982_n2088# 0.234333f
C107 minus.n43 a_n2982_n2088# 0.210377f
C108 minus.n44 a_n2982_n2088# 0.172554f
C109 minus.n45 a_n2982_n2088# 0.040426f
C110 minus.t9 a_n2982_n2088# 0.492482f
C111 minus.n46 a_n2982_n2088# 0.227571f
C112 minus.n47 a_n2982_n2088# 0.009173f
C113 minus.t10 a_n2982_n2088# 0.492482f
C114 minus.n48 a_n2982_n2088# 0.227571f
C115 minus.n49 a_n2982_n2088# 0.040426f
C116 minus.n50 a_n2982_n2088# 0.040426f
C117 minus.n51 a_n2982_n2088# 0.040426f
C118 minus.t12 a_n2982_n2088# 0.492482f
C119 minus.n52 a_n2982_n2088# 0.227571f
C120 minus.n53 a_n2982_n2088# 0.009173f
C121 minus.t5 a_n2982_n2088# 0.492482f
C122 minus.n54 a_n2982_n2088# 0.227571f
C123 minus.n55 a_n2982_n2088# 0.040426f
C124 minus.n56 a_n2982_n2088# 0.040426f
C125 minus.n57 a_n2982_n2088# 0.040426f
C126 minus.t7 a_n2982_n2088# 0.492482f
C127 minus.n58 a_n2982_n2088# 0.227571f
C128 minus.n59 a_n2982_n2088# 0.009173f
C129 minus.t2 a_n2982_n2088# 0.492482f
C130 minus.n60 a_n2982_n2088# 0.227571f
C131 minus.n61 a_n2982_n2088# 0.040426f
C132 minus.n62 a_n2982_n2088# 0.040426f
C133 minus.n63 a_n2982_n2088# 0.040426f
C134 minus.t1 a_n2982_n2088# 0.492482f
C135 minus.n64 a_n2982_n2088# 0.227571f
C136 minus.n65 a_n2982_n2088# 0.009173f
C137 minus.t17 a_n2982_n2088# 0.492482f
C138 minus.n66 a_n2982_n2088# 0.227197f
C139 minus.n67 a_n2982_n2088# 0.280092f
C140 minus.n68 a_n2982_n2088# 1.72556f
C141 source.n0 a_n2982_n2088# 0.036611f
C142 source.n1 a_n2982_n2088# 0.026047f
C143 source.n2 a_n2982_n2088# 0.013996f
C144 source.n3 a_n2982_n2088# 0.033082f
C145 source.n4 a_n2982_n2088# 0.01482f
C146 source.n5 a_n2982_n2088# 0.026047f
C147 source.n6 a_n2982_n2088# 0.013996f
C148 source.n7 a_n2982_n2088# 0.033082f
C149 source.n8 a_n2982_n2088# 0.01482f
C150 source.n9 a_n2982_n2088# 0.111461f
C151 source.t35 a_n2982_n2088# 0.05392f
C152 source.n10 a_n2982_n2088# 0.024812f
C153 source.n11 a_n2982_n2088# 0.019541f
C154 source.n12 a_n2982_n2088# 0.013996f
C155 source.n13 a_n2982_n2088# 0.619755f
C156 source.n14 a_n2982_n2088# 0.026047f
C157 source.n15 a_n2982_n2088# 0.013996f
C158 source.n16 a_n2982_n2088# 0.01482f
C159 source.n17 a_n2982_n2088# 0.033082f
C160 source.n18 a_n2982_n2088# 0.033082f
C161 source.n19 a_n2982_n2088# 0.01482f
C162 source.n20 a_n2982_n2088# 0.013996f
C163 source.n21 a_n2982_n2088# 0.026047f
C164 source.n22 a_n2982_n2088# 0.026047f
C165 source.n23 a_n2982_n2088# 0.013996f
C166 source.n24 a_n2982_n2088# 0.01482f
C167 source.n25 a_n2982_n2088# 0.033082f
C168 source.n26 a_n2982_n2088# 0.071617f
C169 source.n27 a_n2982_n2088# 0.01482f
C170 source.n28 a_n2982_n2088# 0.013996f
C171 source.n29 a_n2982_n2088# 0.060206f
C172 source.n30 a_n2982_n2088# 0.040073f
C173 source.n31 a_n2982_n2088# 0.680432f
C174 source.t28 a_n2982_n2088# 0.123497f
C175 source.t20 a_n2982_n2088# 0.123497f
C176 source.n32 a_n2982_n2088# 0.961806f
C177 source.n33 a_n2982_n2088# 0.393207f
C178 source.t24 a_n2982_n2088# 0.123497f
C179 source.t39 a_n2982_n2088# 0.123497f
C180 source.n34 a_n2982_n2088# 0.961806f
C181 source.n35 a_n2982_n2088# 0.393207f
C182 source.t25 a_n2982_n2088# 0.123497f
C183 source.t34 a_n2982_n2088# 0.123497f
C184 source.n36 a_n2982_n2088# 0.961806f
C185 source.n37 a_n2982_n2088# 0.393207f
C186 source.t23 a_n2982_n2088# 0.123497f
C187 source.t37 a_n2982_n2088# 0.123497f
C188 source.n38 a_n2982_n2088# 0.961806f
C189 source.n39 a_n2982_n2088# 0.393207f
C190 source.n40 a_n2982_n2088# 0.036611f
C191 source.n41 a_n2982_n2088# 0.026047f
C192 source.n42 a_n2982_n2088# 0.013996f
C193 source.n43 a_n2982_n2088# 0.033082f
C194 source.n44 a_n2982_n2088# 0.01482f
C195 source.n45 a_n2982_n2088# 0.026047f
C196 source.n46 a_n2982_n2088# 0.013996f
C197 source.n47 a_n2982_n2088# 0.033082f
C198 source.n48 a_n2982_n2088# 0.01482f
C199 source.n49 a_n2982_n2088# 0.111461f
C200 source.t33 a_n2982_n2088# 0.05392f
C201 source.n50 a_n2982_n2088# 0.024812f
C202 source.n51 a_n2982_n2088# 0.019541f
C203 source.n52 a_n2982_n2088# 0.013996f
C204 source.n53 a_n2982_n2088# 0.619755f
C205 source.n54 a_n2982_n2088# 0.026047f
C206 source.n55 a_n2982_n2088# 0.013996f
C207 source.n56 a_n2982_n2088# 0.01482f
C208 source.n57 a_n2982_n2088# 0.033082f
C209 source.n58 a_n2982_n2088# 0.033082f
C210 source.n59 a_n2982_n2088# 0.01482f
C211 source.n60 a_n2982_n2088# 0.013996f
C212 source.n61 a_n2982_n2088# 0.026047f
C213 source.n62 a_n2982_n2088# 0.026047f
C214 source.n63 a_n2982_n2088# 0.013996f
C215 source.n64 a_n2982_n2088# 0.01482f
C216 source.n65 a_n2982_n2088# 0.033082f
C217 source.n66 a_n2982_n2088# 0.071617f
C218 source.n67 a_n2982_n2088# 0.01482f
C219 source.n68 a_n2982_n2088# 0.013996f
C220 source.n69 a_n2982_n2088# 0.060206f
C221 source.n70 a_n2982_n2088# 0.040073f
C222 source.n71 a_n2982_n2088# 0.1362f
C223 source.n72 a_n2982_n2088# 0.036611f
C224 source.n73 a_n2982_n2088# 0.026047f
C225 source.n74 a_n2982_n2088# 0.013996f
C226 source.n75 a_n2982_n2088# 0.033082f
C227 source.n76 a_n2982_n2088# 0.01482f
C228 source.n77 a_n2982_n2088# 0.026047f
C229 source.n78 a_n2982_n2088# 0.013996f
C230 source.n79 a_n2982_n2088# 0.033082f
C231 source.n80 a_n2982_n2088# 0.01482f
C232 source.n81 a_n2982_n2088# 0.111461f
C233 source.t6 a_n2982_n2088# 0.05392f
C234 source.n82 a_n2982_n2088# 0.024812f
C235 source.n83 a_n2982_n2088# 0.019541f
C236 source.n84 a_n2982_n2088# 0.013996f
C237 source.n85 a_n2982_n2088# 0.619755f
C238 source.n86 a_n2982_n2088# 0.026047f
C239 source.n87 a_n2982_n2088# 0.013996f
C240 source.n88 a_n2982_n2088# 0.01482f
C241 source.n89 a_n2982_n2088# 0.033082f
C242 source.n90 a_n2982_n2088# 0.033082f
C243 source.n91 a_n2982_n2088# 0.01482f
C244 source.n92 a_n2982_n2088# 0.013996f
C245 source.n93 a_n2982_n2088# 0.026047f
C246 source.n94 a_n2982_n2088# 0.026047f
C247 source.n95 a_n2982_n2088# 0.013996f
C248 source.n96 a_n2982_n2088# 0.01482f
C249 source.n97 a_n2982_n2088# 0.033082f
C250 source.n98 a_n2982_n2088# 0.071617f
C251 source.n99 a_n2982_n2088# 0.01482f
C252 source.n100 a_n2982_n2088# 0.013996f
C253 source.n101 a_n2982_n2088# 0.060206f
C254 source.n102 a_n2982_n2088# 0.040073f
C255 source.n103 a_n2982_n2088# 0.1362f
C256 source.t9 a_n2982_n2088# 0.123497f
C257 source.t5 a_n2982_n2088# 0.123497f
C258 source.n104 a_n2982_n2088# 0.961806f
C259 source.n105 a_n2982_n2088# 0.393207f
C260 source.t18 a_n2982_n2088# 0.123497f
C261 source.t0 a_n2982_n2088# 0.123497f
C262 source.n106 a_n2982_n2088# 0.961806f
C263 source.n107 a_n2982_n2088# 0.393207f
C264 source.t13 a_n2982_n2088# 0.123497f
C265 source.t11 a_n2982_n2088# 0.123497f
C266 source.n108 a_n2982_n2088# 0.961806f
C267 source.n109 a_n2982_n2088# 0.393207f
C268 source.t7 a_n2982_n2088# 0.123497f
C269 source.t3 a_n2982_n2088# 0.123497f
C270 source.n110 a_n2982_n2088# 0.961806f
C271 source.n111 a_n2982_n2088# 0.393207f
C272 source.n112 a_n2982_n2088# 0.036611f
C273 source.n113 a_n2982_n2088# 0.026047f
C274 source.n114 a_n2982_n2088# 0.013996f
C275 source.n115 a_n2982_n2088# 0.033082f
C276 source.n116 a_n2982_n2088# 0.01482f
C277 source.n117 a_n2982_n2088# 0.026047f
C278 source.n118 a_n2982_n2088# 0.013996f
C279 source.n119 a_n2982_n2088# 0.033082f
C280 source.n120 a_n2982_n2088# 0.01482f
C281 source.n121 a_n2982_n2088# 0.111461f
C282 source.t14 a_n2982_n2088# 0.05392f
C283 source.n122 a_n2982_n2088# 0.024812f
C284 source.n123 a_n2982_n2088# 0.019541f
C285 source.n124 a_n2982_n2088# 0.013996f
C286 source.n125 a_n2982_n2088# 0.619755f
C287 source.n126 a_n2982_n2088# 0.026047f
C288 source.n127 a_n2982_n2088# 0.013996f
C289 source.n128 a_n2982_n2088# 0.01482f
C290 source.n129 a_n2982_n2088# 0.033082f
C291 source.n130 a_n2982_n2088# 0.033082f
C292 source.n131 a_n2982_n2088# 0.01482f
C293 source.n132 a_n2982_n2088# 0.013996f
C294 source.n133 a_n2982_n2088# 0.026047f
C295 source.n134 a_n2982_n2088# 0.026047f
C296 source.n135 a_n2982_n2088# 0.013996f
C297 source.n136 a_n2982_n2088# 0.01482f
C298 source.n137 a_n2982_n2088# 0.033082f
C299 source.n138 a_n2982_n2088# 0.071617f
C300 source.n139 a_n2982_n2088# 0.01482f
C301 source.n140 a_n2982_n2088# 0.013996f
C302 source.n141 a_n2982_n2088# 0.060206f
C303 source.n142 a_n2982_n2088# 0.040073f
C304 source.n143 a_n2982_n2088# 1.02411f
C305 source.n144 a_n2982_n2088# 0.036611f
C306 source.n145 a_n2982_n2088# 0.026047f
C307 source.n146 a_n2982_n2088# 0.013996f
C308 source.n147 a_n2982_n2088# 0.033082f
C309 source.n148 a_n2982_n2088# 0.01482f
C310 source.n149 a_n2982_n2088# 0.026047f
C311 source.n150 a_n2982_n2088# 0.013996f
C312 source.n151 a_n2982_n2088# 0.033082f
C313 source.n152 a_n2982_n2088# 0.01482f
C314 source.n153 a_n2982_n2088# 0.111461f
C315 source.t31 a_n2982_n2088# 0.05392f
C316 source.n154 a_n2982_n2088# 0.024812f
C317 source.n155 a_n2982_n2088# 0.019541f
C318 source.n156 a_n2982_n2088# 0.013996f
C319 source.n157 a_n2982_n2088# 0.619755f
C320 source.n158 a_n2982_n2088# 0.026047f
C321 source.n159 a_n2982_n2088# 0.013996f
C322 source.n160 a_n2982_n2088# 0.01482f
C323 source.n161 a_n2982_n2088# 0.033082f
C324 source.n162 a_n2982_n2088# 0.033082f
C325 source.n163 a_n2982_n2088# 0.01482f
C326 source.n164 a_n2982_n2088# 0.013996f
C327 source.n165 a_n2982_n2088# 0.026047f
C328 source.n166 a_n2982_n2088# 0.026047f
C329 source.n167 a_n2982_n2088# 0.013996f
C330 source.n168 a_n2982_n2088# 0.01482f
C331 source.n169 a_n2982_n2088# 0.033082f
C332 source.n170 a_n2982_n2088# 0.071617f
C333 source.n171 a_n2982_n2088# 0.01482f
C334 source.n172 a_n2982_n2088# 0.013996f
C335 source.n173 a_n2982_n2088# 0.060206f
C336 source.n174 a_n2982_n2088# 0.040073f
C337 source.n175 a_n2982_n2088# 1.02411f
C338 source.t32 a_n2982_n2088# 0.123497f
C339 source.t29 a_n2982_n2088# 0.123497f
C340 source.n176 a_n2982_n2088# 0.9618f
C341 source.n177 a_n2982_n2088# 0.393214f
C342 source.t21 a_n2982_n2088# 0.123497f
C343 source.t22 a_n2982_n2088# 0.123497f
C344 source.n178 a_n2982_n2088# 0.9618f
C345 source.n179 a_n2982_n2088# 0.393214f
C346 source.t36 a_n2982_n2088# 0.123497f
C347 source.t38 a_n2982_n2088# 0.123497f
C348 source.n180 a_n2982_n2088# 0.9618f
C349 source.n181 a_n2982_n2088# 0.393214f
C350 source.t30 a_n2982_n2088# 0.123497f
C351 source.t26 a_n2982_n2088# 0.123497f
C352 source.n182 a_n2982_n2088# 0.9618f
C353 source.n183 a_n2982_n2088# 0.393214f
C354 source.n184 a_n2982_n2088# 0.036611f
C355 source.n185 a_n2982_n2088# 0.026047f
C356 source.n186 a_n2982_n2088# 0.013996f
C357 source.n187 a_n2982_n2088# 0.033082f
C358 source.n188 a_n2982_n2088# 0.01482f
C359 source.n189 a_n2982_n2088# 0.026047f
C360 source.n190 a_n2982_n2088# 0.013996f
C361 source.n191 a_n2982_n2088# 0.033082f
C362 source.n192 a_n2982_n2088# 0.01482f
C363 source.n193 a_n2982_n2088# 0.111461f
C364 source.t27 a_n2982_n2088# 0.05392f
C365 source.n194 a_n2982_n2088# 0.024812f
C366 source.n195 a_n2982_n2088# 0.019541f
C367 source.n196 a_n2982_n2088# 0.013996f
C368 source.n197 a_n2982_n2088# 0.619755f
C369 source.n198 a_n2982_n2088# 0.026047f
C370 source.n199 a_n2982_n2088# 0.013996f
C371 source.n200 a_n2982_n2088# 0.01482f
C372 source.n201 a_n2982_n2088# 0.033082f
C373 source.n202 a_n2982_n2088# 0.033082f
C374 source.n203 a_n2982_n2088# 0.01482f
C375 source.n204 a_n2982_n2088# 0.013996f
C376 source.n205 a_n2982_n2088# 0.026047f
C377 source.n206 a_n2982_n2088# 0.026047f
C378 source.n207 a_n2982_n2088# 0.013996f
C379 source.n208 a_n2982_n2088# 0.01482f
C380 source.n209 a_n2982_n2088# 0.033082f
C381 source.n210 a_n2982_n2088# 0.071617f
C382 source.n211 a_n2982_n2088# 0.01482f
C383 source.n212 a_n2982_n2088# 0.013996f
C384 source.n213 a_n2982_n2088# 0.060206f
C385 source.n214 a_n2982_n2088# 0.040073f
C386 source.n215 a_n2982_n2088# 0.1362f
C387 source.n216 a_n2982_n2088# 0.036611f
C388 source.n217 a_n2982_n2088# 0.026047f
C389 source.n218 a_n2982_n2088# 0.013996f
C390 source.n219 a_n2982_n2088# 0.033082f
C391 source.n220 a_n2982_n2088# 0.01482f
C392 source.n221 a_n2982_n2088# 0.026047f
C393 source.n222 a_n2982_n2088# 0.013996f
C394 source.n223 a_n2982_n2088# 0.033082f
C395 source.n224 a_n2982_n2088# 0.01482f
C396 source.n225 a_n2982_n2088# 0.111461f
C397 source.t10 a_n2982_n2088# 0.05392f
C398 source.n226 a_n2982_n2088# 0.024812f
C399 source.n227 a_n2982_n2088# 0.019541f
C400 source.n228 a_n2982_n2088# 0.013996f
C401 source.n229 a_n2982_n2088# 0.619755f
C402 source.n230 a_n2982_n2088# 0.026047f
C403 source.n231 a_n2982_n2088# 0.013996f
C404 source.n232 a_n2982_n2088# 0.01482f
C405 source.n233 a_n2982_n2088# 0.033082f
C406 source.n234 a_n2982_n2088# 0.033082f
C407 source.n235 a_n2982_n2088# 0.01482f
C408 source.n236 a_n2982_n2088# 0.013996f
C409 source.n237 a_n2982_n2088# 0.026047f
C410 source.n238 a_n2982_n2088# 0.026047f
C411 source.n239 a_n2982_n2088# 0.013996f
C412 source.n240 a_n2982_n2088# 0.01482f
C413 source.n241 a_n2982_n2088# 0.033082f
C414 source.n242 a_n2982_n2088# 0.071617f
C415 source.n243 a_n2982_n2088# 0.01482f
C416 source.n244 a_n2982_n2088# 0.013996f
C417 source.n245 a_n2982_n2088# 0.060206f
C418 source.n246 a_n2982_n2088# 0.040073f
C419 source.n247 a_n2982_n2088# 0.1362f
C420 source.t12 a_n2982_n2088# 0.123497f
C421 source.t15 a_n2982_n2088# 0.123497f
C422 source.n248 a_n2982_n2088# 0.9618f
C423 source.n249 a_n2982_n2088# 0.393214f
C424 source.t17 a_n2982_n2088# 0.123497f
C425 source.t16 a_n2982_n2088# 0.123497f
C426 source.n250 a_n2982_n2088# 0.9618f
C427 source.n251 a_n2982_n2088# 0.393214f
C428 source.t8 a_n2982_n2088# 0.123497f
C429 source.t19 a_n2982_n2088# 0.123497f
C430 source.n252 a_n2982_n2088# 0.9618f
C431 source.n253 a_n2982_n2088# 0.393214f
C432 source.t2 a_n2982_n2088# 0.123497f
C433 source.t1 a_n2982_n2088# 0.123497f
C434 source.n254 a_n2982_n2088# 0.9618f
C435 source.n255 a_n2982_n2088# 0.393214f
C436 source.n256 a_n2982_n2088# 0.036611f
C437 source.n257 a_n2982_n2088# 0.026047f
C438 source.n258 a_n2982_n2088# 0.013996f
C439 source.n259 a_n2982_n2088# 0.033082f
C440 source.n260 a_n2982_n2088# 0.01482f
C441 source.n261 a_n2982_n2088# 0.026047f
C442 source.n262 a_n2982_n2088# 0.013996f
C443 source.n263 a_n2982_n2088# 0.033082f
C444 source.n264 a_n2982_n2088# 0.01482f
C445 source.n265 a_n2982_n2088# 0.111461f
C446 source.t4 a_n2982_n2088# 0.05392f
C447 source.n266 a_n2982_n2088# 0.024812f
C448 source.n267 a_n2982_n2088# 0.019541f
C449 source.n268 a_n2982_n2088# 0.013996f
C450 source.n269 a_n2982_n2088# 0.619755f
C451 source.n270 a_n2982_n2088# 0.026047f
C452 source.n271 a_n2982_n2088# 0.013996f
C453 source.n272 a_n2982_n2088# 0.01482f
C454 source.n273 a_n2982_n2088# 0.033082f
C455 source.n274 a_n2982_n2088# 0.033082f
C456 source.n275 a_n2982_n2088# 0.01482f
C457 source.n276 a_n2982_n2088# 0.013996f
C458 source.n277 a_n2982_n2088# 0.026047f
C459 source.n278 a_n2982_n2088# 0.026047f
C460 source.n279 a_n2982_n2088# 0.013996f
C461 source.n280 a_n2982_n2088# 0.01482f
C462 source.n281 a_n2982_n2088# 0.033082f
C463 source.n282 a_n2982_n2088# 0.071617f
C464 source.n283 a_n2982_n2088# 0.01482f
C465 source.n284 a_n2982_n2088# 0.013996f
C466 source.n285 a_n2982_n2088# 0.060206f
C467 source.n286 a_n2982_n2088# 0.040073f
C468 source.n287 a_n2982_n2088# 0.306103f
C469 source.n288 a_n2982_n2088# 1.08021f
C470 drain_left.t9 a_n2982_n2088# 0.129288f
C471 drain_left.t17 a_n2982_n2088# 0.129288f
C472 drain_left.n0 a_n2982_n2088# 1.08333f
C473 drain_left.t14 a_n2982_n2088# 0.129288f
C474 drain_left.t7 a_n2982_n2088# 0.129288f
C475 drain_left.n1 a_n2982_n2088# 1.07826f
C476 drain_left.n2 a_n2982_n2088# 0.756516f
C477 drain_left.t13 a_n2982_n2088# 0.129288f
C478 drain_left.t3 a_n2982_n2088# 0.129288f
C479 drain_left.n3 a_n2982_n2088# 1.07826f
C480 drain_left.t18 a_n2982_n2088# 0.129288f
C481 drain_left.t4 a_n2982_n2088# 0.129288f
C482 drain_left.n4 a_n2982_n2088# 1.08333f
C483 drain_left.t5 a_n2982_n2088# 0.129288f
C484 drain_left.t0 a_n2982_n2088# 0.129288f
C485 drain_left.n5 a_n2982_n2088# 1.07826f
C486 drain_left.n6 a_n2982_n2088# 0.756516f
C487 drain_left.n7 a_n2982_n2088# 1.62289f
C488 drain_left.t16 a_n2982_n2088# 0.129288f
C489 drain_left.t12 a_n2982_n2088# 0.129288f
C490 drain_left.n8 a_n2982_n2088# 1.08333f
C491 drain_left.t8 a_n2982_n2088# 0.129288f
C492 drain_left.t15 a_n2982_n2088# 0.129288f
C493 drain_left.n9 a_n2982_n2088# 1.07827f
C494 drain_left.n10 a_n2982_n2088# 0.760609f
C495 drain_left.t6 a_n2982_n2088# 0.129288f
C496 drain_left.t19 a_n2982_n2088# 0.129288f
C497 drain_left.n11 a_n2982_n2088# 1.07827f
C498 drain_left.n12 a_n2982_n2088# 0.377346f
C499 drain_left.t10 a_n2982_n2088# 0.129288f
C500 drain_left.t1 a_n2982_n2088# 0.129288f
C501 drain_left.n13 a_n2982_n2088# 1.07827f
C502 drain_left.n14 a_n2982_n2088# 0.377346f
C503 drain_left.t2 a_n2982_n2088# 0.129288f
C504 drain_left.t11 a_n2982_n2088# 0.129288f
C505 drain_left.n15 a_n2982_n2088# 1.07826f
C506 drain_left.n16 a_n2982_n2088# 0.618538f
C507 plus.n0 a_n2982_n2088# 0.041429f
C508 plus.t4 a_n2982_n2088# 0.5047f
C509 plus.t19 a_n2982_n2088# 0.5047f
C510 plus.n1 a_n2982_n2088# 0.041429f
C511 plus.t11 a_n2982_n2088# 0.5047f
C512 plus.n2 a_n2982_n2088# 0.233217f
C513 plus.n3 a_n2982_n2088# 0.041429f
C514 plus.t0 a_n2982_n2088# 0.5047f
C515 plus.t15 a_n2982_n2088# 0.5047f
C516 plus.n4 a_n2982_n2088# 0.233217f
C517 plus.n5 a_n2982_n2088# 0.041429f
C518 plus.t5 a_n2982_n2088# 0.5047f
C519 plus.t14 a_n2982_n2088# 0.5047f
C520 plus.n6 a_n2982_n2088# 0.233217f
C521 plus.n7 a_n2982_n2088# 0.041429f
C522 plus.t2 a_n2982_n2088# 0.5047f
C523 plus.t16 a_n2982_n2088# 0.5047f
C524 plus.n8 a_n2982_n2088# 0.240146f
C525 plus.t6 a_n2982_n2088# 0.525295f
C526 plus.n9 a_n2982_n2088# 0.215597f
C527 plus.n10 a_n2982_n2088# 0.176835f
C528 plus.n11 a_n2982_n2088# 0.009401f
C529 plus.n12 a_n2982_n2088# 0.233217f
C530 plus.n13 a_n2982_n2088# 0.009401f
C531 plus.n14 a_n2982_n2088# 0.041429f
C532 plus.n15 a_n2982_n2088# 0.041429f
C533 plus.n16 a_n2982_n2088# 0.041429f
C534 plus.n17 a_n2982_n2088# 0.009401f
C535 plus.n18 a_n2982_n2088# 0.233217f
C536 plus.n19 a_n2982_n2088# 0.009401f
C537 plus.n20 a_n2982_n2088# 0.041429f
C538 plus.n21 a_n2982_n2088# 0.041429f
C539 plus.n22 a_n2982_n2088# 0.041429f
C540 plus.n23 a_n2982_n2088# 0.009401f
C541 plus.n24 a_n2982_n2088# 0.233217f
C542 plus.n25 a_n2982_n2088# 0.009401f
C543 plus.n26 a_n2982_n2088# 0.041429f
C544 plus.n27 a_n2982_n2088# 0.041429f
C545 plus.n28 a_n2982_n2088# 0.041429f
C546 plus.n29 a_n2982_n2088# 0.009401f
C547 plus.n30 a_n2982_n2088# 0.233217f
C548 plus.n31 a_n2982_n2088# 0.009401f
C549 plus.n32 a_n2982_n2088# 0.232834f
C550 plus.n33 a_n2982_n2088# 0.371924f
C551 plus.n34 a_n2982_n2088# 0.041429f
C552 plus.t8 a_n2982_n2088# 0.5047f
C553 plus.n35 a_n2982_n2088# 0.041429f
C554 plus.t7 a_n2982_n2088# 0.5047f
C555 plus.t10 a_n2982_n2088# 0.5047f
C556 plus.n36 a_n2982_n2088# 0.233217f
C557 plus.n37 a_n2982_n2088# 0.041429f
C558 plus.t18 a_n2982_n2088# 0.5047f
C559 plus.t17 a_n2982_n2088# 0.5047f
C560 plus.n38 a_n2982_n2088# 0.233217f
C561 plus.n39 a_n2982_n2088# 0.041429f
C562 plus.t3 a_n2982_n2088# 0.5047f
C563 plus.t1 a_n2982_n2088# 0.5047f
C564 plus.n40 a_n2982_n2088# 0.233217f
C565 plus.n41 a_n2982_n2088# 0.041429f
C566 plus.t9 a_n2982_n2088# 0.5047f
C567 plus.t13 a_n2982_n2088# 0.5047f
C568 plus.n42 a_n2982_n2088# 0.240146f
C569 plus.t12 a_n2982_n2088# 0.525295f
C570 plus.n43 a_n2982_n2088# 0.215597f
C571 plus.n44 a_n2982_n2088# 0.176835f
C572 plus.n45 a_n2982_n2088# 0.009401f
C573 plus.n46 a_n2982_n2088# 0.233217f
C574 plus.n47 a_n2982_n2088# 0.009401f
C575 plus.n48 a_n2982_n2088# 0.041429f
C576 plus.n49 a_n2982_n2088# 0.041429f
C577 plus.n50 a_n2982_n2088# 0.041429f
C578 plus.n51 a_n2982_n2088# 0.009401f
C579 plus.n52 a_n2982_n2088# 0.233217f
C580 plus.n53 a_n2982_n2088# 0.009401f
C581 plus.n54 a_n2982_n2088# 0.041429f
C582 plus.n55 a_n2982_n2088# 0.041429f
C583 plus.n56 a_n2982_n2088# 0.041429f
C584 plus.n57 a_n2982_n2088# 0.009401f
C585 plus.n58 a_n2982_n2088# 0.233217f
C586 plus.n59 a_n2982_n2088# 0.009401f
C587 plus.n60 a_n2982_n2088# 0.041429f
C588 plus.n61 a_n2982_n2088# 0.041429f
C589 plus.n62 a_n2982_n2088# 0.041429f
C590 plus.n63 a_n2982_n2088# 0.009401f
C591 plus.n64 a_n2982_n2088# 0.233217f
C592 plus.n65 a_n2982_n2088# 0.009401f
C593 plus.n66 a_n2982_n2088# 0.232834f
C594 plus.n67 a_n2982_n2088# 1.32398f
.ends

