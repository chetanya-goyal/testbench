* NGSPICE file created from diffpair212.ext - technology: sky130A

.subckt diffpair212 minus drain_right drain_left source plus
X0 drain_right.t5 minus.t0 source.t8 a_n1460_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X1 a_n1460_n1488# a_n1460_n1488# a_n1460_n1488# a_n1460_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.6
X2 a_n1460_n1488# a_n1460_n1488# a_n1460_n1488# a_n1460_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X3 a_n1460_n1488# a_n1460_n1488# a_n1460_n1488# a_n1460_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X4 source.t9 minus.t1 drain_right.t4 a_n1460_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X5 drain_left.t5 plus.t0 source.t5 a_n1460_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X6 drain_right.t3 minus.t2 source.t7 a_n1460_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X7 source.t10 minus.t3 drain_right.t2 a_n1460_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X8 drain_left.t4 plus.t1 source.t2 a_n1460_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X9 drain_right.t1 minus.t4 source.t11 a_n1460_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X10 drain_right.t0 minus.t5 source.t6 a_n1460_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X11 source.t0 plus.t2 drain_left.t3 a_n1460_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X12 drain_left.t2 plus.t3 source.t4 a_n1460_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X13 drain_left.t1 plus.t4 source.t1 a_n1460_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X14 a_n1460_n1488# a_n1460_n1488# a_n1460_n1488# a_n1460_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X15 source.t3 plus.t5 drain_left.t0 a_n1460_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
R0 minus.n0 minus.t4 212.793
R1 minus.n4 minus.t5 212.793
R2 minus.n1 minus.t3 185.972
R3 minus.n2 minus.t2 185.972
R4 minus.n5 minus.t1 185.972
R5 minus.n6 minus.t0 185.972
R6 minus.n3 minus.n2 161.3
R7 minus.n7 minus.n6 161.3
R8 minus.n2 minus.n1 48.2005
R9 minus.n6 minus.n5 48.2005
R10 minus.n3 minus.n0 45.1367
R11 minus.n7 minus.n4 45.1367
R12 minus.n8 minus.n3 27.9607
R13 minus.n1 minus.n0 13.3799
R14 minus.n5 minus.n4 13.3799
R15 minus.n8 minus.n7 6.62739
R16 minus minus.n8 0.188
R17 source.n0 source.t2 69.6943
R18 source.n3 source.t11 69.6943
R19 source.n11 source.t8 69.6942
R20 source.n8 source.t5 69.6942
R21 source.n2 source.n1 63.0943
R22 source.n5 source.n4 63.0943
R23 source.n10 source.n9 63.0942
R24 source.n7 source.n6 63.0942
R25 source.n7 source.n5 16.073
R26 source.n12 source.n0 9.60747
R27 source.n9 source.t6 6.6005
R28 source.n9 source.t9 6.6005
R29 source.n6 source.t1 6.6005
R30 source.n6 source.t3 6.6005
R31 source.n1 source.t4 6.6005
R32 source.n1 source.t0 6.6005
R33 source.n4 source.t7 6.6005
R34 source.n4 source.t10 6.6005
R35 source.n12 source.n11 5.66429
R36 source.n3 source.n2 0.87119
R37 source.n10 source.n8 0.87119
R38 source.n5 source.n3 0.802224
R39 source.n2 source.n0 0.802224
R40 source.n8 source.n7 0.802224
R41 source.n11 source.n10 0.802224
R42 source source.n12 0.188
R43 drain_right.n1 drain_right.t0 86.9189
R44 drain_right.n3 drain_right.t3 86.3731
R45 drain_right.n3 drain_right.n2 80.5748
R46 drain_right.n1 drain_right.n0 79.9181
R47 drain_right drain_right.n1 22.2004
R48 drain_right.n0 drain_right.t4 6.6005
R49 drain_right.n0 drain_right.t5 6.6005
R50 drain_right.n2 drain_right.t2 6.6005
R51 drain_right.n2 drain_right.t1 6.6005
R52 drain_right drain_right.n3 6.05408
R53 plus.n0 plus.t3 212.793
R54 plus.n4 plus.t0 212.793
R55 plus.n2 plus.t1 185.972
R56 plus.n1 plus.t2 185.972
R57 plus.n6 plus.t4 185.972
R58 plus.n5 plus.t5 185.972
R59 plus.n3 plus.n2 161.3
R60 plus.n7 plus.n6 161.3
R61 plus.n2 plus.n1 48.2005
R62 plus.n6 plus.n5 48.2005
R63 plus.n3 plus.n0 45.1367
R64 plus.n7 plus.n4 45.1367
R65 plus plus.n7 25.2509
R66 plus.n1 plus.n0 13.3799
R67 plus.n5 plus.n4 13.3799
R68 plus plus.n3 8.86224
R69 drain_left.n3 drain_left.t2 87.1748
R70 drain_left.n1 drain_left.t1 86.9189
R71 drain_left.n1 drain_left.n0 79.9181
R72 drain_left.n3 drain_left.n2 79.7731
R73 drain_left drain_left.n1 22.7536
R74 drain_left.n0 drain_left.t0 6.6005
R75 drain_left.n0 drain_left.t5 6.6005
R76 drain_left.n2 drain_left.t3 6.6005
R77 drain_left.n2 drain_left.t4 6.6005
R78 drain_left drain_left.n3 6.45494
C0 drain_left drain_right 0.671668f
C1 drain_left source 4.05921f
C2 drain_right plus 0.299377f
C3 minus drain_left 0.176422f
C4 source plus 1.37031f
C5 minus plus 3.30107f
C6 source drain_right 4.05714f
C7 minus drain_right 1.25458f
C8 minus source 1.35618f
C9 drain_left plus 1.39297f
C10 drain_right a_n1460_n1488# 3.433244f
C11 drain_left a_n1460_n1488# 3.62875f
C12 source a_n1460_n1488# 2.846137f
C13 minus a_n1460_n1488# 4.850642f
C14 plus a_n1460_n1488# 5.461979f
C15 drain_left.t1 a_n1460_n1488# 0.394208f
C16 drain_left.t0 a_n1460_n1488# 0.042445f
C17 drain_left.t5 a_n1460_n1488# 0.042445f
C18 drain_left.n0 a_n1460_n1488# 0.306489f
C19 drain_left.n1 a_n1460_n1488# 0.902912f
C20 drain_left.t2 a_n1460_n1488# 0.394956f
C21 drain_left.t3 a_n1460_n1488# 0.042445f
C22 drain_left.t4 a_n1460_n1488# 0.042445f
C23 drain_left.n2 a_n1460_n1488# 0.306112f
C24 drain_left.n3 a_n1460_n1488# 0.615646f
C25 plus.t3 a_n1460_n1488# 0.165558f
C26 plus.n0 a_n1460_n1488# 0.080226f
C27 plus.t1 a_n1460_n1488# 0.154064f
C28 plus.t2 a_n1460_n1488# 0.154064f
C29 plus.n1 a_n1460_n1488# 0.097585f
C30 plus.n2 a_n1460_n1488# 0.091108f
C31 plus.n3 a_n1460_n1488# 0.3153f
C32 plus.t0 a_n1460_n1488# 0.165558f
C33 plus.n4 a_n1460_n1488# 0.080226f
C34 plus.t4 a_n1460_n1488# 0.154064f
C35 plus.t5 a_n1460_n1488# 0.154064f
C36 plus.n5 a_n1460_n1488# 0.097585f
C37 plus.n6 a_n1460_n1488# 0.091108f
C38 plus.n7 a_n1460_n1488# 0.716859f
C39 drain_right.t0 a_n1460_n1488# 0.401059f
C40 drain_right.t4 a_n1460_n1488# 0.043183f
C41 drain_right.t5 a_n1460_n1488# 0.043183f
C42 drain_right.n0 a_n1460_n1488# 0.311815f
C43 drain_right.n1 a_n1460_n1488# 0.882326f
C44 drain_right.t2 a_n1460_n1488# 0.043183f
C45 drain_right.t1 a_n1460_n1488# 0.043183f
C46 drain_right.n2 a_n1460_n1488# 0.313893f
C47 drain_right.t3 a_n1460_n1488# 0.399707f
C48 drain_right.n3 a_n1460_n1488# 0.638074f
C49 source.t2 a_n1460_n1488# 0.42751f
C50 source.n0 a_n1460_n1488# 0.615076f
C51 source.t4 a_n1460_n1488# 0.051484f
C52 source.t0 a_n1460_n1488# 0.051484f
C53 source.n1 a_n1460_n1488# 0.326435f
C54 source.n2 a_n1460_n1488# 0.306209f
C55 source.t11 a_n1460_n1488# 0.42751f
C56 source.n3 a_n1460_n1488# 0.345543f
C57 source.t7 a_n1460_n1488# 0.051484f
C58 source.t10 a_n1460_n1488# 0.051484f
C59 source.n4 a_n1460_n1488# 0.326435f
C60 source.n5 a_n1460_n1488# 0.862595f
C61 source.t1 a_n1460_n1488# 0.051484f
C62 source.t3 a_n1460_n1488# 0.051484f
C63 source.n6 a_n1460_n1488# 0.326432f
C64 source.n7 a_n1460_n1488# 0.862597f
C65 source.t5 a_n1460_n1488# 0.427508f
C66 source.n8 a_n1460_n1488# 0.345546f
C67 source.t6 a_n1460_n1488# 0.051484f
C68 source.t9 a_n1460_n1488# 0.051484f
C69 source.n9 a_n1460_n1488# 0.326432f
C70 source.n10 a_n1460_n1488# 0.306211f
C71 source.t8 a_n1460_n1488# 0.427508f
C72 source.n11 a_n1460_n1488# 0.454427f
C73 source.n12 a_n1460_n1488# 0.637602f
C74 minus.t4 a_n1460_n1488# 0.162712f
C75 minus.n0 a_n1460_n1488# 0.078847f
C76 minus.t3 a_n1460_n1488# 0.151416f
C77 minus.n1 a_n1460_n1488# 0.095908f
C78 minus.t2 a_n1460_n1488# 0.151416f
C79 minus.n2 a_n1460_n1488# 0.089542f
C80 minus.n3 a_n1460_n1488# 0.740756f
C81 minus.t5 a_n1460_n1488# 0.162712f
C82 minus.n4 a_n1460_n1488# 0.078847f
C83 minus.t1 a_n1460_n1488# 0.151416f
C84 minus.n5 a_n1460_n1488# 0.095908f
C85 minus.t0 a_n1460_n1488# 0.151416f
C86 minus.n6 a_n1460_n1488# 0.089542f
C87 minus.n7 a_n1460_n1488# 0.283283f
C88 minus.n8 a_n1460_n1488# 0.79786f
.ends

