* NGSPICE file created from diffpair153.ext - technology: sky130A

.subckt diffpair153 minus drain_right drain_left source plus
X0 a_n1846_n1288# a_n1846_n1288# a_n1846_n1288# a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.8
X1 a_n1846_n1288# a_n1846_n1288# a_n1846_n1288# a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X2 drain_right.t7 minus.t0 source.t8 a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X3 drain_right.t6 minus.t1 source.t15 a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X4 a_n1846_n1288# a_n1846_n1288# a_n1846_n1288# a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X5 source.t7 plus.t0 drain_left.t7 a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X6 source.t4 plus.t1 drain_left.t6 a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X7 a_n1846_n1288# a_n1846_n1288# a_n1846_n1288# a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X8 drain_right.t5 minus.t2 source.t14 a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X9 source.t13 minus.t3 drain_right.t4 a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X10 drain_right.t3 minus.t4 source.t11 a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X11 source.t9 minus.t5 drain_right.t2 a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X12 drain_left.t5 plus.t2 source.t5 a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X13 source.t12 minus.t6 drain_right.t1 a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X14 source.t6 plus.t3 drain_left.t4 a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X15 source.t10 minus.t7 drain_right.t0 a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X16 drain_left.t3 plus.t4 source.t2 a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X17 drain_left.t2 plus.t5 source.t0 a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X18 source.t1 plus.t6 drain_left.t1 a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X19 drain_left.t0 plus.t7 source.t3 a_n1846_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
R0 minus.n7 minus.n6 161.3
R1 minus.n5 minus.n0 161.3
R2 minus.n15 minus.n14 161.3
R3 minus.n13 minus.n8 161.3
R4 minus.n2 minus.t4 129.957
R5 minus.n10 minus.t6 129.957
R6 minus.n1 minus.t3 109.355
R7 minus.n4 minus.t2 109.355
R8 minus.n6 minus.t5 109.355
R9 minus.n9 minus.t0 109.355
R10 minus.n12 minus.t7 109.355
R11 minus.n14 minus.t1 109.355
R12 minus.n4 minus.n3 80.6037
R13 minus.n12 minus.n11 80.6037
R14 minus.n4 minus.n1 48.2005
R15 minus.n12 minus.n9 48.2005
R16 minus.n5 minus.n4 41.6278
R17 minus.n13 minus.n12 41.6278
R18 minus.n3 minus.n2 31.6158
R19 minus.n11 minus.n10 31.6158
R20 minus.n16 minus.n7 28.6899
R21 minus.n2 minus.n1 17.6494
R22 minus.n10 minus.n9 17.6494
R23 minus.n16 minus.n15 6.65202
R24 minus.n6 minus.n5 6.57323
R25 minus.n14 minus.n13 6.57323
R26 minus.n3 minus.n0 0.285035
R27 minus.n11 minus.n8 0.285035
R28 minus.n7 minus.n0 0.189894
R29 minus.n15 minus.n8 0.189894
R30 minus minus.n16 0.188
R31 source.n66 source.n64 289.615
R32 source.n56 source.n54 289.615
R33 source.n48 source.n46 289.615
R34 source.n38 source.n36 289.615
R35 source.n2 source.n0 289.615
R36 source.n12 source.n10 289.615
R37 source.n20 source.n18 289.615
R38 source.n30 source.n28 289.615
R39 source.n67 source.n66 185
R40 source.n57 source.n56 185
R41 source.n49 source.n48 185
R42 source.n39 source.n38 185
R43 source.n3 source.n2 185
R44 source.n13 source.n12 185
R45 source.n21 source.n20 185
R46 source.n31 source.n30 185
R47 source.t15 source.n65 167.117
R48 source.t12 source.n55 167.117
R49 source.t0 source.n47 167.117
R50 source.t4 source.n37 167.117
R51 source.t5 source.n1 167.117
R52 source.t1 source.n11 167.117
R53 source.t11 source.n19 167.117
R54 source.t9 source.n29 167.117
R55 source.n9 source.n8 84.1169
R56 source.n27 source.n26 84.1169
R57 source.n63 source.n62 84.1168
R58 source.n45 source.n44 84.1168
R59 source.n66 source.t15 52.3082
R60 source.n56 source.t12 52.3082
R61 source.n48 source.t0 52.3082
R62 source.n38 source.t4 52.3082
R63 source.n2 source.t5 52.3082
R64 source.n12 source.t1 52.3082
R65 source.n20 source.t11 52.3082
R66 source.n30 source.t9 52.3082
R67 source.n71 source.n70 31.4096
R68 source.n61 source.n60 31.4096
R69 source.n53 source.n52 31.4096
R70 source.n43 source.n42 31.4096
R71 source.n7 source.n6 31.4096
R72 source.n17 source.n16 31.4096
R73 source.n25 source.n24 31.4096
R74 source.n35 source.n34 31.4096
R75 source.n43 source.n35 14.6861
R76 source.n62 source.t8 9.9005
R77 source.n62 source.t10 9.9005
R78 source.n44 source.t3 9.9005
R79 source.n44 source.t7 9.9005
R80 source.n8 source.t2 9.9005
R81 source.n8 source.t6 9.9005
R82 source.n26 source.t14 9.9005
R83 source.n26 source.t13 9.9005
R84 source.n67 source.n65 9.71174
R85 source.n57 source.n55 9.71174
R86 source.n49 source.n47 9.71174
R87 source.n39 source.n37 9.71174
R88 source.n3 source.n1 9.71174
R89 source.n13 source.n11 9.71174
R90 source.n21 source.n19 9.71174
R91 source.n31 source.n29 9.71174
R92 source.n70 source.n69 9.45567
R93 source.n60 source.n59 9.45567
R94 source.n52 source.n51 9.45567
R95 source.n42 source.n41 9.45567
R96 source.n6 source.n5 9.45567
R97 source.n16 source.n15 9.45567
R98 source.n24 source.n23 9.45567
R99 source.n34 source.n33 9.45567
R100 source.n69 source.n68 9.3005
R101 source.n59 source.n58 9.3005
R102 source.n51 source.n50 9.3005
R103 source.n41 source.n40 9.3005
R104 source.n5 source.n4 9.3005
R105 source.n15 source.n14 9.3005
R106 source.n23 source.n22 9.3005
R107 source.n33 source.n32 9.3005
R108 source.n72 source.n7 8.93611
R109 source.n70 source.n64 8.14595
R110 source.n60 source.n54 8.14595
R111 source.n52 source.n46 8.14595
R112 source.n42 source.n36 8.14595
R113 source.n6 source.n0 8.14595
R114 source.n16 source.n10 8.14595
R115 source.n24 source.n18 8.14595
R116 source.n34 source.n28 8.14595
R117 source.n68 source.n67 7.3702
R118 source.n58 source.n57 7.3702
R119 source.n50 source.n49 7.3702
R120 source.n40 source.n39 7.3702
R121 source.n4 source.n3 7.3702
R122 source.n14 source.n13 7.3702
R123 source.n22 source.n21 7.3702
R124 source.n32 source.n31 7.3702
R125 source.n68 source.n64 5.81868
R126 source.n58 source.n54 5.81868
R127 source.n50 source.n46 5.81868
R128 source.n40 source.n36 5.81868
R129 source.n4 source.n0 5.81868
R130 source.n14 source.n10 5.81868
R131 source.n22 source.n18 5.81868
R132 source.n32 source.n28 5.81868
R133 source.n72 source.n71 5.7505
R134 source.n69 source.n65 3.44771
R135 source.n59 source.n55 3.44771
R136 source.n51 source.n47 3.44771
R137 source.n41 source.n37 3.44771
R138 source.n5 source.n1 3.44771
R139 source.n15 source.n11 3.44771
R140 source.n23 source.n19 3.44771
R141 source.n33 source.n29 3.44771
R142 source.n35 source.n27 0.974638
R143 source.n27 source.n25 0.974638
R144 source.n17 source.n9 0.974638
R145 source.n9 source.n7 0.974638
R146 source.n45 source.n43 0.974638
R147 source.n53 source.n45 0.974638
R148 source.n63 source.n61 0.974638
R149 source.n71 source.n63 0.974638
R150 source.n25 source.n17 0.470328
R151 source.n61 source.n53 0.470328
R152 source source.n72 0.188
R153 drain_right.n5 drain_right.n3 101.769
R154 drain_right.n2 drain_right.n1 101.228
R155 drain_right.n2 drain_right.n0 101.228
R156 drain_right.n5 drain_right.n4 100.796
R157 drain_right drain_right.n2 22.6476
R158 drain_right.n1 drain_right.t0 9.9005
R159 drain_right.n1 drain_right.t6 9.9005
R160 drain_right.n0 drain_right.t1 9.9005
R161 drain_right.n0 drain_right.t7 9.9005
R162 drain_right.n3 drain_right.t4 9.9005
R163 drain_right.n3 drain_right.t3 9.9005
R164 drain_right.n4 drain_right.t2 9.9005
R165 drain_right.n4 drain_right.t5 9.9005
R166 drain_right drain_right.n5 6.62735
R167 plus.n5 plus.n0 161.3
R168 plus.n7 plus.n6 161.3
R169 plus.n13 plus.n8 161.3
R170 plus.n15 plus.n14 161.3
R171 plus.n2 plus.t6 129.957
R172 plus.n10 plus.t5 129.957
R173 plus.n6 plus.t2 109.355
R174 plus.n4 plus.t3 109.355
R175 plus.n3 plus.t4 109.355
R176 plus.n14 plus.t1 109.355
R177 plus.n12 plus.t7 109.355
R178 plus.n11 plus.t0 109.355
R179 plus.n4 plus.n1 80.6037
R180 plus.n12 plus.n9 80.6037
R181 plus.n4 plus.n3 48.2005
R182 plus.n12 plus.n11 48.2005
R183 plus.n5 plus.n4 41.6278
R184 plus.n13 plus.n12 41.6278
R185 plus.n2 plus.n1 31.6158
R186 plus.n10 plus.n9 31.6158
R187 plus plus.n15 26.3589
R188 plus.n3 plus.n2 17.6494
R189 plus.n11 plus.n10 17.6494
R190 plus plus.n7 8.50808
R191 plus.n6 plus.n5 6.57323
R192 plus.n14 plus.n13 6.57323
R193 plus.n1 plus.n0 0.285035
R194 plus.n9 plus.n8 0.285035
R195 plus.n7 plus.n0 0.189894
R196 plus.n15 plus.n8 0.189894
R197 drain_left.n5 drain_left.n3 101.769
R198 drain_left.n2 drain_left.n1 101.228
R199 drain_left.n2 drain_left.n0 101.228
R200 drain_left.n5 drain_left.n4 100.796
R201 drain_left drain_left.n2 23.2008
R202 drain_left.n1 drain_left.t7 9.9005
R203 drain_left.n1 drain_left.t2 9.9005
R204 drain_left.n0 drain_left.t6 9.9005
R205 drain_left.n0 drain_left.t0 9.9005
R206 drain_left.n4 drain_left.t4 9.9005
R207 drain_left.n4 drain_left.t5 9.9005
R208 drain_left.n3 drain_left.t1 9.9005
R209 drain_left.n3 drain_left.t3 9.9005
R210 drain_left drain_left.n5 6.62735
C0 drain_left minus 0.177367f
C1 drain_right source 3.65952f
C2 drain_left drain_right 0.873724f
C3 drain_right minus 1.31382f
C4 plus source 1.6433f
C5 drain_left plus 1.49299f
C6 plus minus 3.599f
C7 drain_right plus 0.340514f
C8 drain_left source 3.65713f
C9 source minus 1.62934f
C10 drain_right a_n1846_n1288# 3.38502f
C11 drain_left a_n1846_n1288# 3.61f
C12 source a_n1846_n1288# 3.114882f
C13 minus a_n1846_n1288# 6.338142f
C14 plus a_n1846_n1288# 6.878961f
C15 drain_left.t6 a_n1846_n1288# 0.029128f
C16 drain_left.t0 a_n1846_n1288# 0.029128f
C17 drain_left.n0 a_n1846_n1288# 0.183985f
C18 drain_left.t7 a_n1846_n1288# 0.029128f
C19 drain_left.t2 a_n1846_n1288# 0.029128f
C20 drain_left.n1 a_n1846_n1288# 0.183985f
C21 drain_left.n2 a_n1846_n1288# 1.01131f
C22 drain_left.t1 a_n1846_n1288# 0.029128f
C23 drain_left.t3 a_n1846_n1288# 0.029128f
C24 drain_left.n3 a_n1846_n1288# 0.185521f
C25 drain_left.t4 a_n1846_n1288# 0.029128f
C26 drain_left.t5 a_n1846_n1288# 0.029128f
C27 drain_left.n4 a_n1846_n1288# 0.182992f
C28 drain_left.n5 a_n1846_n1288# 0.683679f
C29 plus.n0 a_n1846_n1288# 0.033866f
C30 plus.t2 a_n1846_n1288# 0.125749f
C31 plus.t3 a_n1846_n1288# 0.125749f
C32 plus.n1 a_n1846_n1288# 0.145255f
C33 plus.t4 a_n1846_n1288# 0.125749f
C34 plus.t6 a_n1846_n1288# 0.139605f
C35 plus.n2 a_n1846_n1288# 0.075665f
C36 plus.n3 a_n1846_n1288# 0.092595f
C37 plus.n4 a_n1846_n1288# 0.092181f
C38 plus.n5 a_n1846_n1288# 0.005759f
C39 plus.n6 a_n1846_n1288# 0.082667f
C40 plus.n7 a_n1846_n1288# 0.190954f
C41 plus.n8 a_n1846_n1288# 0.033866f
C42 plus.t1 a_n1846_n1288# 0.125749f
C43 plus.n9 a_n1846_n1288# 0.145255f
C44 plus.t7 a_n1846_n1288# 0.125749f
C45 plus.t5 a_n1846_n1288# 0.139605f
C46 plus.n10 a_n1846_n1288# 0.075665f
C47 plus.t0 a_n1846_n1288# 0.125749f
C48 plus.n11 a_n1846_n1288# 0.092595f
C49 plus.n12 a_n1846_n1288# 0.092181f
C50 plus.n13 a_n1846_n1288# 0.005759f
C51 plus.n14 a_n1846_n1288# 0.082667f
C52 plus.n15 a_n1846_n1288# 0.587436f
C53 drain_right.t1 a_n1846_n1288# 0.029707f
C54 drain_right.t7 a_n1846_n1288# 0.029707f
C55 drain_right.n0 a_n1846_n1288# 0.187641f
C56 drain_right.t0 a_n1846_n1288# 0.029707f
C57 drain_right.t6 a_n1846_n1288# 0.029707f
C58 drain_right.n1 a_n1846_n1288# 0.187641f
C59 drain_right.n2 a_n1846_n1288# 0.994578f
C60 drain_right.t4 a_n1846_n1288# 0.029707f
C61 drain_right.t3 a_n1846_n1288# 0.029707f
C62 drain_right.n3 a_n1846_n1288# 0.189208f
C63 drain_right.t2 a_n1846_n1288# 0.029707f
C64 drain_right.t5 a_n1846_n1288# 0.029707f
C65 drain_right.n4 a_n1846_n1288# 0.186629f
C66 drain_right.n5 a_n1846_n1288# 0.697266f
C67 source.n0 a_n1846_n1288# 0.027453f
C68 source.n1 a_n1846_n1288# 0.060743f
C69 source.t5 a_n1846_n1288# 0.045584f
C70 source.n2 a_n1846_n1288# 0.04754f
C71 source.n3 a_n1846_n1288# 0.015325f
C72 source.n4 a_n1846_n1288# 0.010107f
C73 source.n5 a_n1846_n1288# 0.133892f
C74 source.n6 a_n1846_n1288# 0.030095f
C75 source.n7 a_n1846_n1288# 0.330234f
C76 source.t2 a_n1846_n1288# 0.029727f
C77 source.t6 a_n1846_n1288# 0.029727f
C78 source.n8 a_n1846_n1288# 0.158918f
C79 source.n9 a_n1846_n1288# 0.264309f
C80 source.n10 a_n1846_n1288# 0.027453f
C81 source.n11 a_n1846_n1288# 0.060743f
C82 source.t1 a_n1846_n1288# 0.045584f
C83 source.n12 a_n1846_n1288# 0.04754f
C84 source.n13 a_n1846_n1288# 0.015325f
C85 source.n14 a_n1846_n1288# 0.010107f
C86 source.n15 a_n1846_n1288# 0.133892f
C87 source.n16 a_n1846_n1288# 0.030095f
C88 source.n17 a_n1846_n1288# 0.102998f
C89 source.n18 a_n1846_n1288# 0.027453f
C90 source.n19 a_n1846_n1288# 0.060743f
C91 source.t11 a_n1846_n1288# 0.045584f
C92 source.n20 a_n1846_n1288# 0.04754f
C93 source.n21 a_n1846_n1288# 0.015325f
C94 source.n22 a_n1846_n1288# 0.010107f
C95 source.n23 a_n1846_n1288# 0.133892f
C96 source.n24 a_n1846_n1288# 0.030095f
C97 source.n25 a_n1846_n1288# 0.102998f
C98 source.t14 a_n1846_n1288# 0.029727f
C99 source.t13 a_n1846_n1288# 0.029727f
C100 source.n26 a_n1846_n1288# 0.158918f
C101 source.n27 a_n1846_n1288# 0.264309f
C102 source.n28 a_n1846_n1288# 0.027453f
C103 source.n29 a_n1846_n1288# 0.060743f
C104 source.t9 a_n1846_n1288# 0.045584f
C105 source.n30 a_n1846_n1288# 0.04754f
C106 source.n31 a_n1846_n1288# 0.015325f
C107 source.n32 a_n1846_n1288# 0.010107f
C108 source.n33 a_n1846_n1288# 0.133892f
C109 source.n34 a_n1846_n1288# 0.030095f
C110 source.n35 a_n1846_n1288# 0.511587f
C111 source.n36 a_n1846_n1288# 0.027453f
C112 source.n37 a_n1846_n1288# 0.060743f
C113 source.t4 a_n1846_n1288# 0.045584f
C114 source.n38 a_n1846_n1288# 0.04754f
C115 source.n39 a_n1846_n1288# 0.015325f
C116 source.n40 a_n1846_n1288# 0.010107f
C117 source.n41 a_n1846_n1288# 0.133892f
C118 source.n42 a_n1846_n1288# 0.030095f
C119 source.n43 a_n1846_n1288# 0.511587f
C120 source.t3 a_n1846_n1288# 0.029727f
C121 source.t7 a_n1846_n1288# 0.029727f
C122 source.n44 a_n1846_n1288# 0.158917f
C123 source.n45 a_n1846_n1288# 0.26431f
C124 source.n46 a_n1846_n1288# 0.027453f
C125 source.n47 a_n1846_n1288# 0.060743f
C126 source.t0 a_n1846_n1288# 0.045584f
C127 source.n48 a_n1846_n1288# 0.04754f
C128 source.n49 a_n1846_n1288# 0.015325f
C129 source.n50 a_n1846_n1288# 0.010107f
C130 source.n51 a_n1846_n1288# 0.133892f
C131 source.n52 a_n1846_n1288# 0.030095f
C132 source.n53 a_n1846_n1288# 0.102998f
C133 source.n54 a_n1846_n1288# 0.027453f
C134 source.n55 a_n1846_n1288# 0.060743f
C135 source.t12 a_n1846_n1288# 0.045584f
C136 source.n56 a_n1846_n1288# 0.04754f
C137 source.n57 a_n1846_n1288# 0.015325f
C138 source.n58 a_n1846_n1288# 0.010107f
C139 source.n59 a_n1846_n1288# 0.133892f
C140 source.n60 a_n1846_n1288# 0.030095f
C141 source.n61 a_n1846_n1288# 0.102998f
C142 source.t8 a_n1846_n1288# 0.029727f
C143 source.t10 a_n1846_n1288# 0.029727f
C144 source.n62 a_n1846_n1288# 0.158917f
C145 source.n63 a_n1846_n1288# 0.26431f
C146 source.n64 a_n1846_n1288# 0.027453f
C147 source.n65 a_n1846_n1288# 0.060743f
C148 source.t15 a_n1846_n1288# 0.045584f
C149 source.n66 a_n1846_n1288# 0.04754f
C150 source.n67 a_n1846_n1288# 0.015325f
C151 source.n68 a_n1846_n1288# 0.010107f
C152 source.n69 a_n1846_n1288# 0.133892f
C153 source.n70 a_n1846_n1288# 0.030095f
C154 source.n71 a_n1846_n1288# 0.229761f
C155 source.n72 a_n1846_n1288# 0.476557f
C156 minus.n0 a_n1846_n1288# 0.03339f
C157 minus.t3 a_n1846_n1288# 0.123982f
C158 minus.n1 a_n1846_n1288# 0.091293f
C159 minus.t2 a_n1846_n1288# 0.123982f
C160 minus.t4 a_n1846_n1288# 0.137642f
C161 minus.n2 a_n1846_n1288# 0.074601f
C162 minus.n3 a_n1846_n1288# 0.143214f
C163 minus.n4 a_n1846_n1288# 0.090885f
C164 minus.n5 a_n1846_n1288# 0.005678f
C165 minus.t5 a_n1846_n1288# 0.123982f
C166 minus.n6 a_n1846_n1288# 0.081505f
C167 minus.n7 a_n1846_n1288# 0.606327f
C168 minus.n8 a_n1846_n1288# 0.03339f
C169 minus.t0 a_n1846_n1288# 0.123982f
C170 minus.n9 a_n1846_n1288# 0.091293f
C171 minus.t6 a_n1846_n1288# 0.137642f
C172 minus.n10 a_n1846_n1288# 0.074601f
C173 minus.n11 a_n1846_n1288# 0.143214f
C174 minus.t7 a_n1846_n1288# 0.123982f
C175 minus.n12 a_n1846_n1288# 0.090885f
C176 minus.n13 a_n1846_n1288# 0.005678f
C177 minus.t1 a_n1846_n1288# 0.123982f
C178 minus.n14 a_n1846_n1288# 0.081505f
C179 minus.n15 a_n1846_n1288# 0.17249f
C180 minus.n16 a_n1846_n1288# 0.744445f
.ends

