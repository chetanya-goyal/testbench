* NGSPICE file created from diffpair449.ext - technology: sky130A

.subckt diffpair449 minus drain_right drain_left source plus
X0 drain_right.t23 minus.t0 source.t36 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.5
X1 source.t3 plus.t0 drain_left.t23 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X2 drain_left.t22 plus.t1 source.t10 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X3 a_n2874_n3288# a_n2874_n3288# a_n2874_n3288# a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.5
X4 drain_right.t22 minus.t1 source.t22 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X5 drain_right.t21 minus.t2 source.t45 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X6 drain_left.t21 plus.t2 source.t2 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.5
X7 source.t6 plus.t3 drain_left.t20 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X8 source.t33 minus.t3 drain_right.t20 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.5
X9 drain_left.t19 plus.t4 source.t13 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X10 source.t43 minus.t4 drain_right.t19 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X11 source.t19 plus.t5 drain_left.t18 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X12 source.t12 plus.t6 drain_left.t17 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.5
X13 source.t42 minus.t5 drain_right.t18 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X14 source.t30 minus.t6 drain_right.t17 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X15 drain_left.t16 plus.t7 source.t11 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X16 drain_right.t16 minus.t7 source.t29 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X17 drain_left.t15 plus.t8 source.t46 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X18 drain_right.t15 minus.t8 source.t37 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X19 drain_right.t14 minus.t9 source.t25 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X20 a_n2874_n3288# a_n2874_n3288# a_n2874_n3288# a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.5
X21 drain_left.t14 plus.t9 source.t47 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X22 source.t5 plus.t10 drain_left.t13 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X23 drain_left.t12 plus.t11 source.t0 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X24 source.t4 plus.t12 drain_left.t11 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X25 source.t27 minus.t10 drain_right.t13 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X26 drain_right.t12 minus.t11 source.t39 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X27 source.t38 minus.t12 drain_right.t11 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X28 source.t20 plus.t13 drain_left.t10 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X29 source.t40 minus.t13 drain_right.t10 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X30 source.t23 minus.t14 drain_right.t9 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X31 source.t34 minus.t15 drain_right.t8 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X32 drain_right.t7 minus.t16 source.t35 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X33 drain_left.t9 plus.t14 source.t18 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X34 drain_right.t6 minus.t17 source.t28 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.5
X35 drain_right.t5 minus.t18 source.t26 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X36 a_n2874_n3288# a_n2874_n3288# a_n2874_n3288# a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.5
X37 a_n2874_n3288# a_n2874_n3288# a_n2874_n3288# a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.5
X38 drain_left.t8 plus.t15 source.t8 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X39 drain_right.t4 minus.t19 source.t24 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X40 drain_right.t3 minus.t20 source.t41 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X41 source.t32 minus.t21 drain_right.t2 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X42 source.t14 plus.t16 drain_left.t7 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.5
X43 source.t17 plus.t17 drain_left.t6 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X44 drain_left.t5 plus.t18 source.t7 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.5
X45 source.t9 plus.t19 drain_left.t4 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X46 source.t31 minus.t22 drain_right.t1 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.5
X47 drain_left.t3 plus.t20 source.t21 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X48 source.t15 plus.t21 drain_left.t2 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X49 source.t1 plus.t22 drain_left.t1 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X50 drain_left.t0 plus.t23 source.t16 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X51 source.t44 minus.t23 drain_right.t0 a_n2874_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
R0 minus.n9 minus.t17 683.324
R1 minus.n43 minus.t3 683.324
R2 minus.n8 minus.t4 656.966
R3 minus.n7 minus.t8 656.966
R4 minus.n13 minus.t21 656.966
R5 minus.n5 minus.t7 656.966
R6 minus.n18 minus.t13 656.966
R7 minus.n20 minus.t1 656.966
R8 minus.n3 minus.t14 656.966
R9 minus.n25 minus.t19 656.966
R10 minus.n1 minus.t5 656.966
R11 minus.n30 minus.t18 656.966
R12 minus.n32 minus.t22 656.966
R13 minus.n42 minus.t2 656.966
R14 minus.n41 minus.t12 656.966
R15 minus.n47 minus.t11 656.966
R16 minus.n39 minus.t6 656.966
R17 minus.n52 minus.t16 656.966
R18 minus.n54 minus.t15 656.966
R19 minus.n37 minus.t9 656.966
R20 minus.n59 minus.t23 656.966
R21 minus.n35 minus.t20 656.966
R22 minus.n64 minus.t10 656.966
R23 minus.n66 minus.t0 656.966
R24 minus.n33 minus.n32 161.3
R25 minus.n31 minus.n0 161.3
R26 minus.n30 minus.n29 161.3
R27 minus.n28 minus.n1 161.3
R28 minus.n27 minus.n26 161.3
R29 minus.n25 minus.n2 161.3
R30 minus.n24 minus.n23 161.3
R31 minus.n22 minus.n3 161.3
R32 minus.n21 minus.n20 161.3
R33 minus.n19 minus.n4 161.3
R34 minus.n18 minus.n17 161.3
R35 minus.n16 minus.n5 161.3
R36 minus.n15 minus.n14 161.3
R37 minus.n13 minus.n6 161.3
R38 minus.n12 minus.n11 161.3
R39 minus.n10 minus.n7 161.3
R40 minus.n67 minus.n66 161.3
R41 minus.n65 minus.n34 161.3
R42 minus.n64 minus.n63 161.3
R43 minus.n62 minus.n35 161.3
R44 minus.n61 minus.n60 161.3
R45 minus.n59 minus.n36 161.3
R46 minus.n58 minus.n57 161.3
R47 minus.n56 minus.n37 161.3
R48 minus.n55 minus.n54 161.3
R49 minus.n53 minus.n38 161.3
R50 minus.n52 minus.n51 161.3
R51 minus.n50 minus.n39 161.3
R52 minus.n49 minus.n48 161.3
R53 minus.n47 minus.n40 161.3
R54 minus.n46 minus.n45 161.3
R55 minus.n44 minus.n41 161.3
R56 minus.n8 minus.n7 48.2005
R57 minus.n18 minus.n5 48.2005
R58 minus.n20 minus.n3 48.2005
R59 minus.n30 minus.n1 48.2005
R60 minus.n42 minus.n41 48.2005
R61 minus.n52 minus.n39 48.2005
R62 minus.n54 minus.n37 48.2005
R63 minus.n64 minus.n35 48.2005
R64 minus.n14 minus.n13 47.4702
R65 minus.n25 minus.n24 47.4702
R66 minus.n48 minus.n47 47.4702
R67 minus.n59 minus.n58 47.4702
R68 minus.n32 minus.n31 46.0096
R69 minus.n66 minus.n65 46.0096
R70 minus.n10 minus.n9 45.0871
R71 minus.n44 minus.n43 45.0871
R72 minus.n68 minus.n33 40.0346
R73 minus.n13 minus.n12 25.5611
R74 minus.n26 minus.n25 25.5611
R75 minus.n47 minus.n46 25.5611
R76 minus.n60 minus.n59 25.5611
R77 minus.n20 minus.n19 24.1005
R78 minus.n19 minus.n18 24.1005
R79 minus.n53 minus.n52 24.1005
R80 minus.n54 minus.n53 24.1005
R81 minus.n12 minus.n7 22.6399
R82 minus.n26 minus.n1 22.6399
R83 minus.n46 minus.n41 22.6399
R84 minus.n60 minus.n35 22.6399
R85 minus.n9 minus.n8 14.1472
R86 minus.n43 minus.n42 14.1472
R87 minus.n68 minus.n67 6.52702
R88 minus.n31 minus.n30 2.19141
R89 minus.n65 minus.n64 2.19141
R90 minus.n14 minus.n5 0.730803
R91 minus.n24 minus.n3 0.730803
R92 minus.n48 minus.n39 0.730803
R93 minus.n58 minus.n37 0.730803
R94 minus.n33 minus.n0 0.189894
R95 minus.n29 minus.n0 0.189894
R96 minus.n29 minus.n28 0.189894
R97 minus.n28 minus.n27 0.189894
R98 minus.n27 minus.n2 0.189894
R99 minus.n23 minus.n2 0.189894
R100 minus.n23 minus.n22 0.189894
R101 minus.n22 minus.n21 0.189894
R102 minus.n21 minus.n4 0.189894
R103 minus.n17 minus.n4 0.189894
R104 minus.n17 minus.n16 0.189894
R105 minus.n16 minus.n15 0.189894
R106 minus.n15 minus.n6 0.189894
R107 minus.n11 minus.n6 0.189894
R108 minus.n11 minus.n10 0.189894
R109 minus.n45 minus.n44 0.189894
R110 minus.n45 minus.n40 0.189894
R111 minus.n49 minus.n40 0.189894
R112 minus.n50 minus.n49 0.189894
R113 minus.n51 minus.n50 0.189894
R114 minus.n51 minus.n38 0.189894
R115 minus.n55 minus.n38 0.189894
R116 minus.n56 minus.n55 0.189894
R117 minus.n57 minus.n56 0.189894
R118 minus.n57 minus.n36 0.189894
R119 minus.n61 minus.n36 0.189894
R120 minus.n62 minus.n61 0.189894
R121 minus.n63 minus.n62 0.189894
R122 minus.n63 minus.n34 0.189894
R123 minus.n67 minus.n34 0.189894
R124 minus minus.n68 0.188
R125 source.n562 source.n502 289.615
R126 source.n486 source.n426 289.615
R127 source.n420 source.n360 289.615
R128 source.n344 source.n284 289.615
R129 source.n60 source.n0 289.615
R130 source.n136 source.n76 289.615
R131 source.n202 source.n142 289.615
R132 source.n278 source.n218 289.615
R133 source.n522 source.n521 185
R134 source.n527 source.n526 185
R135 source.n529 source.n528 185
R136 source.n518 source.n517 185
R137 source.n535 source.n534 185
R138 source.n537 source.n536 185
R139 source.n514 source.n513 185
R140 source.n544 source.n543 185
R141 source.n545 source.n512 185
R142 source.n547 source.n546 185
R143 source.n510 source.n509 185
R144 source.n553 source.n552 185
R145 source.n555 source.n554 185
R146 source.n506 source.n505 185
R147 source.n561 source.n560 185
R148 source.n563 source.n562 185
R149 source.n446 source.n445 185
R150 source.n451 source.n450 185
R151 source.n453 source.n452 185
R152 source.n442 source.n441 185
R153 source.n459 source.n458 185
R154 source.n461 source.n460 185
R155 source.n438 source.n437 185
R156 source.n468 source.n467 185
R157 source.n469 source.n436 185
R158 source.n471 source.n470 185
R159 source.n434 source.n433 185
R160 source.n477 source.n476 185
R161 source.n479 source.n478 185
R162 source.n430 source.n429 185
R163 source.n485 source.n484 185
R164 source.n487 source.n486 185
R165 source.n380 source.n379 185
R166 source.n385 source.n384 185
R167 source.n387 source.n386 185
R168 source.n376 source.n375 185
R169 source.n393 source.n392 185
R170 source.n395 source.n394 185
R171 source.n372 source.n371 185
R172 source.n402 source.n401 185
R173 source.n403 source.n370 185
R174 source.n405 source.n404 185
R175 source.n368 source.n367 185
R176 source.n411 source.n410 185
R177 source.n413 source.n412 185
R178 source.n364 source.n363 185
R179 source.n419 source.n418 185
R180 source.n421 source.n420 185
R181 source.n304 source.n303 185
R182 source.n309 source.n308 185
R183 source.n311 source.n310 185
R184 source.n300 source.n299 185
R185 source.n317 source.n316 185
R186 source.n319 source.n318 185
R187 source.n296 source.n295 185
R188 source.n326 source.n325 185
R189 source.n327 source.n294 185
R190 source.n329 source.n328 185
R191 source.n292 source.n291 185
R192 source.n335 source.n334 185
R193 source.n337 source.n336 185
R194 source.n288 source.n287 185
R195 source.n343 source.n342 185
R196 source.n345 source.n344 185
R197 source.n61 source.n60 185
R198 source.n59 source.n58 185
R199 source.n4 source.n3 185
R200 source.n53 source.n52 185
R201 source.n51 source.n50 185
R202 source.n8 source.n7 185
R203 source.n45 source.n44 185
R204 source.n43 source.n10 185
R205 source.n42 source.n41 185
R206 source.n13 source.n11 185
R207 source.n36 source.n35 185
R208 source.n34 source.n33 185
R209 source.n17 source.n16 185
R210 source.n28 source.n27 185
R211 source.n26 source.n25 185
R212 source.n21 source.n20 185
R213 source.n137 source.n136 185
R214 source.n135 source.n134 185
R215 source.n80 source.n79 185
R216 source.n129 source.n128 185
R217 source.n127 source.n126 185
R218 source.n84 source.n83 185
R219 source.n121 source.n120 185
R220 source.n119 source.n86 185
R221 source.n118 source.n117 185
R222 source.n89 source.n87 185
R223 source.n112 source.n111 185
R224 source.n110 source.n109 185
R225 source.n93 source.n92 185
R226 source.n104 source.n103 185
R227 source.n102 source.n101 185
R228 source.n97 source.n96 185
R229 source.n203 source.n202 185
R230 source.n201 source.n200 185
R231 source.n146 source.n145 185
R232 source.n195 source.n194 185
R233 source.n193 source.n192 185
R234 source.n150 source.n149 185
R235 source.n187 source.n186 185
R236 source.n185 source.n152 185
R237 source.n184 source.n183 185
R238 source.n155 source.n153 185
R239 source.n178 source.n177 185
R240 source.n176 source.n175 185
R241 source.n159 source.n158 185
R242 source.n170 source.n169 185
R243 source.n168 source.n167 185
R244 source.n163 source.n162 185
R245 source.n279 source.n278 185
R246 source.n277 source.n276 185
R247 source.n222 source.n221 185
R248 source.n271 source.n270 185
R249 source.n269 source.n268 185
R250 source.n226 source.n225 185
R251 source.n263 source.n262 185
R252 source.n261 source.n228 185
R253 source.n260 source.n259 185
R254 source.n231 source.n229 185
R255 source.n254 source.n253 185
R256 source.n252 source.n251 185
R257 source.n235 source.n234 185
R258 source.n246 source.n245 185
R259 source.n244 source.n243 185
R260 source.n239 source.n238 185
R261 source.n523 source.t36 149.524
R262 source.n447 source.t33 149.524
R263 source.n381 source.t7 149.524
R264 source.n305 source.t14 149.524
R265 source.n22 source.t2 149.524
R266 source.n98 source.t12 149.524
R267 source.n164 source.t28 149.524
R268 source.n240 source.t31 149.524
R269 source.n527 source.n521 104.615
R270 source.n528 source.n527 104.615
R271 source.n528 source.n517 104.615
R272 source.n535 source.n517 104.615
R273 source.n536 source.n535 104.615
R274 source.n536 source.n513 104.615
R275 source.n544 source.n513 104.615
R276 source.n545 source.n544 104.615
R277 source.n546 source.n545 104.615
R278 source.n546 source.n509 104.615
R279 source.n553 source.n509 104.615
R280 source.n554 source.n553 104.615
R281 source.n554 source.n505 104.615
R282 source.n561 source.n505 104.615
R283 source.n562 source.n561 104.615
R284 source.n451 source.n445 104.615
R285 source.n452 source.n451 104.615
R286 source.n452 source.n441 104.615
R287 source.n459 source.n441 104.615
R288 source.n460 source.n459 104.615
R289 source.n460 source.n437 104.615
R290 source.n468 source.n437 104.615
R291 source.n469 source.n468 104.615
R292 source.n470 source.n469 104.615
R293 source.n470 source.n433 104.615
R294 source.n477 source.n433 104.615
R295 source.n478 source.n477 104.615
R296 source.n478 source.n429 104.615
R297 source.n485 source.n429 104.615
R298 source.n486 source.n485 104.615
R299 source.n385 source.n379 104.615
R300 source.n386 source.n385 104.615
R301 source.n386 source.n375 104.615
R302 source.n393 source.n375 104.615
R303 source.n394 source.n393 104.615
R304 source.n394 source.n371 104.615
R305 source.n402 source.n371 104.615
R306 source.n403 source.n402 104.615
R307 source.n404 source.n403 104.615
R308 source.n404 source.n367 104.615
R309 source.n411 source.n367 104.615
R310 source.n412 source.n411 104.615
R311 source.n412 source.n363 104.615
R312 source.n419 source.n363 104.615
R313 source.n420 source.n419 104.615
R314 source.n309 source.n303 104.615
R315 source.n310 source.n309 104.615
R316 source.n310 source.n299 104.615
R317 source.n317 source.n299 104.615
R318 source.n318 source.n317 104.615
R319 source.n318 source.n295 104.615
R320 source.n326 source.n295 104.615
R321 source.n327 source.n326 104.615
R322 source.n328 source.n327 104.615
R323 source.n328 source.n291 104.615
R324 source.n335 source.n291 104.615
R325 source.n336 source.n335 104.615
R326 source.n336 source.n287 104.615
R327 source.n343 source.n287 104.615
R328 source.n344 source.n343 104.615
R329 source.n60 source.n59 104.615
R330 source.n59 source.n3 104.615
R331 source.n52 source.n3 104.615
R332 source.n52 source.n51 104.615
R333 source.n51 source.n7 104.615
R334 source.n44 source.n7 104.615
R335 source.n44 source.n43 104.615
R336 source.n43 source.n42 104.615
R337 source.n42 source.n11 104.615
R338 source.n35 source.n11 104.615
R339 source.n35 source.n34 104.615
R340 source.n34 source.n16 104.615
R341 source.n27 source.n16 104.615
R342 source.n27 source.n26 104.615
R343 source.n26 source.n20 104.615
R344 source.n136 source.n135 104.615
R345 source.n135 source.n79 104.615
R346 source.n128 source.n79 104.615
R347 source.n128 source.n127 104.615
R348 source.n127 source.n83 104.615
R349 source.n120 source.n83 104.615
R350 source.n120 source.n119 104.615
R351 source.n119 source.n118 104.615
R352 source.n118 source.n87 104.615
R353 source.n111 source.n87 104.615
R354 source.n111 source.n110 104.615
R355 source.n110 source.n92 104.615
R356 source.n103 source.n92 104.615
R357 source.n103 source.n102 104.615
R358 source.n102 source.n96 104.615
R359 source.n202 source.n201 104.615
R360 source.n201 source.n145 104.615
R361 source.n194 source.n145 104.615
R362 source.n194 source.n193 104.615
R363 source.n193 source.n149 104.615
R364 source.n186 source.n149 104.615
R365 source.n186 source.n185 104.615
R366 source.n185 source.n184 104.615
R367 source.n184 source.n153 104.615
R368 source.n177 source.n153 104.615
R369 source.n177 source.n176 104.615
R370 source.n176 source.n158 104.615
R371 source.n169 source.n158 104.615
R372 source.n169 source.n168 104.615
R373 source.n168 source.n162 104.615
R374 source.n278 source.n277 104.615
R375 source.n277 source.n221 104.615
R376 source.n270 source.n221 104.615
R377 source.n270 source.n269 104.615
R378 source.n269 source.n225 104.615
R379 source.n262 source.n225 104.615
R380 source.n262 source.n261 104.615
R381 source.n261 source.n260 104.615
R382 source.n260 source.n229 104.615
R383 source.n253 source.n229 104.615
R384 source.n253 source.n252 104.615
R385 source.n252 source.n234 104.615
R386 source.n245 source.n234 104.615
R387 source.n245 source.n244 104.615
R388 source.n244 source.n238 104.615
R389 source.t36 source.n521 52.3082
R390 source.t33 source.n445 52.3082
R391 source.t7 source.n379 52.3082
R392 source.t14 source.n303 52.3082
R393 source.t2 source.n20 52.3082
R394 source.t12 source.n96 52.3082
R395 source.t28 source.n162 52.3082
R396 source.t31 source.n238 52.3082
R397 source.n67 source.n66 42.8739
R398 source.n69 source.n68 42.8739
R399 source.n71 source.n70 42.8739
R400 source.n73 source.n72 42.8739
R401 source.n75 source.n74 42.8739
R402 source.n209 source.n208 42.8739
R403 source.n211 source.n210 42.8739
R404 source.n213 source.n212 42.8739
R405 source.n215 source.n214 42.8739
R406 source.n217 source.n216 42.8739
R407 source.n501 source.n500 42.8737
R408 source.n499 source.n498 42.8737
R409 source.n497 source.n496 42.8737
R410 source.n495 source.n494 42.8737
R411 source.n493 source.n492 42.8737
R412 source.n359 source.n358 42.8737
R413 source.n357 source.n356 42.8737
R414 source.n355 source.n354 42.8737
R415 source.n353 source.n352 42.8737
R416 source.n351 source.n350 42.8737
R417 source.n567 source.n566 29.8581
R418 source.n491 source.n490 29.8581
R419 source.n425 source.n424 29.8581
R420 source.n349 source.n348 29.8581
R421 source.n65 source.n64 29.8581
R422 source.n141 source.n140 29.8581
R423 source.n207 source.n206 29.8581
R424 source.n283 source.n282 29.8581
R425 source.n349 source.n283 22.0032
R426 source.n568 source.n65 16.3826
R427 source.n547 source.n512 13.1884
R428 source.n471 source.n436 13.1884
R429 source.n405 source.n370 13.1884
R430 source.n329 source.n294 13.1884
R431 source.n45 source.n10 13.1884
R432 source.n121 source.n86 13.1884
R433 source.n187 source.n152 13.1884
R434 source.n263 source.n228 13.1884
R435 source.n543 source.n542 12.8005
R436 source.n548 source.n510 12.8005
R437 source.n467 source.n466 12.8005
R438 source.n472 source.n434 12.8005
R439 source.n401 source.n400 12.8005
R440 source.n406 source.n368 12.8005
R441 source.n325 source.n324 12.8005
R442 source.n330 source.n292 12.8005
R443 source.n46 source.n8 12.8005
R444 source.n41 source.n12 12.8005
R445 source.n122 source.n84 12.8005
R446 source.n117 source.n88 12.8005
R447 source.n188 source.n150 12.8005
R448 source.n183 source.n154 12.8005
R449 source.n264 source.n226 12.8005
R450 source.n259 source.n230 12.8005
R451 source.n541 source.n514 12.0247
R452 source.n552 source.n551 12.0247
R453 source.n465 source.n438 12.0247
R454 source.n476 source.n475 12.0247
R455 source.n399 source.n372 12.0247
R456 source.n410 source.n409 12.0247
R457 source.n323 source.n296 12.0247
R458 source.n334 source.n333 12.0247
R459 source.n50 source.n49 12.0247
R460 source.n40 source.n13 12.0247
R461 source.n126 source.n125 12.0247
R462 source.n116 source.n89 12.0247
R463 source.n192 source.n191 12.0247
R464 source.n182 source.n155 12.0247
R465 source.n268 source.n267 12.0247
R466 source.n258 source.n231 12.0247
R467 source.n538 source.n537 11.249
R468 source.n555 source.n508 11.249
R469 source.n462 source.n461 11.249
R470 source.n479 source.n432 11.249
R471 source.n396 source.n395 11.249
R472 source.n413 source.n366 11.249
R473 source.n320 source.n319 11.249
R474 source.n337 source.n290 11.249
R475 source.n53 source.n6 11.249
R476 source.n37 source.n36 11.249
R477 source.n129 source.n82 11.249
R478 source.n113 source.n112 11.249
R479 source.n195 source.n148 11.249
R480 source.n179 source.n178 11.249
R481 source.n271 source.n224 11.249
R482 source.n255 source.n254 11.249
R483 source.n534 source.n516 10.4732
R484 source.n556 source.n506 10.4732
R485 source.n458 source.n440 10.4732
R486 source.n480 source.n430 10.4732
R487 source.n392 source.n374 10.4732
R488 source.n414 source.n364 10.4732
R489 source.n316 source.n298 10.4732
R490 source.n338 source.n288 10.4732
R491 source.n54 source.n4 10.4732
R492 source.n33 source.n15 10.4732
R493 source.n130 source.n80 10.4732
R494 source.n109 source.n91 10.4732
R495 source.n196 source.n146 10.4732
R496 source.n175 source.n157 10.4732
R497 source.n272 source.n222 10.4732
R498 source.n251 source.n233 10.4732
R499 source.n523 source.n522 10.2747
R500 source.n447 source.n446 10.2747
R501 source.n381 source.n380 10.2747
R502 source.n305 source.n304 10.2747
R503 source.n22 source.n21 10.2747
R504 source.n98 source.n97 10.2747
R505 source.n164 source.n163 10.2747
R506 source.n240 source.n239 10.2747
R507 source.n533 source.n518 9.69747
R508 source.n560 source.n559 9.69747
R509 source.n457 source.n442 9.69747
R510 source.n484 source.n483 9.69747
R511 source.n391 source.n376 9.69747
R512 source.n418 source.n417 9.69747
R513 source.n315 source.n300 9.69747
R514 source.n342 source.n341 9.69747
R515 source.n58 source.n57 9.69747
R516 source.n32 source.n17 9.69747
R517 source.n134 source.n133 9.69747
R518 source.n108 source.n93 9.69747
R519 source.n200 source.n199 9.69747
R520 source.n174 source.n159 9.69747
R521 source.n276 source.n275 9.69747
R522 source.n250 source.n235 9.69747
R523 source.n566 source.n565 9.45567
R524 source.n490 source.n489 9.45567
R525 source.n424 source.n423 9.45567
R526 source.n348 source.n347 9.45567
R527 source.n64 source.n63 9.45567
R528 source.n140 source.n139 9.45567
R529 source.n206 source.n205 9.45567
R530 source.n282 source.n281 9.45567
R531 source.n565 source.n564 9.3005
R532 source.n504 source.n503 9.3005
R533 source.n559 source.n558 9.3005
R534 source.n557 source.n556 9.3005
R535 source.n508 source.n507 9.3005
R536 source.n551 source.n550 9.3005
R537 source.n549 source.n548 9.3005
R538 source.n525 source.n524 9.3005
R539 source.n520 source.n519 9.3005
R540 source.n531 source.n530 9.3005
R541 source.n533 source.n532 9.3005
R542 source.n516 source.n515 9.3005
R543 source.n539 source.n538 9.3005
R544 source.n541 source.n540 9.3005
R545 source.n542 source.n511 9.3005
R546 source.n489 source.n488 9.3005
R547 source.n428 source.n427 9.3005
R548 source.n483 source.n482 9.3005
R549 source.n481 source.n480 9.3005
R550 source.n432 source.n431 9.3005
R551 source.n475 source.n474 9.3005
R552 source.n473 source.n472 9.3005
R553 source.n449 source.n448 9.3005
R554 source.n444 source.n443 9.3005
R555 source.n455 source.n454 9.3005
R556 source.n457 source.n456 9.3005
R557 source.n440 source.n439 9.3005
R558 source.n463 source.n462 9.3005
R559 source.n465 source.n464 9.3005
R560 source.n466 source.n435 9.3005
R561 source.n423 source.n422 9.3005
R562 source.n362 source.n361 9.3005
R563 source.n417 source.n416 9.3005
R564 source.n415 source.n414 9.3005
R565 source.n366 source.n365 9.3005
R566 source.n409 source.n408 9.3005
R567 source.n407 source.n406 9.3005
R568 source.n383 source.n382 9.3005
R569 source.n378 source.n377 9.3005
R570 source.n389 source.n388 9.3005
R571 source.n391 source.n390 9.3005
R572 source.n374 source.n373 9.3005
R573 source.n397 source.n396 9.3005
R574 source.n399 source.n398 9.3005
R575 source.n400 source.n369 9.3005
R576 source.n347 source.n346 9.3005
R577 source.n286 source.n285 9.3005
R578 source.n341 source.n340 9.3005
R579 source.n339 source.n338 9.3005
R580 source.n290 source.n289 9.3005
R581 source.n333 source.n332 9.3005
R582 source.n331 source.n330 9.3005
R583 source.n307 source.n306 9.3005
R584 source.n302 source.n301 9.3005
R585 source.n313 source.n312 9.3005
R586 source.n315 source.n314 9.3005
R587 source.n298 source.n297 9.3005
R588 source.n321 source.n320 9.3005
R589 source.n323 source.n322 9.3005
R590 source.n324 source.n293 9.3005
R591 source.n24 source.n23 9.3005
R592 source.n19 source.n18 9.3005
R593 source.n30 source.n29 9.3005
R594 source.n32 source.n31 9.3005
R595 source.n15 source.n14 9.3005
R596 source.n38 source.n37 9.3005
R597 source.n40 source.n39 9.3005
R598 source.n12 source.n9 9.3005
R599 source.n63 source.n62 9.3005
R600 source.n2 source.n1 9.3005
R601 source.n57 source.n56 9.3005
R602 source.n55 source.n54 9.3005
R603 source.n6 source.n5 9.3005
R604 source.n49 source.n48 9.3005
R605 source.n47 source.n46 9.3005
R606 source.n100 source.n99 9.3005
R607 source.n95 source.n94 9.3005
R608 source.n106 source.n105 9.3005
R609 source.n108 source.n107 9.3005
R610 source.n91 source.n90 9.3005
R611 source.n114 source.n113 9.3005
R612 source.n116 source.n115 9.3005
R613 source.n88 source.n85 9.3005
R614 source.n139 source.n138 9.3005
R615 source.n78 source.n77 9.3005
R616 source.n133 source.n132 9.3005
R617 source.n131 source.n130 9.3005
R618 source.n82 source.n81 9.3005
R619 source.n125 source.n124 9.3005
R620 source.n123 source.n122 9.3005
R621 source.n166 source.n165 9.3005
R622 source.n161 source.n160 9.3005
R623 source.n172 source.n171 9.3005
R624 source.n174 source.n173 9.3005
R625 source.n157 source.n156 9.3005
R626 source.n180 source.n179 9.3005
R627 source.n182 source.n181 9.3005
R628 source.n154 source.n151 9.3005
R629 source.n205 source.n204 9.3005
R630 source.n144 source.n143 9.3005
R631 source.n199 source.n198 9.3005
R632 source.n197 source.n196 9.3005
R633 source.n148 source.n147 9.3005
R634 source.n191 source.n190 9.3005
R635 source.n189 source.n188 9.3005
R636 source.n242 source.n241 9.3005
R637 source.n237 source.n236 9.3005
R638 source.n248 source.n247 9.3005
R639 source.n250 source.n249 9.3005
R640 source.n233 source.n232 9.3005
R641 source.n256 source.n255 9.3005
R642 source.n258 source.n257 9.3005
R643 source.n230 source.n227 9.3005
R644 source.n281 source.n280 9.3005
R645 source.n220 source.n219 9.3005
R646 source.n275 source.n274 9.3005
R647 source.n273 source.n272 9.3005
R648 source.n224 source.n223 9.3005
R649 source.n267 source.n266 9.3005
R650 source.n265 source.n264 9.3005
R651 source.n530 source.n529 8.92171
R652 source.n563 source.n504 8.92171
R653 source.n454 source.n453 8.92171
R654 source.n487 source.n428 8.92171
R655 source.n388 source.n387 8.92171
R656 source.n421 source.n362 8.92171
R657 source.n312 source.n311 8.92171
R658 source.n345 source.n286 8.92171
R659 source.n61 source.n2 8.92171
R660 source.n29 source.n28 8.92171
R661 source.n137 source.n78 8.92171
R662 source.n105 source.n104 8.92171
R663 source.n203 source.n144 8.92171
R664 source.n171 source.n170 8.92171
R665 source.n279 source.n220 8.92171
R666 source.n247 source.n246 8.92171
R667 source.n526 source.n520 8.14595
R668 source.n564 source.n502 8.14595
R669 source.n450 source.n444 8.14595
R670 source.n488 source.n426 8.14595
R671 source.n384 source.n378 8.14595
R672 source.n422 source.n360 8.14595
R673 source.n308 source.n302 8.14595
R674 source.n346 source.n284 8.14595
R675 source.n62 source.n0 8.14595
R676 source.n25 source.n19 8.14595
R677 source.n138 source.n76 8.14595
R678 source.n101 source.n95 8.14595
R679 source.n204 source.n142 8.14595
R680 source.n167 source.n161 8.14595
R681 source.n280 source.n218 8.14595
R682 source.n243 source.n237 8.14595
R683 source.n525 source.n522 7.3702
R684 source.n449 source.n446 7.3702
R685 source.n383 source.n380 7.3702
R686 source.n307 source.n304 7.3702
R687 source.n24 source.n21 7.3702
R688 source.n100 source.n97 7.3702
R689 source.n166 source.n163 7.3702
R690 source.n242 source.n239 7.3702
R691 source.n526 source.n525 5.81868
R692 source.n566 source.n502 5.81868
R693 source.n450 source.n449 5.81868
R694 source.n490 source.n426 5.81868
R695 source.n384 source.n383 5.81868
R696 source.n424 source.n360 5.81868
R697 source.n308 source.n307 5.81868
R698 source.n348 source.n284 5.81868
R699 source.n64 source.n0 5.81868
R700 source.n25 source.n24 5.81868
R701 source.n140 source.n76 5.81868
R702 source.n101 source.n100 5.81868
R703 source.n206 source.n142 5.81868
R704 source.n167 source.n166 5.81868
R705 source.n282 source.n218 5.81868
R706 source.n243 source.n242 5.81868
R707 source.n568 source.n567 5.62119
R708 source.n529 source.n520 5.04292
R709 source.n564 source.n563 5.04292
R710 source.n453 source.n444 5.04292
R711 source.n488 source.n487 5.04292
R712 source.n387 source.n378 5.04292
R713 source.n422 source.n421 5.04292
R714 source.n311 source.n302 5.04292
R715 source.n346 source.n345 5.04292
R716 source.n62 source.n61 5.04292
R717 source.n28 source.n19 5.04292
R718 source.n138 source.n137 5.04292
R719 source.n104 source.n95 5.04292
R720 source.n204 source.n203 5.04292
R721 source.n170 source.n161 5.04292
R722 source.n280 source.n279 5.04292
R723 source.n246 source.n237 5.04292
R724 source.n530 source.n518 4.26717
R725 source.n560 source.n504 4.26717
R726 source.n454 source.n442 4.26717
R727 source.n484 source.n428 4.26717
R728 source.n388 source.n376 4.26717
R729 source.n418 source.n362 4.26717
R730 source.n312 source.n300 4.26717
R731 source.n342 source.n286 4.26717
R732 source.n58 source.n2 4.26717
R733 source.n29 source.n17 4.26717
R734 source.n134 source.n78 4.26717
R735 source.n105 source.n93 4.26717
R736 source.n200 source.n144 4.26717
R737 source.n171 source.n159 4.26717
R738 source.n276 source.n220 4.26717
R739 source.n247 source.n235 4.26717
R740 source.n534 source.n533 3.49141
R741 source.n559 source.n506 3.49141
R742 source.n458 source.n457 3.49141
R743 source.n483 source.n430 3.49141
R744 source.n392 source.n391 3.49141
R745 source.n417 source.n364 3.49141
R746 source.n316 source.n315 3.49141
R747 source.n341 source.n288 3.49141
R748 source.n57 source.n4 3.49141
R749 source.n33 source.n32 3.49141
R750 source.n133 source.n80 3.49141
R751 source.n109 source.n108 3.49141
R752 source.n199 source.n146 3.49141
R753 source.n175 source.n174 3.49141
R754 source.n275 source.n222 3.49141
R755 source.n251 source.n250 3.49141
R756 source.n524 source.n523 2.84303
R757 source.n448 source.n447 2.84303
R758 source.n382 source.n381 2.84303
R759 source.n306 source.n305 2.84303
R760 source.n23 source.n22 2.84303
R761 source.n99 source.n98 2.84303
R762 source.n165 source.n164 2.84303
R763 source.n241 source.n240 2.84303
R764 source.n537 source.n516 2.71565
R765 source.n556 source.n555 2.71565
R766 source.n461 source.n440 2.71565
R767 source.n480 source.n479 2.71565
R768 source.n395 source.n374 2.71565
R769 source.n414 source.n413 2.71565
R770 source.n319 source.n298 2.71565
R771 source.n338 source.n337 2.71565
R772 source.n54 source.n53 2.71565
R773 source.n36 source.n15 2.71565
R774 source.n130 source.n129 2.71565
R775 source.n112 source.n91 2.71565
R776 source.n196 source.n195 2.71565
R777 source.n178 source.n157 2.71565
R778 source.n272 source.n271 2.71565
R779 source.n254 source.n233 2.71565
R780 source.n538 source.n514 1.93989
R781 source.n552 source.n508 1.93989
R782 source.n462 source.n438 1.93989
R783 source.n476 source.n432 1.93989
R784 source.n396 source.n372 1.93989
R785 source.n410 source.n366 1.93989
R786 source.n320 source.n296 1.93989
R787 source.n334 source.n290 1.93989
R788 source.n50 source.n6 1.93989
R789 source.n37 source.n13 1.93989
R790 source.n126 source.n82 1.93989
R791 source.n113 source.n89 1.93989
R792 source.n192 source.n148 1.93989
R793 source.n179 source.n155 1.93989
R794 source.n268 source.n224 1.93989
R795 source.n255 source.n231 1.93989
R796 source.n500 source.t41 1.6505
R797 source.n500 source.t27 1.6505
R798 source.n498 source.t25 1.6505
R799 source.n498 source.t44 1.6505
R800 source.n496 source.t35 1.6505
R801 source.n496 source.t34 1.6505
R802 source.n494 source.t39 1.6505
R803 source.n494 source.t30 1.6505
R804 source.n492 source.t45 1.6505
R805 source.n492 source.t38 1.6505
R806 source.n358 source.t46 1.6505
R807 source.n358 source.t9 1.6505
R808 source.n356 source.t10 1.6505
R809 source.n356 source.t3 1.6505
R810 source.n354 source.t11 1.6505
R811 source.n354 source.t4 1.6505
R812 source.n352 source.t47 1.6505
R813 source.n352 source.t1 1.6505
R814 source.n350 source.t13 1.6505
R815 source.n350 source.t5 1.6505
R816 source.n66 source.t18 1.6505
R817 source.n66 source.t6 1.6505
R818 source.n68 source.t21 1.6505
R819 source.n68 source.t19 1.6505
R820 source.n70 source.t16 1.6505
R821 source.n70 source.t20 1.6505
R822 source.n72 source.t0 1.6505
R823 source.n72 source.t17 1.6505
R824 source.n74 source.t8 1.6505
R825 source.n74 source.t15 1.6505
R826 source.n208 source.t37 1.6505
R827 source.n208 source.t43 1.6505
R828 source.n210 source.t29 1.6505
R829 source.n210 source.t32 1.6505
R830 source.n212 source.t22 1.6505
R831 source.n212 source.t40 1.6505
R832 source.n214 source.t24 1.6505
R833 source.n214 source.t23 1.6505
R834 source.n216 source.t26 1.6505
R835 source.n216 source.t42 1.6505
R836 source.n543 source.n541 1.16414
R837 source.n551 source.n510 1.16414
R838 source.n467 source.n465 1.16414
R839 source.n475 source.n434 1.16414
R840 source.n401 source.n399 1.16414
R841 source.n409 source.n368 1.16414
R842 source.n325 source.n323 1.16414
R843 source.n333 source.n292 1.16414
R844 source.n49 source.n8 1.16414
R845 source.n41 source.n40 1.16414
R846 source.n125 source.n84 1.16414
R847 source.n117 source.n116 1.16414
R848 source.n191 source.n150 1.16414
R849 source.n183 source.n182 1.16414
R850 source.n267 source.n226 1.16414
R851 source.n259 source.n258 1.16414
R852 source.n283 source.n217 0.716017
R853 source.n217 source.n215 0.716017
R854 source.n215 source.n213 0.716017
R855 source.n213 source.n211 0.716017
R856 source.n211 source.n209 0.716017
R857 source.n209 source.n207 0.716017
R858 source.n141 source.n75 0.716017
R859 source.n75 source.n73 0.716017
R860 source.n73 source.n71 0.716017
R861 source.n71 source.n69 0.716017
R862 source.n69 source.n67 0.716017
R863 source.n67 source.n65 0.716017
R864 source.n351 source.n349 0.716017
R865 source.n353 source.n351 0.716017
R866 source.n355 source.n353 0.716017
R867 source.n357 source.n355 0.716017
R868 source.n359 source.n357 0.716017
R869 source.n425 source.n359 0.716017
R870 source.n493 source.n491 0.716017
R871 source.n495 source.n493 0.716017
R872 source.n497 source.n495 0.716017
R873 source.n499 source.n497 0.716017
R874 source.n501 source.n499 0.716017
R875 source.n567 source.n501 0.716017
R876 source.n207 source.n141 0.470328
R877 source.n491 source.n425 0.470328
R878 source.n542 source.n512 0.388379
R879 source.n548 source.n547 0.388379
R880 source.n466 source.n436 0.388379
R881 source.n472 source.n471 0.388379
R882 source.n400 source.n370 0.388379
R883 source.n406 source.n405 0.388379
R884 source.n324 source.n294 0.388379
R885 source.n330 source.n329 0.388379
R886 source.n46 source.n45 0.388379
R887 source.n12 source.n10 0.388379
R888 source.n122 source.n121 0.388379
R889 source.n88 source.n86 0.388379
R890 source.n188 source.n187 0.388379
R891 source.n154 source.n152 0.388379
R892 source.n264 source.n263 0.388379
R893 source.n230 source.n228 0.388379
R894 source source.n568 0.188
R895 source.n524 source.n519 0.155672
R896 source.n531 source.n519 0.155672
R897 source.n532 source.n531 0.155672
R898 source.n532 source.n515 0.155672
R899 source.n539 source.n515 0.155672
R900 source.n540 source.n539 0.155672
R901 source.n540 source.n511 0.155672
R902 source.n549 source.n511 0.155672
R903 source.n550 source.n549 0.155672
R904 source.n550 source.n507 0.155672
R905 source.n557 source.n507 0.155672
R906 source.n558 source.n557 0.155672
R907 source.n558 source.n503 0.155672
R908 source.n565 source.n503 0.155672
R909 source.n448 source.n443 0.155672
R910 source.n455 source.n443 0.155672
R911 source.n456 source.n455 0.155672
R912 source.n456 source.n439 0.155672
R913 source.n463 source.n439 0.155672
R914 source.n464 source.n463 0.155672
R915 source.n464 source.n435 0.155672
R916 source.n473 source.n435 0.155672
R917 source.n474 source.n473 0.155672
R918 source.n474 source.n431 0.155672
R919 source.n481 source.n431 0.155672
R920 source.n482 source.n481 0.155672
R921 source.n482 source.n427 0.155672
R922 source.n489 source.n427 0.155672
R923 source.n382 source.n377 0.155672
R924 source.n389 source.n377 0.155672
R925 source.n390 source.n389 0.155672
R926 source.n390 source.n373 0.155672
R927 source.n397 source.n373 0.155672
R928 source.n398 source.n397 0.155672
R929 source.n398 source.n369 0.155672
R930 source.n407 source.n369 0.155672
R931 source.n408 source.n407 0.155672
R932 source.n408 source.n365 0.155672
R933 source.n415 source.n365 0.155672
R934 source.n416 source.n415 0.155672
R935 source.n416 source.n361 0.155672
R936 source.n423 source.n361 0.155672
R937 source.n306 source.n301 0.155672
R938 source.n313 source.n301 0.155672
R939 source.n314 source.n313 0.155672
R940 source.n314 source.n297 0.155672
R941 source.n321 source.n297 0.155672
R942 source.n322 source.n321 0.155672
R943 source.n322 source.n293 0.155672
R944 source.n331 source.n293 0.155672
R945 source.n332 source.n331 0.155672
R946 source.n332 source.n289 0.155672
R947 source.n339 source.n289 0.155672
R948 source.n340 source.n339 0.155672
R949 source.n340 source.n285 0.155672
R950 source.n347 source.n285 0.155672
R951 source.n63 source.n1 0.155672
R952 source.n56 source.n1 0.155672
R953 source.n56 source.n55 0.155672
R954 source.n55 source.n5 0.155672
R955 source.n48 source.n5 0.155672
R956 source.n48 source.n47 0.155672
R957 source.n47 source.n9 0.155672
R958 source.n39 source.n9 0.155672
R959 source.n39 source.n38 0.155672
R960 source.n38 source.n14 0.155672
R961 source.n31 source.n14 0.155672
R962 source.n31 source.n30 0.155672
R963 source.n30 source.n18 0.155672
R964 source.n23 source.n18 0.155672
R965 source.n139 source.n77 0.155672
R966 source.n132 source.n77 0.155672
R967 source.n132 source.n131 0.155672
R968 source.n131 source.n81 0.155672
R969 source.n124 source.n81 0.155672
R970 source.n124 source.n123 0.155672
R971 source.n123 source.n85 0.155672
R972 source.n115 source.n85 0.155672
R973 source.n115 source.n114 0.155672
R974 source.n114 source.n90 0.155672
R975 source.n107 source.n90 0.155672
R976 source.n107 source.n106 0.155672
R977 source.n106 source.n94 0.155672
R978 source.n99 source.n94 0.155672
R979 source.n205 source.n143 0.155672
R980 source.n198 source.n143 0.155672
R981 source.n198 source.n197 0.155672
R982 source.n197 source.n147 0.155672
R983 source.n190 source.n147 0.155672
R984 source.n190 source.n189 0.155672
R985 source.n189 source.n151 0.155672
R986 source.n181 source.n151 0.155672
R987 source.n181 source.n180 0.155672
R988 source.n180 source.n156 0.155672
R989 source.n173 source.n156 0.155672
R990 source.n173 source.n172 0.155672
R991 source.n172 source.n160 0.155672
R992 source.n165 source.n160 0.155672
R993 source.n281 source.n219 0.155672
R994 source.n274 source.n219 0.155672
R995 source.n274 source.n273 0.155672
R996 source.n273 source.n223 0.155672
R997 source.n266 source.n223 0.155672
R998 source.n266 source.n265 0.155672
R999 source.n265 source.n227 0.155672
R1000 source.n257 source.n227 0.155672
R1001 source.n257 source.n256 0.155672
R1002 source.n256 source.n232 0.155672
R1003 source.n249 source.n232 0.155672
R1004 source.n249 source.n248 0.155672
R1005 source.n248 source.n236 0.155672
R1006 source.n241 source.n236 0.155672
R1007 drain_right.n7 drain_right.n5 60.268
R1008 drain_right.n2 drain_right.n0 60.268
R1009 drain_right.n13 drain_right.n11 60.268
R1010 drain_right.n13 drain_right.n12 59.5527
R1011 drain_right.n15 drain_right.n14 59.5527
R1012 drain_right.n17 drain_right.n16 59.5527
R1013 drain_right.n19 drain_right.n18 59.5527
R1014 drain_right.n21 drain_right.n20 59.5527
R1015 drain_right.n7 drain_right.n6 59.5525
R1016 drain_right.n9 drain_right.n8 59.5525
R1017 drain_right.n4 drain_right.n3 59.5525
R1018 drain_right.n2 drain_right.n1 59.5525
R1019 drain_right drain_right.n10 33.6113
R1020 drain_right drain_right.n21 6.36873
R1021 drain_right.n5 drain_right.t13 1.6505
R1022 drain_right.n5 drain_right.t23 1.6505
R1023 drain_right.n6 drain_right.t0 1.6505
R1024 drain_right.n6 drain_right.t3 1.6505
R1025 drain_right.n8 drain_right.t8 1.6505
R1026 drain_right.n8 drain_right.t14 1.6505
R1027 drain_right.n3 drain_right.t17 1.6505
R1028 drain_right.n3 drain_right.t7 1.6505
R1029 drain_right.n1 drain_right.t11 1.6505
R1030 drain_right.n1 drain_right.t12 1.6505
R1031 drain_right.n0 drain_right.t20 1.6505
R1032 drain_right.n0 drain_right.t21 1.6505
R1033 drain_right.n11 drain_right.t19 1.6505
R1034 drain_right.n11 drain_right.t6 1.6505
R1035 drain_right.n12 drain_right.t2 1.6505
R1036 drain_right.n12 drain_right.t15 1.6505
R1037 drain_right.n14 drain_right.t10 1.6505
R1038 drain_right.n14 drain_right.t16 1.6505
R1039 drain_right.n16 drain_right.t9 1.6505
R1040 drain_right.n16 drain_right.t22 1.6505
R1041 drain_right.n18 drain_right.t18 1.6505
R1042 drain_right.n18 drain_right.t4 1.6505
R1043 drain_right.n20 drain_right.t1 1.6505
R1044 drain_right.n20 drain_right.t5 1.6505
R1045 drain_right.n9 drain_right.n7 0.716017
R1046 drain_right.n4 drain_right.n2 0.716017
R1047 drain_right.n21 drain_right.n19 0.716017
R1048 drain_right.n19 drain_right.n17 0.716017
R1049 drain_right.n17 drain_right.n15 0.716017
R1050 drain_right.n15 drain_right.n13 0.716017
R1051 drain_right.n10 drain_right.n9 0.302913
R1052 drain_right.n10 drain_right.n4 0.302913
R1053 plus.n11 plus.t6 683.324
R1054 plus.n45 plus.t18 683.324
R1055 plus.n32 plus.t2 656.966
R1056 plus.n30 plus.t3 656.966
R1057 plus.n29 plus.t14 656.966
R1058 plus.n3 plus.t5 656.966
R1059 plus.n23 plus.t20 656.966
R1060 plus.n22 plus.t13 656.966
R1061 plus.n6 plus.t23 656.966
R1062 plus.n17 plus.t17 656.966
R1063 plus.n15 plus.t11 656.966
R1064 plus.n9 plus.t21 656.966
R1065 plus.n10 plus.t15 656.966
R1066 plus.n66 plus.t16 656.966
R1067 plus.n64 plus.t4 656.966
R1068 plus.n63 plus.t10 656.966
R1069 plus.n37 plus.t9 656.966
R1070 plus.n57 plus.t22 656.966
R1071 plus.n56 plus.t7 656.966
R1072 plus.n40 plus.t12 656.966
R1073 plus.n51 plus.t1 656.966
R1074 plus.n49 plus.t0 656.966
R1075 plus.n43 plus.t8 656.966
R1076 plus.n44 plus.t19 656.966
R1077 plus.n12 plus.n9 161.3
R1078 plus.n14 plus.n13 161.3
R1079 plus.n15 plus.n8 161.3
R1080 plus.n16 plus.n7 161.3
R1081 plus.n18 plus.n17 161.3
R1082 plus.n19 plus.n6 161.3
R1083 plus.n21 plus.n20 161.3
R1084 plus.n22 plus.n5 161.3
R1085 plus.n23 plus.n4 161.3
R1086 plus.n25 plus.n24 161.3
R1087 plus.n26 plus.n3 161.3
R1088 plus.n28 plus.n27 161.3
R1089 plus.n29 plus.n2 161.3
R1090 plus.n30 plus.n1 161.3
R1091 plus.n31 plus.n0 161.3
R1092 plus.n33 plus.n32 161.3
R1093 plus.n46 plus.n43 161.3
R1094 plus.n48 plus.n47 161.3
R1095 plus.n49 plus.n42 161.3
R1096 plus.n50 plus.n41 161.3
R1097 plus.n52 plus.n51 161.3
R1098 plus.n53 plus.n40 161.3
R1099 plus.n55 plus.n54 161.3
R1100 plus.n56 plus.n39 161.3
R1101 plus.n57 plus.n38 161.3
R1102 plus.n59 plus.n58 161.3
R1103 plus.n60 plus.n37 161.3
R1104 plus.n62 plus.n61 161.3
R1105 plus.n63 plus.n36 161.3
R1106 plus.n64 plus.n35 161.3
R1107 plus.n65 plus.n34 161.3
R1108 plus.n67 plus.n66 161.3
R1109 plus.n30 plus.n29 48.2005
R1110 plus.n23 plus.n22 48.2005
R1111 plus.n17 plus.n6 48.2005
R1112 plus.n10 plus.n9 48.2005
R1113 plus.n64 plus.n63 48.2005
R1114 plus.n57 plus.n56 48.2005
R1115 plus.n51 plus.n40 48.2005
R1116 plus.n44 plus.n43 48.2005
R1117 plus.n24 plus.n3 47.4702
R1118 plus.n16 plus.n15 47.4702
R1119 plus.n58 plus.n37 47.4702
R1120 plus.n50 plus.n49 47.4702
R1121 plus.n32 plus.n31 46.0096
R1122 plus.n66 plus.n65 46.0096
R1123 plus.n12 plus.n11 45.0871
R1124 plus.n46 plus.n45 45.0871
R1125 plus plus.n67 33.9157
R1126 plus.n28 plus.n3 25.5611
R1127 plus.n15 plus.n14 25.5611
R1128 plus.n62 plus.n37 25.5611
R1129 plus.n49 plus.n48 25.5611
R1130 plus.n21 plus.n6 24.1005
R1131 plus.n22 plus.n21 24.1005
R1132 plus.n56 plus.n55 24.1005
R1133 plus.n55 plus.n40 24.1005
R1134 plus.n29 plus.n28 22.6399
R1135 plus.n14 plus.n9 22.6399
R1136 plus.n63 plus.n62 22.6399
R1137 plus.n48 plus.n43 22.6399
R1138 plus.n11 plus.n10 14.1472
R1139 plus.n45 plus.n44 14.1472
R1140 plus plus.n33 12.171
R1141 plus.n31 plus.n30 2.19141
R1142 plus.n65 plus.n64 2.19141
R1143 plus.n24 plus.n23 0.730803
R1144 plus.n17 plus.n16 0.730803
R1145 plus.n58 plus.n57 0.730803
R1146 plus.n51 plus.n50 0.730803
R1147 plus.n13 plus.n12 0.189894
R1148 plus.n13 plus.n8 0.189894
R1149 plus.n8 plus.n7 0.189894
R1150 plus.n18 plus.n7 0.189894
R1151 plus.n19 plus.n18 0.189894
R1152 plus.n20 plus.n19 0.189894
R1153 plus.n20 plus.n5 0.189894
R1154 plus.n5 plus.n4 0.189894
R1155 plus.n25 plus.n4 0.189894
R1156 plus.n26 plus.n25 0.189894
R1157 plus.n27 plus.n26 0.189894
R1158 plus.n27 plus.n2 0.189894
R1159 plus.n2 plus.n1 0.189894
R1160 plus.n1 plus.n0 0.189894
R1161 plus.n33 plus.n0 0.189894
R1162 plus.n67 plus.n34 0.189894
R1163 plus.n35 plus.n34 0.189894
R1164 plus.n36 plus.n35 0.189894
R1165 plus.n61 plus.n36 0.189894
R1166 plus.n61 plus.n60 0.189894
R1167 plus.n60 plus.n59 0.189894
R1168 plus.n59 plus.n38 0.189894
R1169 plus.n39 plus.n38 0.189894
R1170 plus.n54 plus.n39 0.189894
R1171 plus.n54 plus.n53 0.189894
R1172 plus.n53 plus.n52 0.189894
R1173 plus.n52 plus.n41 0.189894
R1174 plus.n42 plus.n41 0.189894
R1175 plus.n47 plus.n42 0.189894
R1176 plus.n47 plus.n46 0.189894
R1177 drain_left.n13 drain_left.n11 60.2682
R1178 drain_left.n7 drain_left.n5 60.268
R1179 drain_left.n2 drain_left.n0 60.268
R1180 drain_left.n19 drain_left.n18 59.5527
R1181 drain_left.n17 drain_left.n16 59.5527
R1182 drain_left.n15 drain_left.n14 59.5527
R1183 drain_left.n13 drain_left.n12 59.5527
R1184 drain_left.n7 drain_left.n6 59.5525
R1185 drain_left.n9 drain_left.n8 59.5525
R1186 drain_left.n4 drain_left.n3 59.5525
R1187 drain_left.n2 drain_left.n1 59.5525
R1188 drain_left.n21 drain_left.n20 59.5525
R1189 drain_left drain_left.n10 34.1645
R1190 drain_left drain_left.n21 6.36873
R1191 drain_left.n5 drain_left.t4 1.6505
R1192 drain_left.n5 drain_left.t5 1.6505
R1193 drain_left.n6 drain_left.t23 1.6505
R1194 drain_left.n6 drain_left.t15 1.6505
R1195 drain_left.n8 drain_left.t11 1.6505
R1196 drain_left.n8 drain_left.t22 1.6505
R1197 drain_left.n3 drain_left.t1 1.6505
R1198 drain_left.n3 drain_left.t16 1.6505
R1199 drain_left.n1 drain_left.t13 1.6505
R1200 drain_left.n1 drain_left.t14 1.6505
R1201 drain_left.n0 drain_left.t7 1.6505
R1202 drain_left.n0 drain_left.t19 1.6505
R1203 drain_left.n20 drain_left.t20 1.6505
R1204 drain_left.n20 drain_left.t21 1.6505
R1205 drain_left.n18 drain_left.t18 1.6505
R1206 drain_left.n18 drain_left.t9 1.6505
R1207 drain_left.n16 drain_left.t10 1.6505
R1208 drain_left.n16 drain_left.t3 1.6505
R1209 drain_left.n14 drain_left.t6 1.6505
R1210 drain_left.n14 drain_left.t0 1.6505
R1211 drain_left.n12 drain_left.t2 1.6505
R1212 drain_left.n12 drain_left.t12 1.6505
R1213 drain_left.n11 drain_left.t17 1.6505
R1214 drain_left.n11 drain_left.t8 1.6505
R1215 drain_left.n9 drain_left.n7 0.716017
R1216 drain_left.n4 drain_left.n2 0.716017
R1217 drain_left.n15 drain_left.n13 0.716017
R1218 drain_left.n17 drain_left.n15 0.716017
R1219 drain_left.n19 drain_left.n17 0.716017
R1220 drain_left.n21 drain_left.n19 0.716017
R1221 drain_left.n10 drain_left.n9 0.302913
R1222 drain_left.n10 drain_left.n4 0.302913
C0 plus minus 6.74153f
C1 drain_right plus 0.443411f
C2 minus source 12.190701f
C3 drain_right source 33.9729f
C4 minus drain_left 0.173624f
C5 drain_right drain_left 1.55979f
C6 plus source 12.2047f
C7 plus drain_left 12.4201f
C8 source drain_left 33.9713f
C9 drain_right minus 12.1337f
C10 drain_right a_n2874_n3288# 7.5204f
C11 drain_left a_n2874_n3288# 7.93102f
C12 source a_n2874_n3288# 9.277133f
C13 minus a_n2874_n3288# 11.520677f
C14 plus a_n2874_n3288# 13.48404f
C15 drain_left.t7 a_n2874_n3288# 0.279702f
C16 drain_left.t19 a_n2874_n3288# 0.279702f
C17 drain_left.n0 a_n2874_n3288# 2.49361f
C18 drain_left.t13 a_n2874_n3288# 0.279702f
C19 drain_left.t14 a_n2874_n3288# 0.279702f
C20 drain_left.n1 a_n2874_n3288# 2.48891f
C21 drain_left.n2 a_n2874_n3288# 0.774293f
C22 drain_left.t1 a_n2874_n3288# 0.279702f
C23 drain_left.t16 a_n2874_n3288# 0.279702f
C24 drain_left.n3 a_n2874_n3288# 2.48891f
C25 drain_left.n4 a_n2874_n3288# 0.346553f
C26 drain_left.t4 a_n2874_n3288# 0.279702f
C27 drain_left.t5 a_n2874_n3288# 0.279702f
C28 drain_left.n5 a_n2874_n3288# 2.49361f
C29 drain_left.t23 a_n2874_n3288# 0.279702f
C30 drain_left.t15 a_n2874_n3288# 0.279702f
C31 drain_left.n6 a_n2874_n3288# 2.48891f
C32 drain_left.n7 a_n2874_n3288# 0.774293f
C33 drain_left.t11 a_n2874_n3288# 0.279702f
C34 drain_left.t22 a_n2874_n3288# 0.279702f
C35 drain_left.n8 a_n2874_n3288# 2.48891f
C36 drain_left.n9 a_n2874_n3288# 0.346553f
C37 drain_left.n10 a_n2874_n3288# 1.77374f
C38 drain_left.t17 a_n2874_n3288# 0.279702f
C39 drain_left.t8 a_n2874_n3288# 0.279702f
C40 drain_left.n11 a_n2874_n3288# 2.49362f
C41 drain_left.t2 a_n2874_n3288# 0.279702f
C42 drain_left.t12 a_n2874_n3288# 0.279702f
C43 drain_left.n12 a_n2874_n3288# 2.48892f
C44 drain_left.n13 a_n2874_n3288# 0.774273f
C45 drain_left.t6 a_n2874_n3288# 0.279702f
C46 drain_left.t0 a_n2874_n3288# 0.279702f
C47 drain_left.n14 a_n2874_n3288# 2.48892f
C48 drain_left.n15 a_n2874_n3288# 0.383544f
C49 drain_left.t10 a_n2874_n3288# 0.279702f
C50 drain_left.t3 a_n2874_n3288# 0.279702f
C51 drain_left.n16 a_n2874_n3288# 2.48892f
C52 drain_left.n17 a_n2874_n3288# 0.383544f
C53 drain_left.t18 a_n2874_n3288# 0.279702f
C54 drain_left.t9 a_n2874_n3288# 0.279702f
C55 drain_left.n18 a_n2874_n3288# 2.48892f
C56 drain_left.n19 a_n2874_n3288# 0.383544f
C57 drain_left.t20 a_n2874_n3288# 0.279702f
C58 drain_left.t21 a_n2874_n3288# 0.279702f
C59 drain_left.n20 a_n2874_n3288# 2.48891f
C60 drain_left.n21 a_n2874_n3288# 0.636964f
C61 plus.n0 a_n2874_n3288# 0.043909f
C62 plus.t2 a_n2874_n3288# 0.751235f
C63 plus.t3 a_n2874_n3288# 0.751235f
C64 plus.n1 a_n2874_n3288# 0.043909f
C65 plus.t14 a_n2874_n3288# 0.751235f
C66 plus.n2 a_n2874_n3288# 0.043909f
C67 plus.t5 a_n2874_n3288# 0.751235f
C68 plus.n3 a_n2874_n3288# 0.307636f
C69 plus.n4 a_n2874_n3288# 0.043909f
C70 plus.t20 a_n2874_n3288# 0.751235f
C71 plus.t13 a_n2874_n3288# 0.751235f
C72 plus.n5 a_n2874_n3288# 0.043909f
C73 plus.t23 a_n2874_n3288# 0.751235f
C74 plus.n6 a_n2874_n3288# 0.3075f
C75 plus.n7 a_n2874_n3288# 0.043909f
C76 plus.t17 a_n2874_n3288# 0.751235f
C77 plus.t11 a_n2874_n3288# 0.751235f
C78 plus.n8 a_n2874_n3288# 0.043909f
C79 plus.t21 a_n2874_n3288# 0.751235f
C80 plus.n9 a_n2874_n3288# 0.30723f
C81 plus.t15 a_n2874_n3288# 0.751235f
C82 plus.n10 a_n2874_n3288# 0.312425f
C83 plus.t6 a_n2874_n3288# 0.762922f
C84 plus.n11 a_n2874_n3288# 0.292786f
C85 plus.n12 a_n2874_n3288# 0.178287f
C86 plus.n13 a_n2874_n3288# 0.043909f
C87 plus.n14 a_n2874_n3288# 0.009964f
C88 plus.n15 a_n2874_n3288# 0.307636f
C89 plus.n16 a_n2874_n3288# 0.009964f
C90 plus.n17 a_n2874_n3288# 0.303169f
C91 plus.n18 a_n2874_n3288# 0.043909f
C92 plus.n19 a_n2874_n3288# 0.043909f
C93 plus.n20 a_n2874_n3288# 0.043909f
C94 plus.n21 a_n2874_n3288# 0.009964f
C95 plus.n22 a_n2874_n3288# 0.3075f
C96 plus.n23 a_n2874_n3288# 0.303169f
C97 plus.n24 a_n2874_n3288# 0.009964f
C98 plus.n25 a_n2874_n3288# 0.043909f
C99 plus.n26 a_n2874_n3288# 0.043909f
C100 plus.n27 a_n2874_n3288# 0.043909f
C101 plus.n28 a_n2874_n3288# 0.009964f
C102 plus.n29 a_n2874_n3288# 0.30723f
C103 plus.n30 a_n2874_n3288# 0.30344f
C104 plus.n31 a_n2874_n3288# 0.009964f
C105 plus.n32 a_n2874_n3288# 0.302628f
C106 plus.n33 a_n2874_n3288# 0.494105f
C107 plus.n34 a_n2874_n3288# 0.043909f
C108 plus.t16 a_n2874_n3288# 0.751235f
C109 plus.n35 a_n2874_n3288# 0.043909f
C110 plus.t4 a_n2874_n3288# 0.751235f
C111 plus.n36 a_n2874_n3288# 0.043909f
C112 plus.t10 a_n2874_n3288# 0.751235f
C113 plus.t9 a_n2874_n3288# 0.751235f
C114 plus.n37 a_n2874_n3288# 0.307636f
C115 plus.n38 a_n2874_n3288# 0.043909f
C116 plus.t22 a_n2874_n3288# 0.751235f
C117 plus.n39 a_n2874_n3288# 0.043909f
C118 plus.t7 a_n2874_n3288# 0.751235f
C119 plus.t12 a_n2874_n3288# 0.751235f
C120 plus.n40 a_n2874_n3288# 0.3075f
C121 plus.n41 a_n2874_n3288# 0.043909f
C122 plus.t1 a_n2874_n3288# 0.751235f
C123 plus.n42 a_n2874_n3288# 0.043909f
C124 plus.t0 a_n2874_n3288# 0.751235f
C125 plus.t8 a_n2874_n3288# 0.751235f
C126 plus.n43 a_n2874_n3288# 0.30723f
C127 plus.t18 a_n2874_n3288# 0.762922f
C128 plus.t19 a_n2874_n3288# 0.751235f
C129 plus.n44 a_n2874_n3288# 0.312425f
C130 plus.n45 a_n2874_n3288# 0.292786f
C131 plus.n46 a_n2874_n3288# 0.178287f
C132 plus.n47 a_n2874_n3288# 0.043909f
C133 plus.n48 a_n2874_n3288# 0.009964f
C134 plus.n49 a_n2874_n3288# 0.307636f
C135 plus.n50 a_n2874_n3288# 0.009964f
C136 plus.n51 a_n2874_n3288# 0.303169f
C137 plus.n52 a_n2874_n3288# 0.043909f
C138 plus.n53 a_n2874_n3288# 0.043909f
C139 plus.n54 a_n2874_n3288# 0.043909f
C140 plus.n55 a_n2874_n3288# 0.009964f
C141 plus.n56 a_n2874_n3288# 0.3075f
C142 plus.n57 a_n2874_n3288# 0.303169f
C143 plus.n58 a_n2874_n3288# 0.009964f
C144 plus.n59 a_n2874_n3288# 0.043909f
C145 plus.n60 a_n2874_n3288# 0.043909f
C146 plus.n61 a_n2874_n3288# 0.043909f
C147 plus.n62 a_n2874_n3288# 0.009964f
C148 plus.n63 a_n2874_n3288# 0.30723f
C149 plus.n64 a_n2874_n3288# 0.30344f
C150 plus.n65 a_n2874_n3288# 0.009964f
C151 plus.n66 a_n2874_n3288# 0.302628f
C152 plus.n67 a_n2874_n3288# 1.54726f
C153 drain_right.t20 a_n2874_n3288# 0.278586f
C154 drain_right.t21 a_n2874_n3288# 0.278586f
C155 drain_right.n0 a_n2874_n3288# 2.48366f
C156 drain_right.t11 a_n2874_n3288# 0.278586f
C157 drain_right.t12 a_n2874_n3288# 0.278586f
C158 drain_right.n1 a_n2874_n3288# 2.47899f
C159 drain_right.n2 a_n2874_n3288# 0.771205f
C160 drain_right.t17 a_n2874_n3288# 0.278586f
C161 drain_right.t7 a_n2874_n3288# 0.278586f
C162 drain_right.n3 a_n2874_n3288# 2.47899f
C163 drain_right.n4 a_n2874_n3288# 0.34517f
C164 drain_right.t13 a_n2874_n3288# 0.278586f
C165 drain_right.t23 a_n2874_n3288# 0.278586f
C166 drain_right.n5 a_n2874_n3288# 2.48366f
C167 drain_right.t0 a_n2874_n3288# 0.278586f
C168 drain_right.t3 a_n2874_n3288# 0.278586f
C169 drain_right.n6 a_n2874_n3288# 2.47899f
C170 drain_right.n7 a_n2874_n3288# 0.771205f
C171 drain_right.t8 a_n2874_n3288# 0.278586f
C172 drain_right.t14 a_n2874_n3288# 0.278586f
C173 drain_right.n8 a_n2874_n3288# 2.47899f
C174 drain_right.n9 a_n2874_n3288# 0.34517f
C175 drain_right.n10 a_n2874_n3288# 1.70674f
C176 drain_right.t19 a_n2874_n3288# 0.278586f
C177 drain_right.t6 a_n2874_n3288# 0.278586f
C178 drain_right.n11 a_n2874_n3288# 2.48366f
C179 drain_right.t2 a_n2874_n3288# 0.278586f
C180 drain_right.t15 a_n2874_n3288# 0.278586f
C181 drain_right.n12 a_n2874_n3288# 2.479f
C182 drain_right.n13 a_n2874_n3288# 0.771195f
C183 drain_right.t10 a_n2874_n3288# 0.278586f
C184 drain_right.t16 a_n2874_n3288# 0.278586f
C185 drain_right.n14 a_n2874_n3288# 2.479f
C186 drain_right.n15 a_n2874_n3288# 0.382014f
C187 drain_right.t9 a_n2874_n3288# 0.278586f
C188 drain_right.t22 a_n2874_n3288# 0.278586f
C189 drain_right.n16 a_n2874_n3288# 2.479f
C190 drain_right.n17 a_n2874_n3288# 0.382014f
C191 drain_right.t18 a_n2874_n3288# 0.278586f
C192 drain_right.t4 a_n2874_n3288# 0.278586f
C193 drain_right.n18 a_n2874_n3288# 2.479f
C194 drain_right.n19 a_n2874_n3288# 0.382014f
C195 drain_right.t1 a_n2874_n3288# 0.278586f
C196 drain_right.t5 a_n2874_n3288# 0.278586f
C197 drain_right.n20 a_n2874_n3288# 2.479f
C198 drain_right.n21 a_n2874_n3288# 0.634413f
C199 source.n0 a_n2874_n3288# 0.035161f
C200 source.n1 a_n2874_n3288# 0.026544f
C201 source.n2 a_n2874_n3288# 0.014264f
C202 source.n3 a_n2874_n3288# 0.033714f
C203 source.n4 a_n2874_n3288# 0.015103f
C204 source.n5 a_n2874_n3288# 0.026544f
C205 source.n6 a_n2874_n3288# 0.014264f
C206 source.n7 a_n2874_n3288# 0.033714f
C207 source.n8 a_n2874_n3288# 0.015103f
C208 source.n9 a_n2874_n3288# 0.026544f
C209 source.n10 a_n2874_n3288# 0.014683f
C210 source.n11 a_n2874_n3288# 0.033714f
C211 source.n12 a_n2874_n3288# 0.014264f
C212 source.n13 a_n2874_n3288# 0.015103f
C213 source.n14 a_n2874_n3288# 0.026544f
C214 source.n15 a_n2874_n3288# 0.014264f
C215 source.n16 a_n2874_n3288# 0.033714f
C216 source.n17 a_n2874_n3288# 0.015103f
C217 source.n18 a_n2874_n3288# 0.026544f
C218 source.n19 a_n2874_n3288# 0.014264f
C219 source.n20 a_n2874_n3288# 0.025286f
C220 source.n21 a_n2874_n3288# 0.023833f
C221 source.t2 a_n2874_n3288# 0.056941f
C222 source.n22 a_n2874_n3288# 0.19138f
C223 source.n23 a_n2874_n3288# 1.3391f
C224 source.n24 a_n2874_n3288# 0.014264f
C225 source.n25 a_n2874_n3288# 0.015103f
C226 source.n26 a_n2874_n3288# 0.033714f
C227 source.n27 a_n2874_n3288# 0.033714f
C228 source.n28 a_n2874_n3288# 0.015103f
C229 source.n29 a_n2874_n3288# 0.014264f
C230 source.n30 a_n2874_n3288# 0.026544f
C231 source.n31 a_n2874_n3288# 0.026544f
C232 source.n32 a_n2874_n3288# 0.014264f
C233 source.n33 a_n2874_n3288# 0.015103f
C234 source.n34 a_n2874_n3288# 0.033714f
C235 source.n35 a_n2874_n3288# 0.033714f
C236 source.n36 a_n2874_n3288# 0.015103f
C237 source.n37 a_n2874_n3288# 0.014264f
C238 source.n38 a_n2874_n3288# 0.026544f
C239 source.n39 a_n2874_n3288# 0.026544f
C240 source.n40 a_n2874_n3288# 0.014264f
C241 source.n41 a_n2874_n3288# 0.015103f
C242 source.n42 a_n2874_n3288# 0.033714f
C243 source.n43 a_n2874_n3288# 0.033714f
C244 source.n44 a_n2874_n3288# 0.033714f
C245 source.n45 a_n2874_n3288# 0.014683f
C246 source.n46 a_n2874_n3288# 0.014264f
C247 source.n47 a_n2874_n3288# 0.026544f
C248 source.n48 a_n2874_n3288# 0.026544f
C249 source.n49 a_n2874_n3288# 0.014264f
C250 source.n50 a_n2874_n3288# 0.015103f
C251 source.n51 a_n2874_n3288# 0.033714f
C252 source.n52 a_n2874_n3288# 0.033714f
C253 source.n53 a_n2874_n3288# 0.015103f
C254 source.n54 a_n2874_n3288# 0.014264f
C255 source.n55 a_n2874_n3288# 0.026544f
C256 source.n56 a_n2874_n3288# 0.026544f
C257 source.n57 a_n2874_n3288# 0.014264f
C258 source.n58 a_n2874_n3288# 0.015103f
C259 source.n59 a_n2874_n3288# 0.033714f
C260 source.n60 a_n2874_n3288# 0.069185f
C261 source.n61 a_n2874_n3288# 0.015103f
C262 source.n62 a_n2874_n3288# 0.014264f
C263 source.n63 a_n2874_n3288# 0.057004f
C264 source.n64 a_n2874_n3288# 0.038182f
C265 source.n65 a_n2874_n3288# 1.09245f
C266 source.t18 a_n2874_n3288# 0.251711f
C267 source.t6 a_n2874_n3288# 0.251711f
C268 source.n66 a_n2874_n3288# 2.15515f
C269 source.n67 a_n2874_n3288# 0.393777f
C270 source.t21 a_n2874_n3288# 0.251711f
C271 source.t19 a_n2874_n3288# 0.251711f
C272 source.n68 a_n2874_n3288# 2.15515f
C273 source.n69 a_n2874_n3288# 0.393777f
C274 source.t16 a_n2874_n3288# 0.251711f
C275 source.t20 a_n2874_n3288# 0.251711f
C276 source.n70 a_n2874_n3288# 2.15515f
C277 source.n71 a_n2874_n3288# 0.393777f
C278 source.t0 a_n2874_n3288# 0.251711f
C279 source.t17 a_n2874_n3288# 0.251711f
C280 source.n72 a_n2874_n3288# 2.15515f
C281 source.n73 a_n2874_n3288# 0.393777f
C282 source.t8 a_n2874_n3288# 0.251711f
C283 source.t15 a_n2874_n3288# 0.251711f
C284 source.n74 a_n2874_n3288# 2.15515f
C285 source.n75 a_n2874_n3288# 0.393777f
C286 source.n76 a_n2874_n3288# 0.035161f
C287 source.n77 a_n2874_n3288# 0.026544f
C288 source.n78 a_n2874_n3288# 0.014264f
C289 source.n79 a_n2874_n3288# 0.033714f
C290 source.n80 a_n2874_n3288# 0.015103f
C291 source.n81 a_n2874_n3288# 0.026544f
C292 source.n82 a_n2874_n3288# 0.014264f
C293 source.n83 a_n2874_n3288# 0.033714f
C294 source.n84 a_n2874_n3288# 0.015103f
C295 source.n85 a_n2874_n3288# 0.026544f
C296 source.n86 a_n2874_n3288# 0.014683f
C297 source.n87 a_n2874_n3288# 0.033714f
C298 source.n88 a_n2874_n3288# 0.014264f
C299 source.n89 a_n2874_n3288# 0.015103f
C300 source.n90 a_n2874_n3288# 0.026544f
C301 source.n91 a_n2874_n3288# 0.014264f
C302 source.n92 a_n2874_n3288# 0.033714f
C303 source.n93 a_n2874_n3288# 0.015103f
C304 source.n94 a_n2874_n3288# 0.026544f
C305 source.n95 a_n2874_n3288# 0.014264f
C306 source.n96 a_n2874_n3288# 0.025286f
C307 source.n97 a_n2874_n3288# 0.023833f
C308 source.t12 a_n2874_n3288# 0.056941f
C309 source.n98 a_n2874_n3288# 0.19138f
C310 source.n99 a_n2874_n3288# 1.3391f
C311 source.n100 a_n2874_n3288# 0.014264f
C312 source.n101 a_n2874_n3288# 0.015103f
C313 source.n102 a_n2874_n3288# 0.033714f
C314 source.n103 a_n2874_n3288# 0.033714f
C315 source.n104 a_n2874_n3288# 0.015103f
C316 source.n105 a_n2874_n3288# 0.014264f
C317 source.n106 a_n2874_n3288# 0.026544f
C318 source.n107 a_n2874_n3288# 0.026544f
C319 source.n108 a_n2874_n3288# 0.014264f
C320 source.n109 a_n2874_n3288# 0.015103f
C321 source.n110 a_n2874_n3288# 0.033714f
C322 source.n111 a_n2874_n3288# 0.033714f
C323 source.n112 a_n2874_n3288# 0.015103f
C324 source.n113 a_n2874_n3288# 0.014264f
C325 source.n114 a_n2874_n3288# 0.026544f
C326 source.n115 a_n2874_n3288# 0.026544f
C327 source.n116 a_n2874_n3288# 0.014264f
C328 source.n117 a_n2874_n3288# 0.015103f
C329 source.n118 a_n2874_n3288# 0.033714f
C330 source.n119 a_n2874_n3288# 0.033714f
C331 source.n120 a_n2874_n3288# 0.033714f
C332 source.n121 a_n2874_n3288# 0.014683f
C333 source.n122 a_n2874_n3288# 0.014264f
C334 source.n123 a_n2874_n3288# 0.026544f
C335 source.n124 a_n2874_n3288# 0.026544f
C336 source.n125 a_n2874_n3288# 0.014264f
C337 source.n126 a_n2874_n3288# 0.015103f
C338 source.n127 a_n2874_n3288# 0.033714f
C339 source.n128 a_n2874_n3288# 0.033714f
C340 source.n129 a_n2874_n3288# 0.015103f
C341 source.n130 a_n2874_n3288# 0.014264f
C342 source.n131 a_n2874_n3288# 0.026544f
C343 source.n132 a_n2874_n3288# 0.026544f
C344 source.n133 a_n2874_n3288# 0.014264f
C345 source.n134 a_n2874_n3288# 0.015103f
C346 source.n135 a_n2874_n3288# 0.033714f
C347 source.n136 a_n2874_n3288# 0.069185f
C348 source.n137 a_n2874_n3288# 0.015103f
C349 source.n138 a_n2874_n3288# 0.014264f
C350 source.n139 a_n2874_n3288# 0.057004f
C351 source.n140 a_n2874_n3288# 0.038182f
C352 source.n141 a_n2874_n3288# 0.121603f
C353 source.n142 a_n2874_n3288# 0.035161f
C354 source.n143 a_n2874_n3288# 0.026544f
C355 source.n144 a_n2874_n3288# 0.014264f
C356 source.n145 a_n2874_n3288# 0.033714f
C357 source.n146 a_n2874_n3288# 0.015103f
C358 source.n147 a_n2874_n3288# 0.026544f
C359 source.n148 a_n2874_n3288# 0.014264f
C360 source.n149 a_n2874_n3288# 0.033714f
C361 source.n150 a_n2874_n3288# 0.015103f
C362 source.n151 a_n2874_n3288# 0.026544f
C363 source.n152 a_n2874_n3288# 0.014683f
C364 source.n153 a_n2874_n3288# 0.033714f
C365 source.n154 a_n2874_n3288# 0.014264f
C366 source.n155 a_n2874_n3288# 0.015103f
C367 source.n156 a_n2874_n3288# 0.026544f
C368 source.n157 a_n2874_n3288# 0.014264f
C369 source.n158 a_n2874_n3288# 0.033714f
C370 source.n159 a_n2874_n3288# 0.015103f
C371 source.n160 a_n2874_n3288# 0.026544f
C372 source.n161 a_n2874_n3288# 0.014264f
C373 source.n162 a_n2874_n3288# 0.025286f
C374 source.n163 a_n2874_n3288# 0.023833f
C375 source.t28 a_n2874_n3288# 0.056941f
C376 source.n164 a_n2874_n3288# 0.19138f
C377 source.n165 a_n2874_n3288# 1.3391f
C378 source.n166 a_n2874_n3288# 0.014264f
C379 source.n167 a_n2874_n3288# 0.015103f
C380 source.n168 a_n2874_n3288# 0.033714f
C381 source.n169 a_n2874_n3288# 0.033714f
C382 source.n170 a_n2874_n3288# 0.015103f
C383 source.n171 a_n2874_n3288# 0.014264f
C384 source.n172 a_n2874_n3288# 0.026544f
C385 source.n173 a_n2874_n3288# 0.026544f
C386 source.n174 a_n2874_n3288# 0.014264f
C387 source.n175 a_n2874_n3288# 0.015103f
C388 source.n176 a_n2874_n3288# 0.033714f
C389 source.n177 a_n2874_n3288# 0.033714f
C390 source.n178 a_n2874_n3288# 0.015103f
C391 source.n179 a_n2874_n3288# 0.014264f
C392 source.n180 a_n2874_n3288# 0.026544f
C393 source.n181 a_n2874_n3288# 0.026544f
C394 source.n182 a_n2874_n3288# 0.014264f
C395 source.n183 a_n2874_n3288# 0.015103f
C396 source.n184 a_n2874_n3288# 0.033714f
C397 source.n185 a_n2874_n3288# 0.033714f
C398 source.n186 a_n2874_n3288# 0.033714f
C399 source.n187 a_n2874_n3288# 0.014683f
C400 source.n188 a_n2874_n3288# 0.014264f
C401 source.n189 a_n2874_n3288# 0.026544f
C402 source.n190 a_n2874_n3288# 0.026544f
C403 source.n191 a_n2874_n3288# 0.014264f
C404 source.n192 a_n2874_n3288# 0.015103f
C405 source.n193 a_n2874_n3288# 0.033714f
C406 source.n194 a_n2874_n3288# 0.033714f
C407 source.n195 a_n2874_n3288# 0.015103f
C408 source.n196 a_n2874_n3288# 0.014264f
C409 source.n197 a_n2874_n3288# 0.026544f
C410 source.n198 a_n2874_n3288# 0.026544f
C411 source.n199 a_n2874_n3288# 0.014264f
C412 source.n200 a_n2874_n3288# 0.015103f
C413 source.n201 a_n2874_n3288# 0.033714f
C414 source.n202 a_n2874_n3288# 0.069185f
C415 source.n203 a_n2874_n3288# 0.015103f
C416 source.n204 a_n2874_n3288# 0.014264f
C417 source.n205 a_n2874_n3288# 0.057004f
C418 source.n206 a_n2874_n3288# 0.038182f
C419 source.n207 a_n2874_n3288# 0.121603f
C420 source.t37 a_n2874_n3288# 0.251711f
C421 source.t43 a_n2874_n3288# 0.251711f
C422 source.n208 a_n2874_n3288# 2.15515f
C423 source.n209 a_n2874_n3288# 0.393777f
C424 source.t29 a_n2874_n3288# 0.251711f
C425 source.t32 a_n2874_n3288# 0.251711f
C426 source.n210 a_n2874_n3288# 2.15515f
C427 source.n211 a_n2874_n3288# 0.393777f
C428 source.t22 a_n2874_n3288# 0.251711f
C429 source.t40 a_n2874_n3288# 0.251711f
C430 source.n212 a_n2874_n3288# 2.15515f
C431 source.n213 a_n2874_n3288# 0.393777f
C432 source.t24 a_n2874_n3288# 0.251711f
C433 source.t23 a_n2874_n3288# 0.251711f
C434 source.n214 a_n2874_n3288# 2.15515f
C435 source.n215 a_n2874_n3288# 0.393777f
C436 source.t26 a_n2874_n3288# 0.251711f
C437 source.t42 a_n2874_n3288# 0.251711f
C438 source.n216 a_n2874_n3288# 2.15515f
C439 source.n217 a_n2874_n3288# 0.393777f
C440 source.n218 a_n2874_n3288# 0.035161f
C441 source.n219 a_n2874_n3288# 0.026544f
C442 source.n220 a_n2874_n3288# 0.014264f
C443 source.n221 a_n2874_n3288# 0.033714f
C444 source.n222 a_n2874_n3288# 0.015103f
C445 source.n223 a_n2874_n3288# 0.026544f
C446 source.n224 a_n2874_n3288# 0.014264f
C447 source.n225 a_n2874_n3288# 0.033714f
C448 source.n226 a_n2874_n3288# 0.015103f
C449 source.n227 a_n2874_n3288# 0.026544f
C450 source.n228 a_n2874_n3288# 0.014683f
C451 source.n229 a_n2874_n3288# 0.033714f
C452 source.n230 a_n2874_n3288# 0.014264f
C453 source.n231 a_n2874_n3288# 0.015103f
C454 source.n232 a_n2874_n3288# 0.026544f
C455 source.n233 a_n2874_n3288# 0.014264f
C456 source.n234 a_n2874_n3288# 0.033714f
C457 source.n235 a_n2874_n3288# 0.015103f
C458 source.n236 a_n2874_n3288# 0.026544f
C459 source.n237 a_n2874_n3288# 0.014264f
C460 source.n238 a_n2874_n3288# 0.025286f
C461 source.n239 a_n2874_n3288# 0.023833f
C462 source.t31 a_n2874_n3288# 0.056941f
C463 source.n240 a_n2874_n3288# 0.19138f
C464 source.n241 a_n2874_n3288# 1.3391f
C465 source.n242 a_n2874_n3288# 0.014264f
C466 source.n243 a_n2874_n3288# 0.015103f
C467 source.n244 a_n2874_n3288# 0.033714f
C468 source.n245 a_n2874_n3288# 0.033714f
C469 source.n246 a_n2874_n3288# 0.015103f
C470 source.n247 a_n2874_n3288# 0.014264f
C471 source.n248 a_n2874_n3288# 0.026544f
C472 source.n249 a_n2874_n3288# 0.026544f
C473 source.n250 a_n2874_n3288# 0.014264f
C474 source.n251 a_n2874_n3288# 0.015103f
C475 source.n252 a_n2874_n3288# 0.033714f
C476 source.n253 a_n2874_n3288# 0.033714f
C477 source.n254 a_n2874_n3288# 0.015103f
C478 source.n255 a_n2874_n3288# 0.014264f
C479 source.n256 a_n2874_n3288# 0.026544f
C480 source.n257 a_n2874_n3288# 0.026544f
C481 source.n258 a_n2874_n3288# 0.014264f
C482 source.n259 a_n2874_n3288# 0.015103f
C483 source.n260 a_n2874_n3288# 0.033714f
C484 source.n261 a_n2874_n3288# 0.033714f
C485 source.n262 a_n2874_n3288# 0.033714f
C486 source.n263 a_n2874_n3288# 0.014683f
C487 source.n264 a_n2874_n3288# 0.014264f
C488 source.n265 a_n2874_n3288# 0.026544f
C489 source.n266 a_n2874_n3288# 0.026544f
C490 source.n267 a_n2874_n3288# 0.014264f
C491 source.n268 a_n2874_n3288# 0.015103f
C492 source.n269 a_n2874_n3288# 0.033714f
C493 source.n270 a_n2874_n3288# 0.033714f
C494 source.n271 a_n2874_n3288# 0.015103f
C495 source.n272 a_n2874_n3288# 0.014264f
C496 source.n273 a_n2874_n3288# 0.026544f
C497 source.n274 a_n2874_n3288# 0.026544f
C498 source.n275 a_n2874_n3288# 0.014264f
C499 source.n276 a_n2874_n3288# 0.015103f
C500 source.n277 a_n2874_n3288# 0.033714f
C501 source.n278 a_n2874_n3288# 0.069185f
C502 source.n279 a_n2874_n3288# 0.015103f
C503 source.n280 a_n2874_n3288# 0.014264f
C504 source.n281 a_n2874_n3288# 0.057004f
C505 source.n282 a_n2874_n3288# 0.038182f
C506 source.n283 a_n2874_n3288# 1.51514f
C507 source.n284 a_n2874_n3288# 0.035161f
C508 source.n285 a_n2874_n3288# 0.026544f
C509 source.n286 a_n2874_n3288# 0.014264f
C510 source.n287 a_n2874_n3288# 0.033714f
C511 source.n288 a_n2874_n3288# 0.015103f
C512 source.n289 a_n2874_n3288# 0.026544f
C513 source.n290 a_n2874_n3288# 0.014264f
C514 source.n291 a_n2874_n3288# 0.033714f
C515 source.n292 a_n2874_n3288# 0.015103f
C516 source.n293 a_n2874_n3288# 0.026544f
C517 source.n294 a_n2874_n3288# 0.014683f
C518 source.n295 a_n2874_n3288# 0.033714f
C519 source.n296 a_n2874_n3288# 0.015103f
C520 source.n297 a_n2874_n3288# 0.026544f
C521 source.n298 a_n2874_n3288# 0.014264f
C522 source.n299 a_n2874_n3288# 0.033714f
C523 source.n300 a_n2874_n3288# 0.015103f
C524 source.n301 a_n2874_n3288# 0.026544f
C525 source.n302 a_n2874_n3288# 0.014264f
C526 source.n303 a_n2874_n3288# 0.025286f
C527 source.n304 a_n2874_n3288# 0.023833f
C528 source.t14 a_n2874_n3288# 0.056941f
C529 source.n305 a_n2874_n3288# 0.19138f
C530 source.n306 a_n2874_n3288# 1.3391f
C531 source.n307 a_n2874_n3288# 0.014264f
C532 source.n308 a_n2874_n3288# 0.015103f
C533 source.n309 a_n2874_n3288# 0.033714f
C534 source.n310 a_n2874_n3288# 0.033714f
C535 source.n311 a_n2874_n3288# 0.015103f
C536 source.n312 a_n2874_n3288# 0.014264f
C537 source.n313 a_n2874_n3288# 0.026544f
C538 source.n314 a_n2874_n3288# 0.026544f
C539 source.n315 a_n2874_n3288# 0.014264f
C540 source.n316 a_n2874_n3288# 0.015103f
C541 source.n317 a_n2874_n3288# 0.033714f
C542 source.n318 a_n2874_n3288# 0.033714f
C543 source.n319 a_n2874_n3288# 0.015103f
C544 source.n320 a_n2874_n3288# 0.014264f
C545 source.n321 a_n2874_n3288# 0.026544f
C546 source.n322 a_n2874_n3288# 0.026544f
C547 source.n323 a_n2874_n3288# 0.014264f
C548 source.n324 a_n2874_n3288# 0.014264f
C549 source.n325 a_n2874_n3288# 0.015103f
C550 source.n326 a_n2874_n3288# 0.033714f
C551 source.n327 a_n2874_n3288# 0.033714f
C552 source.n328 a_n2874_n3288# 0.033714f
C553 source.n329 a_n2874_n3288# 0.014683f
C554 source.n330 a_n2874_n3288# 0.014264f
C555 source.n331 a_n2874_n3288# 0.026544f
C556 source.n332 a_n2874_n3288# 0.026544f
C557 source.n333 a_n2874_n3288# 0.014264f
C558 source.n334 a_n2874_n3288# 0.015103f
C559 source.n335 a_n2874_n3288# 0.033714f
C560 source.n336 a_n2874_n3288# 0.033714f
C561 source.n337 a_n2874_n3288# 0.015103f
C562 source.n338 a_n2874_n3288# 0.014264f
C563 source.n339 a_n2874_n3288# 0.026544f
C564 source.n340 a_n2874_n3288# 0.026544f
C565 source.n341 a_n2874_n3288# 0.014264f
C566 source.n342 a_n2874_n3288# 0.015103f
C567 source.n343 a_n2874_n3288# 0.033714f
C568 source.n344 a_n2874_n3288# 0.069185f
C569 source.n345 a_n2874_n3288# 0.015103f
C570 source.n346 a_n2874_n3288# 0.014264f
C571 source.n347 a_n2874_n3288# 0.057004f
C572 source.n348 a_n2874_n3288# 0.038182f
C573 source.n349 a_n2874_n3288# 1.51514f
C574 source.t13 a_n2874_n3288# 0.251711f
C575 source.t5 a_n2874_n3288# 0.251711f
C576 source.n350 a_n2874_n3288# 2.15514f
C577 source.n351 a_n2874_n3288# 0.39379f
C578 source.t47 a_n2874_n3288# 0.251711f
C579 source.t1 a_n2874_n3288# 0.251711f
C580 source.n352 a_n2874_n3288# 2.15514f
C581 source.n353 a_n2874_n3288# 0.39379f
C582 source.t11 a_n2874_n3288# 0.251711f
C583 source.t4 a_n2874_n3288# 0.251711f
C584 source.n354 a_n2874_n3288# 2.15514f
C585 source.n355 a_n2874_n3288# 0.39379f
C586 source.t10 a_n2874_n3288# 0.251711f
C587 source.t3 a_n2874_n3288# 0.251711f
C588 source.n356 a_n2874_n3288# 2.15514f
C589 source.n357 a_n2874_n3288# 0.39379f
C590 source.t46 a_n2874_n3288# 0.251711f
C591 source.t9 a_n2874_n3288# 0.251711f
C592 source.n358 a_n2874_n3288# 2.15514f
C593 source.n359 a_n2874_n3288# 0.39379f
C594 source.n360 a_n2874_n3288# 0.035161f
C595 source.n361 a_n2874_n3288# 0.026544f
C596 source.n362 a_n2874_n3288# 0.014264f
C597 source.n363 a_n2874_n3288# 0.033714f
C598 source.n364 a_n2874_n3288# 0.015103f
C599 source.n365 a_n2874_n3288# 0.026544f
C600 source.n366 a_n2874_n3288# 0.014264f
C601 source.n367 a_n2874_n3288# 0.033714f
C602 source.n368 a_n2874_n3288# 0.015103f
C603 source.n369 a_n2874_n3288# 0.026544f
C604 source.n370 a_n2874_n3288# 0.014683f
C605 source.n371 a_n2874_n3288# 0.033714f
C606 source.n372 a_n2874_n3288# 0.015103f
C607 source.n373 a_n2874_n3288# 0.026544f
C608 source.n374 a_n2874_n3288# 0.014264f
C609 source.n375 a_n2874_n3288# 0.033714f
C610 source.n376 a_n2874_n3288# 0.015103f
C611 source.n377 a_n2874_n3288# 0.026544f
C612 source.n378 a_n2874_n3288# 0.014264f
C613 source.n379 a_n2874_n3288# 0.025286f
C614 source.n380 a_n2874_n3288# 0.023833f
C615 source.t7 a_n2874_n3288# 0.056941f
C616 source.n381 a_n2874_n3288# 0.19138f
C617 source.n382 a_n2874_n3288# 1.3391f
C618 source.n383 a_n2874_n3288# 0.014264f
C619 source.n384 a_n2874_n3288# 0.015103f
C620 source.n385 a_n2874_n3288# 0.033714f
C621 source.n386 a_n2874_n3288# 0.033714f
C622 source.n387 a_n2874_n3288# 0.015103f
C623 source.n388 a_n2874_n3288# 0.014264f
C624 source.n389 a_n2874_n3288# 0.026544f
C625 source.n390 a_n2874_n3288# 0.026544f
C626 source.n391 a_n2874_n3288# 0.014264f
C627 source.n392 a_n2874_n3288# 0.015103f
C628 source.n393 a_n2874_n3288# 0.033714f
C629 source.n394 a_n2874_n3288# 0.033714f
C630 source.n395 a_n2874_n3288# 0.015103f
C631 source.n396 a_n2874_n3288# 0.014264f
C632 source.n397 a_n2874_n3288# 0.026544f
C633 source.n398 a_n2874_n3288# 0.026544f
C634 source.n399 a_n2874_n3288# 0.014264f
C635 source.n400 a_n2874_n3288# 0.014264f
C636 source.n401 a_n2874_n3288# 0.015103f
C637 source.n402 a_n2874_n3288# 0.033714f
C638 source.n403 a_n2874_n3288# 0.033714f
C639 source.n404 a_n2874_n3288# 0.033714f
C640 source.n405 a_n2874_n3288# 0.014683f
C641 source.n406 a_n2874_n3288# 0.014264f
C642 source.n407 a_n2874_n3288# 0.026544f
C643 source.n408 a_n2874_n3288# 0.026544f
C644 source.n409 a_n2874_n3288# 0.014264f
C645 source.n410 a_n2874_n3288# 0.015103f
C646 source.n411 a_n2874_n3288# 0.033714f
C647 source.n412 a_n2874_n3288# 0.033714f
C648 source.n413 a_n2874_n3288# 0.015103f
C649 source.n414 a_n2874_n3288# 0.014264f
C650 source.n415 a_n2874_n3288# 0.026544f
C651 source.n416 a_n2874_n3288# 0.026544f
C652 source.n417 a_n2874_n3288# 0.014264f
C653 source.n418 a_n2874_n3288# 0.015103f
C654 source.n419 a_n2874_n3288# 0.033714f
C655 source.n420 a_n2874_n3288# 0.069185f
C656 source.n421 a_n2874_n3288# 0.015103f
C657 source.n422 a_n2874_n3288# 0.014264f
C658 source.n423 a_n2874_n3288# 0.057004f
C659 source.n424 a_n2874_n3288# 0.038182f
C660 source.n425 a_n2874_n3288# 0.121603f
C661 source.n426 a_n2874_n3288# 0.035161f
C662 source.n427 a_n2874_n3288# 0.026544f
C663 source.n428 a_n2874_n3288# 0.014264f
C664 source.n429 a_n2874_n3288# 0.033714f
C665 source.n430 a_n2874_n3288# 0.015103f
C666 source.n431 a_n2874_n3288# 0.026544f
C667 source.n432 a_n2874_n3288# 0.014264f
C668 source.n433 a_n2874_n3288# 0.033714f
C669 source.n434 a_n2874_n3288# 0.015103f
C670 source.n435 a_n2874_n3288# 0.026544f
C671 source.n436 a_n2874_n3288# 0.014683f
C672 source.n437 a_n2874_n3288# 0.033714f
C673 source.n438 a_n2874_n3288# 0.015103f
C674 source.n439 a_n2874_n3288# 0.026544f
C675 source.n440 a_n2874_n3288# 0.014264f
C676 source.n441 a_n2874_n3288# 0.033714f
C677 source.n442 a_n2874_n3288# 0.015103f
C678 source.n443 a_n2874_n3288# 0.026544f
C679 source.n444 a_n2874_n3288# 0.014264f
C680 source.n445 a_n2874_n3288# 0.025286f
C681 source.n446 a_n2874_n3288# 0.023833f
C682 source.t33 a_n2874_n3288# 0.056941f
C683 source.n447 a_n2874_n3288# 0.19138f
C684 source.n448 a_n2874_n3288# 1.3391f
C685 source.n449 a_n2874_n3288# 0.014264f
C686 source.n450 a_n2874_n3288# 0.015103f
C687 source.n451 a_n2874_n3288# 0.033714f
C688 source.n452 a_n2874_n3288# 0.033714f
C689 source.n453 a_n2874_n3288# 0.015103f
C690 source.n454 a_n2874_n3288# 0.014264f
C691 source.n455 a_n2874_n3288# 0.026544f
C692 source.n456 a_n2874_n3288# 0.026544f
C693 source.n457 a_n2874_n3288# 0.014264f
C694 source.n458 a_n2874_n3288# 0.015103f
C695 source.n459 a_n2874_n3288# 0.033714f
C696 source.n460 a_n2874_n3288# 0.033714f
C697 source.n461 a_n2874_n3288# 0.015103f
C698 source.n462 a_n2874_n3288# 0.014264f
C699 source.n463 a_n2874_n3288# 0.026544f
C700 source.n464 a_n2874_n3288# 0.026544f
C701 source.n465 a_n2874_n3288# 0.014264f
C702 source.n466 a_n2874_n3288# 0.014264f
C703 source.n467 a_n2874_n3288# 0.015103f
C704 source.n468 a_n2874_n3288# 0.033714f
C705 source.n469 a_n2874_n3288# 0.033714f
C706 source.n470 a_n2874_n3288# 0.033714f
C707 source.n471 a_n2874_n3288# 0.014683f
C708 source.n472 a_n2874_n3288# 0.014264f
C709 source.n473 a_n2874_n3288# 0.026544f
C710 source.n474 a_n2874_n3288# 0.026544f
C711 source.n475 a_n2874_n3288# 0.014264f
C712 source.n476 a_n2874_n3288# 0.015103f
C713 source.n477 a_n2874_n3288# 0.033714f
C714 source.n478 a_n2874_n3288# 0.033714f
C715 source.n479 a_n2874_n3288# 0.015103f
C716 source.n480 a_n2874_n3288# 0.014264f
C717 source.n481 a_n2874_n3288# 0.026544f
C718 source.n482 a_n2874_n3288# 0.026544f
C719 source.n483 a_n2874_n3288# 0.014264f
C720 source.n484 a_n2874_n3288# 0.015103f
C721 source.n485 a_n2874_n3288# 0.033714f
C722 source.n486 a_n2874_n3288# 0.069185f
C723 source.n487 a_n2874_n3288# 0.015103f
C724 source.n488 a_n2874_n3288# 0.014264f
C725 source.n489 a_n2874_n3288# 0.057004f
C726 source.n490 a_n2874_n3288# 0.038182f
C727 source.n491 a_n2874_n3288# 0.121603f
C728 source.t45 a_n2874_n3288# 0.251711f
C729 source.t38 a_n2874_n3288# 0.251711f
C730 source.n492 a_n2874_n3288# 2.15514f
C731 source.n493 a_n2874_n3288# 0.39379f
C732 source.t39 a_n2874_n3288# 0.251711f
C733 source.t30 a_n2874_n3288# 0.251711f
C734 source.n494 a_n2874_n3288# 2.15514f
C735 source.n495 a_n2874_n3288# 0.39379f
C736 source.t35 a_n2874_n3288# 0.251711f
C737 source.t34 a_n2874_n3288# 0.251711f
C738 source.n496 a_n2874_n3288# 2.15514f
C739 source.n497 a_n2874_n3288# 0.39379f
C740 source.t25 a_n2874_n3288# 0.251711f
C741 source.t44 a_n2874_n3288# 0.251711f
C742 source.n498 a_n2874_n3288# 2.15514f
C743 source.n499 a_n2874_n3288# 0.39379f
C744 source.t41 a_n2874_n3288# 0.251711f
C745 source.t27 a_n2874_n3288# 0.251711f
C746 source.n500 a_n2874_n3288# 2.15514f
C747 source.n501 a_n2874_n3288# 0.39379f
C748 source.n502 a_n2874_n3288# 0.035161f
C749 source.n503 a_n2874_n3288# 0.026544f
C750 source.n504 a_n2874_n3288# 0.014264f
C751 source.n505 a_n2874_n3288# 0.033714f
C752 source.n506 a_n2874_n3288# 0.015103f
C753 source.n507 a_n2874_n3288# 0.026544f
C754 source.n508 a_n2874_n3288# 0.014264f
C755 source.n509 a_n2874_n3288# 0.033714f
C756 source.n510 a_n2874_n3288# 0.015103f
C757 source.n511 a_n2874_n3288# 0.026544f
C758 source.n512 a_n2874_n3288# 0.014683f
C759 source.n513 a_n2874_n3288# 0.033714f
C760 source.n514 a_n2874_n3288# 0.015103f
C761 source.n515 a_n2874_n3288# 0.026544f
C762 source.n516 a_n2874_n3288# 0.014264f
C763 source.n517 a_n2874_n3288# 0.033714f
C764 source.n518 a_n2874_n3288# 0.015103f
C765 source.n519 a_n2874_n3288# 0.026544f
C766 source.n520 a_n2874_n3288# 0.014264f
C767 source.n521 a_n2874_n3288# 0.025286f
C768 source.n522 a_n2874_n3288# 0.023833f
C769 source.t36 a_n2874_n3288# 0.056941f
C770 source.n523 a_n2874_n3288# 0.19138f
C771 source.n524 a_n2874_n3288# 1.3391f
C772 source.n525 a_n2874_n3288# 0.014264f
C773 source.n526 a_n2874_n3288# 0.015103f
C774 source.n527 a_n2874_n3288# 0.033714f
C775 source.n528 a_n2874_n3288# 0.033714f
C776 source.n529 a_n2874_n3288# 0.015103f
C777 source.n530 a_n2874_n3288# 0.014264f
C778 source.n531 a_n2874_n3288# 0.026544f
C779 source.n532 a_n2874_n3288# 0.026544f
C780 source.n533 a_n2874_n3288# 0.014264f
C781 source.n534 a_n2874_n3288# 0.015103f
C782 source.n535 a_n2874_n3288# 0.033714f
C783 source.n536 a_n2874_n3288# 0.033714f
C784 source.n537 a_n2874_n3288# 0.015103f
C785 source.n538 a_n2874_n3288# 0.014264f
C786 source.n539 a_n2874_n3288# 0.026544f
C787 source.n540 a_n2874_n3288# 0.026544f
C788 source.n541 a_n2874_n3288# 0.014264f
C789 source.n542 a_n2874_n3288# 0.014264f
C790 source.n543 a_n2874_n3288# 0.015103f
C791 source.n544 a_n2874_n3288# 0.033714f
C792 source.n545 a_n2874_n3288# 0.033714f
C793 source.n546 a_n2874_n3288# 0.033714f
C794 source.n547 a_n2874_n3288# 0.014683f
C795 source.n548 a_n2874_n3288# 0.014264f
C796 source.n549 a_n2874_n3288# 0.026544f
C797 source.n550 a_n2874_n3288# 0.026544f
C798 source.n551 a_n2874_n3288# 0.014264f
C799 source.n552 a_n2874_n3288# 0.015103f
C800 source.n553 a_n2874_n3288# 0.033714f
C801 source.n554 a_n2874_n3288# 0.033714f
C802 source.n555 a_n2874_n3288# 0.015103f
C803 source.n556 a_n2874_n3288# 0.014264f
C804 source.n557 a_n2874_n3288# 0.026544f
C805 source.n558 a_n2874_n3288# 0.026544f
C806 source.n559 a_n2874_n3288# 0.014264f
C807 source.n560 a_n2874_n3288# 0.015103f
C808 source.n561 a_n2874_n3288# 0.033714f
C809 source.n562 a_n2874_n3288# 0.069185f
C810 source.n563 a_n2874_n3288# 0.015103f
C811 source.n564 a_n2874_n3288# 0.014264f
C812 source.n565 a_n2874_n3288# 0.057004f
C813 source.n566 a_n2874_n3288# 0.038182f
C814 source.n567 a_n2874_n3288# 0.283163f
C815 source.n568 a_n2874_n3288# 1.67355f
C816 minus.n0 a_n2874_n3288# 0.043365f
C817 minus.t5 a_n2874_n3288# 0.74193f
C818 minus.n1 a_n2874_n3288# 0.303424f
C819 minus.t18 a_n2874_n3288# 0.74193f
C820 minus.n2 a_n2874_n3288# 0.043365f
C821 minus.t14 a_n2874_n3288# 0.74193f
C822 minus.n3 a_n2874_n3288# 0.299414f
C823 minus.n4 a_n2874_n3288# 0.043365f
C824 minus.t7 a_n2874_n3288# 0.74193f
C825 minus.n5 a_n2874_n3288# 0.299414f
C826 minus.t13 a_n2874_n3288# 0.74193f
C827 minus.n6 a_n2874_n3288# 0.043365f
C828 minus.t8 a_n2874_n3288# 0.74193f
C829 minus.n7 a_n2874_n3288# 0.303424f
C830 minus.t17 a_n2874_n3288# 0.753472f
C831 minus.t4 a_n2874_n3288# 0.74193f
C832 minus.n8 a_n2874_n3288# 0.308555f
C833 minus.n9 a_n2874_n3288# 0.289159f
C834 minus.n10 a_n2874_n3288# 0.176079f
C835 minus.n11 a_n2874_n3288# 0.043365f
C836 minus.n12 a_n2874_n3288# 0.00984f
C837 minus.t21 a_n2874_n3288# 0.74193f
C838 minus.n13 a_n2874_n3288# 0.303825f
C839 minus.n14 a_n2874_n3288# 0.00984f
C840 minus.n15 a_n2874_n3288# 0.043365f
C841 minus.n16 a_n2874_n3288# 0.043365f
C842 minus.n17 a_n2874_n3288# 0.043365f
C843 minus.n18 a_n2874_n3288# 0.303692f
C844 minus.n19 a_n2874_n3288# 0.00984f
C845 minus.t1 a_n2874_n3288# 0.74193f
C846 minus.n20 a_n2874_n3288# 0.303692f
C847 minus.n21 a_n2874_n3288# 0.043365f
C848 minus.n22 a_n2874_n3288# 0.043365f
C849 minus.n23 a_n2874_n3288# 0.043365f
C850 minus.n24 a_n2874_n3288# 0.00984f
C851 minus.t19 a_n2874_n3288# 0.74193f
C852 minus.n25 a_n2874_n3288# 0.303825f
C853 minus.n26 a_n2874_n3288# 0.00984f
C854 minus.n27 a_n2874_n3288# 0.043365f
C855 minus.n28 a_n2874_n3288# 0.043365f
C856 minus.n29 a_n2874_n3288# 0.043365f
C857 minus.n30 a_n2874_n3288# 0.299681f
C858 minus.n31 a_n2874_n3288# 0.00984f
C859 minus.t22 a_n2874_n3288# 0.74193f
C860 minus.n32 a_n2874_n3288# 0.298879f
C861 minus.n33 a_n2874_n3288# 1.78927f
C862 minus.n34 a_n2874_n3288# 0.043365f
C863 minus.t20 a_n2874_n3288# 0.74193f
C864 minus.n35 a_n2874_n3288# 0.303424f
C865 minus.n36 a_n2874_n3288# 0.043365f
C866 minus.t9 a_n2874_n3288# 0.74193f
C867 minus.n37 a_n2874_n3288# 0.299414f
C868 minus.n38 a_n2874_n3288# 0.043365f
C869 minus.t6 a_n2874_n3288# 0.74193f
C870 minus.n39 a_n2874_n3288# 0.299414f
C871 minus.n40 a_n2874_n3288# 0.043365f
C872 minus.t12 a_n2874_n3288# 0.74193f
C873 minus.n41 a_n2874_n3288# 0.303424f
C874 minus.t3 a_n2874_n3288# 0.753472f
C875 minus.t2 a_n2874_n3288# 0.74193f
C876 minus.n42 a_n2874_n3288# 0.308555f
C877 minus.n43 a_n2874_n3288# 0.289159f
C878 minus.n44 a_n2874_n3288# 0.176079f
C879 minus.n45 a_n2874_n3288# 0.043365f
C880 minus.n46 a_n2874_n3288# 0.00984f
C881 minus.t11 a_n2874_n3288# 0.74193f
C882 minus.n47 a_n2874_n3288# 0.303825f
C883 minus.n48 a_n2874_n3288# 0.00984f
C884 minus.n49 a_n2874_n3288# 0.043365f
C885 minus.n50 a_n2874_n3288# 0.043365f
C886 minus.n51 a_n2874_n3288# 0.043365f
C887 minus.t16 a_n2874_n3288# 0.74193f
C888 minus.n52 a_n2874_n3288# 0.303692f
C889 minus.n53 a_n2874_n3288# 0.00984f
C890 minus.t15 a_n2874_n3288# 0.74193f
C891 minus.n54 a_n2874_n3288# 0.303692f
C892 minus.n55 a_n2874_n3288# 0.043365f
C893 minus.n56 a_n2874_n3288# 0.043365f
C894 minus.n57 a_n2874_n3288# 0.043365f
C895 minus.n58 a_n2874_n3288# 0.00984f
C896 minus.t23 a_n2874_n3288# 0.74193f
C897 minus.n59 a_n2874_n3288# 0.303825f
C898 minus.n60 a_n2874_n3288# 0.00984f
C899 minus.n61 a_n2874_n3288# 0.043365f
C900 minus.n62 a_n2874_n3288# 0.043365f
C901 minus.n63 a_n2874_n3288# 0.043365f
C902 minus.t10 a_n2874_n3288# 0.74193f
C903 minus.n64 a_n2874_n3288# 0.299681f
C904 minus.n65 a_n2874_n3288# 0.00984f
C905 minus.t0 a_n2874_n3288# 0.74193f
C906 minus.n66 a_n2874_n3288# 0.298879f
C907 minus.n67 a_n2874_n3288# 0.286264f
C908 minus.n68 a_n2874_n3288# 2.14816f
.ends

