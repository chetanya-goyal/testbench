* NGSPICE file created from diffpair329.ext - technology: sky130A

.subckt diffpair329 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t40 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X1 drain_left.t22 plus.t1 source.t34 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X2 drain_left.t21 plus.t2 source.t32 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X3 source.t29 plus.t3 drain_left.t20 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X4 source.t43 plus.t4 drain_left.t19 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X5 drain_right.t23 minus.t0 source.t0 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X6 source.t25 plus.t5 drain_left.t18 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X7 drain_left.t17 plus.t6 source.t46 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X8 source.t15 minus.t1 drain_right.t22 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X9 a_n2406_n2688# a_n2406_n2688# a_n2406_n2688# a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=34.2 ps=151.6 w=9 l=0.15
X10 source.t19 minus.t2 drain_right.t21 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X11 drain_left.t16 plus.t7 source.t27 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X12 a_n2406_n2688# a_n2406_n2688# a_n2406_n2688# a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X13 drain_right.t20 minus.t3 source.t23 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X14 drain_left.t15 plus.t8 source.t38 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X15 a_n2406_n2688# a_n2406_n2688# a_n2406_n2688# a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X16 drain_right.t19 minus.t4 source.t16 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X17 source.t1 minus.t5 drain_right.t18 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X18 drain_right.t17 minus.t6 source.t5 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X19 source.t41 plus.t9 drain_left.t14 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X20 drain_right.t16 minus.t7 source.t6 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X21 drain_right.t15 minus.t8 source.t11 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X22 source.t8 minus.t9 drain_right.t14 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X23 a_n2406_n2688# a_n2406_n2688# a_n2406_n2688# a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X24 source.t2 minus.t10 drain_right.t13 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X25 drain_right.t12 minus.t11 source.t10 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X26 source.t13 minus.t12 drain_right.t11 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X27 drain_left.t13 plus.t10 source.t35 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X28 source.t33 plus.t11 drain_left.t12 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X29 drain_right.t10 minus.t13 source.t18 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X30 drain_right.t9 minus.t14 source.t20 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X31 source.t12 minus.t15 drain_right.t8 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X32 source.t30 plus.t12 drain_left.t11 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X33 source.t17 minus.t16 drain_right.t7 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X34 source.t21 minus.t17 drain_right.t6 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X35 drain_left.t10 plus.t13 source.t44 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X36 source.t22 minus.t18 drain_right.t5 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X37 drain_right.t4 minus.t19 source.t4 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X38 drain_right.t3 minus.t20 source.t9 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X39 source.t36 plus.t14 drain_left.t9 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X40 drain_left.t8 plus.t15 source.t26 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X41 source.t47 plus.t16 drain_left.t7 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X42 source.t28 plus.t17 drain_left.t6 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X43 drain_right.t2 minus.t21 source.t3 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X44 source.t7 minus.t22 drain_right.t1 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X45 source.t39 plus.t18 drain_left.t5 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X46 drain_left.t4 plus.t19 source.t42 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X47 drain_left.t3 plus.t20 source.t37 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X48 source.t14 minus.t23 drain_right.t0 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X49 source.t31 plus.t21 drain_left.t2 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X50 drain_left.t1 plus.t22 source.t45 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X51 source.t24 plus.t23 drain_left.t0 a_n2406_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
R0 plus.n6 plus.t11 1702.34
R1 plus.n35 plus.t22 1702.34
R2 plus.n45 plus.t7 1702.34
R3 plus.n72 plus.t4 1702.34
R4 plus.n7 plus.t20 1654.87
R5 plus.n8 plus.t17 1654.87
R6 plus.n14 plus.t13 1654.87
R7 plus.n16 plus.t23 1654.87
R8 plus.n17 plus.t19 1654.87
R9 plus.n23 plus.t16 1654.87
R10 plus.n25 plus.t10 1654.87
R11 plus.n26 plus.t18 1654.87
R12 plus.n32 plus.t15 1654.87
R13 plus.n34 plus.t12 1654.87
R14 plus.n47 plus.t9 1654.87
R15 plus.n46 plus.t1 1654.87
R16 plus.n53 plus.t5 1654.87
R17 plus.n55 plus.t8 1654.87
R18 plus.n43 plus.t21 1654.87
R19 plus.n61 plus.t2 1654.87
R20 plus.n63 plus.t3 1654.87
R21 plus.n40 plus.t6 1654.87
R22 plus.n69 plus.t14 1654.87
R23 plus.n71 plus.t0 1654.87
R24 plus.n10 plus.n6 161.489
R25 plus.n49 plus.n45 161.489
R26 plus.n10 plus.n9 161.3
R27 plus.n11 plus.n5 161.3
R28 plus.n13 plus.n12 161.3
R29 plus.n15 plus.n4 161.3
R30 plus.n19 plus.n18 161.3
R31 plus.n20 plus.n3 161.3
R32 plus.n22 plus.n21 161.3
R33 plus.n24 plus.n2 161.3
R34 plus.n28 plus.n27 161.3
R35 plus.n29 plus.n1 161.3
R36 plus.n31 plus.n30 161.3
R37 plus.n33 plus.n0 161.3
R38 plus.n36 plus.n35 161.3
R39 plus.n49 plus.n48 161.3
R40 plus.n50 plus.n44 161.3
R41 plus.n52 plus.n51 161.3
R42 plus.n54 plus.n42 161.3
R43 plus.n57 plus.n56 161.3
R44 plus.n58 plus.n41 161.3
R45 plus.n60 plus.n59 161.3
R46 plus.n62 plus.n39 161.3
R47 plus.n65 plus.n64 161.3
R48 plus.n66 plus.n38 161.3
R49 plus.n68 plus.n67 161.3
R50 plus.n70 plus.n37 161.3
R51 plus.n73 plus.n72 161.3
R52 plus.n13 plus.n5 73.0308
R53 plus.n22 plus.n3 73.0308
R54 plus.n31 plus.n1 73.0308
R55 plus.n68 plus.n38 73.0308
R56 plus.n60 plus.n41 73.0308
R57 plus.n52 plus.n44 73.0308
R58 plus.n9 plus.n8 69.3793
R59 plus.n33 plus.n32 69.3793
R60 plus.n70 plus.n69 69.3793
R61 plus.n48 plus.n46 69.3793
R62 plus.n18 plus.n17 62.0763
R63 plus.n24 plus.n23 62.0763
R64 plus.n62 plus.n61 62.0763
R65 plus.n56 plus.n43 62.0763
R66 plus.n15 plus.n14 54.7732
R67 plus.n27 plus.n26 54.7732
R68 plus.n64 plus.n40 54.7732
R69 plus.n54 plus.n53 54.7732
R70 plus.n7 plus.n6 47.4702
R71 plus.n35 plus.n34 47.4702
R72 plus.n72 plus.n71 47.4702
R73 plus.n47 plus.n45 47.4702
R74 plus.n16 plus.n15 40.1672
R75 plus.n27 plus.n25 40.1672
R76 plus.n64 plus.n63 40.1672
R77 plus.n55 plus.n54 40.1672
R78 plus.n18 plus.n16 32.8641
R79 plus.n25 plus.n24 32.8641
R80 plus.n63 plus.n62 32.8641
R81 plus.n56 plus.n55 32.8641
R82 plus plus.n73 31.0028
R83 plus.n9 plus.n7 25.5611
R84 plus.n34 plus.n33 25.5611
R85 plus.n71 plus.n70 25.5611
R86 plus.n48 plus.n47 25.5611
R87 plus.n14 plus.n13 18.2581
R88 plus.n26 plus.n1 18.2581
R89 plus.n40 plus.n38 18.2581
R90 plus.n53 plus.n52 18.2581
R91 plus plus.n36 11.0308
R92 plus.n17 plus.n3 10.955
R93 plus.n23 plus.n22 10.955
R94 plus.n61 plus.n60 10.955
R95 plus.n43 plus.n41 10.955
R96 plus.n8 plus.n5 3.65202
R97 plus.n32 plus.n31 3.65202
R98 plus.n69 plus.n68 3.65202
R99 plus.n46 plus.n44 3.65202
R100 plus.n11 plus.n10 0.189894
R101 plus.n12 plus.n11 0.189894
R102 plus.n12 plus.n4 0.189894
R103 plus.n19 plus.n4 0.189894
R104 plus.n20 plus.n19 0.189894
R105 plus.n21 plus.n20 0.189894
R106 plus.n21 plus.n2 0.189894
R107 plus.n28 plus.n2 0.189894
R108 plus.n29 plus.n28 0.189894
R109 plus.n30 plus.n29 0.189894
R110 plus.n30 plus.n0 0.189894
R111 plus.n36 plus.n0 0.189894
R112 plus.n73 plus.n37 0.189894
R113 plus.n67 plus.n37 0.189894
R114 plus.n67 plus.n66 0.189894
R115 plus.n66 plus.n65 0.189894
R116 plus.n65 plus.n39 0.189894
R117 plus.n59 plus.n39 0.189894
R118 plus.n59 plus.n58 0.189894
R119 plus.n58 plus.n57 0.189894
R120 plus.n57 plus.n42 0.189894
R121 plus.n51 plus.n42 0.189894
R122 plus.n51 plus.n50 0.189894
R123 plus.n50 plus.n49 0.189894
R124 source.n11 source.t33 52.1921
R125 source.n12 source.t6 52.1921
R126 source.n23 source.t21 52.1921
R127 source.n47 source.t0 52.1919
R128 source.n36 source.t14 52.1919
R129 source.n35 source.t27 52.1919
R130 source.n24 source.t43 52.1919
R131 source.n0 source.t45 52.1919
R132 source.n2 source.n1 48.8588
R133 source.n4 source.n3 48.8588
R134 source.n6 source.n5 48.8588
R135 source.n8 source.n7 48.8588
R136 source.n10 source.n9 48.8588
R137 source.n14 source.n13 48.8588
R138 source.n16 source.n15 48.8588
R139 source.n18 source.n17 48.8588
R140 source.n20 source.n19 48.8588
R141 source.n22 source.n21 48.8588
R142 source.n46 source.n45 48.8586
R143 source.n44 source.n43 48.8586
R144 source.n42 source.n41 48.8586
R145 source.n40 source.n39 48.8586
R146 source.n38 source.n37 48.8586
R147 source.n34 source.n33 48.8586
R148 source.n32 source.n31 48.8586
R149 source.n30 source.n29 48.8586
R150 source.n28 source.n27 48.8586
R151 source.n26 source.n25 48.8586
R152 source.n24 source.n23 19.5753
R153 source.n48 source.n0 14.0322
R154 source.n48 source.n47 5.5436
R155 source.n45 source.t5 3.33383
R156 source.n45 source.t12 3.33383
R157 source.n43 source.t3 3.33383
R158 source.n43 source.t19 3.33383
R159 source.n41 source.t16 3.33383
R160 source.n41 source.t13 3.33383
R161 source.n39 source.t9 3.33383
R162 source.n39 source.t15 3.33383
R163 source.n37 source.t23 3.33383
R164 source.n37 source.t8 3.33383
R165 source.n33 source.t34 3.33383
R166 source.n33 source.t41 3.33383
R167 source.n31 source.t38 3.33383
R168 source.n31 source.t25 3.33383
R169 source.n29 source.t32 3.33383
R170 source.n29 source.t31 3.33383
R171 source.n27 source.t46 3.33383
R172 source.n27 source.t29 3.33383
R173 source.n25 source.t40 3.33383
R174 source.n25 source.t36 3.33383
R175 source.n1 source.t26 3.33383
R176 source.n1 source.t30 3.33383
R177 source.n3 source.t35 3.33383
R178 source.n3 source.t39 3.33383
R179 source.n5 source.t42 3.33383
R180 source.n5 source.t47 3.33383
R181 source.n7 source.t44 3.33383
R182 source.n7 source.t24 3.33383
R183 source.n9 source.t37 3.33383
R184 source.n9 source.t28 3.33383
R185 source.n13 source.t18 3.33383
R186 source.n13 source.t1 3.33383
R187 source.n15 source.t11 3.33383
R188 source.n15 source.t2 3.33383
R189 source.n17 source.t20 3.33383
R190 source.n17 source.t22 3.33383
R191 source.n19 source.t10 3.33383
R192 source.n19 source.t17 3.33383
R193 source.n21 source.t4 3.33383
R194 source.n21 source.t7 3.33383
R195 source.n23 source.n22 0.560845
R196 source.n22 source.n20 0.560845
R197 source.n20 source.n18 0.560845
R198 source.n18 source.n16 0.560845
R199 source.n16 source.n14 0.560845
R200 source.n14 source.n12 0.560845
R201 source.n11 source.n10 0.560845
R202 source.n10 source.n8 0.560845
R203 source.n8 source.n6 0.560845
R204 source.n6 source.n4 0.560845
R205 source.n4 source.n2 0.560845
R206 source.n2 source.n0 0.560845
R207 source.n26 source.n24 0.560845
R208 source.n28 source.n26 0.560845
R209 source.n30 source.n28 0.560845
R210 source.n32 source.n30 0.560845
R211 source.n34 source.n32 0.560845
R212 source.n35 source.n34 0.560845
R213 source.n38 source.n36 0.560845
R214 source.n40 source.n38 0.560845
R215 source.n42 source.n40 0.560845
R216 source.n44 source.n42 0.560845
R217 source.n46 source.n44 0.560845
R218 source.n47 source.n46 0.560845
R219 source.n12 source.n11 0.470328
R220 source.n36 source.n35 0.470328
R221 source source.n48 0.188
R222 drain_left.n13 drain_left.n11 66.0979
R223 drain_left.n7 drain_left.n5 66.0977
R224 drain_left.n2 drain_left.n0 66.0977
R225 drain_left.n19 drain_left.n18 65.5376
R226 drain_left.n17 drain_left.n16 65.5376
R227 drain_left.n15 drain_left.n14 65.5376
R228 drain_left.n13 drain_left.n12 65.5376
R229 drain_left.n21 drain_left.n20 65.5374
R230 drain_left.n7 drain_left.n6 65.5373
R231 drain_left.n9 drain_left.n8 65.5373
R232 drain_left.n4 drain_left.n3 65.5373
R233 drain_left.n2 drain_left.n1 65.5373
R234 drain_left drain_left.n10 30.4176
R235 drain_left drain_left.n21 6.21356
R236 drain_left.n5 drain_left.t14 3.33383
R237 drain_left.n5 drain_left.t16 3.33383
R238 drain_left.n6 drain_left.t18 3.33383
R239 drain_left.n6 drain_left.t22 3.33383
R240 drain_left.n8 drain_left.t2 3.33383
R241 drain_left.n8 drain_left.t15 3.33383
R242 drain_left.n3 drain_left.t20 3.33383
R243 drain_left.n3 drain_left.t21 3.33383
R244 drain_left.n1 drain_left.t9 3.33383
R245 drain_left.n1 drain_left.t17 3.33383
R246 drain_left.n0 drain_left.t19 3.33383
R247 drain_left.n0 drain_left.t23 3.33383
R248 drain_left.n20 drain_left.t11 3.33383
R249 drain_left.n20 drain_left.t1 3.33383
R250 drain_left.n18 drain_left.t5 3.33383
R251 drain_left.n18 drain_left.t8 3.33383
R252 drain_left.n16 drain_left.t7 3.33383
R253 drain_left.n16 drain_left.t13 3.33383
R254 drain_left.n14 drain_left.t0 3.33383
R255 drain_left.n14 drain_left.t4 3.33383
R256 drain_left.n12 drain_left.t6 3.33383
R257 drain_left.n12 drain_left.t10 3.33383
R258 drain_left.n11 drain_left.t12 3.33383
R259 drain_left.n11 drain_left.t3 3.33383
R260 drain_left.n9 drain_left.n7 0.560845
R261 drain_left.n4 drain_left.n2 0.560845
R262 drain_left.n15 drain_left.n13 0.560845
R263 drain_left.n17 drain_left.n15 0.560845
R264 drain_left.n19 drain_left.n17 0.560845
R265 drain_left.n21 drain_left.n19 0.560845
R266 drain_left.n10 drain_left.n9 0.225326
R267 drain_left.n10 drain_left.n4 0.225326
R268 minus.n35 minus.t17 1702.34
R269 minus.n8 minus.t7 1702.34
R270 minus.n72 minus.t0 1702.34
R271 minus.n43 minus.t23 1702.34
R272 minus.n34 minus.t19 1654.87
R273 minus.n32 minus.t22 1654.87
R274 minus.n3 minus.t11 1654.87
R275 minus.n26 minus.t16 1654.87
R276 minus.n24 minus.t14 1654.87
R277 minus.n6 minus.t18 1654.87
R278 minus.n18 minus.t8 1654.87
R279 minus.n16 minus.t10 1654.87
R280 minus.n9 minus.t13 1654.87
R281 minus.n10 minus.t5 1654.87
R282 minus.n71 minus.t15 1654.87
R283 minus.n69 minus.t6 1654.87
R284 minus.n63 minus.t2 1654.87
R285 minus.n62 minus.t21 1654.87
R286 minus.n60 minus.t12 1654.87
R287 minus.n54 minus.t4 1654.87
R288 minus.n53 minus.t1 1654.87
R289 minus.n51 minus.t20 1654.87
R290 minus.n45 minus.t9 1654.87
R291 minus.n44 minus.t3 1654.87
R292 minus.n12 minus.n8 161.489
R293 minus.n47 minus.n43 161.489
R294 minus.n36 minus.n35 161.3
R295 minus.n33 minus.n0 161.3
R296 minus.n31 minus.n30 161.3
R297 minus.n29 minus.n1 161.3
R298 minus.n28 minus.n27 161.3
R299 minus.n25 minus.n2 161.3
R300 minus.n23 minus.n22 161.3
R301 minus.n21 minus.n4 161.3
R302 minus.n20 minus.n19 161.3
R303 minus.n17 minus.n5 161.3
R304 minus.n15 minus.n14 161.3
R305 minus.n13 minus.n7 161.3
R306 minus.n12 minus.n11 161.3
R307 minus.n73 minus.n72 161.3
R308 minus.n70 minus.n37 161.3
R309 minus.n68 minus.n67 161.3
R310 minus.n66 minus.n38 161.3
R311 minus.n65 minus.n64 161.3
R312 minus.n61 minus.n39 161.3
R313 minus.n59 minus.n58 161.3
R314 minus.n57 minus.n40 161.3
R315 minus.n56 minus.n55 161.3
R316 minus.n52 minus.n41 161.3
R317 minus.n50 minus.n49 161.3
R318 minus.n48 minus.n42 161.3
R319 minus.n47 minus.n46 161.3
R320 minus.n31 minus.n1 73.0308
R321 minus.n23 minus.n4 73.0308
R322 minus.n15 minus.n7 73.0308
R323 minus.n50 minus.n42 73.0308
R324 minus.n59 minus.n40 73.0308
R325 minus.n68 minus.n38 73.0308
R326 minus.n33 minus.n32 69.3793
R327 minus.n11 minus.n9 69.3793
R328 minus.n46 minus.n45 69.3793
R329 minus.n70 minus.n69 69.3793
R330 minus.n25 minus.n24 62.0763
R331 minus.n19 minus.n6 62.0763
R332 minus.n55 minus.n54 62.0763
R333 minus.n61 minus.n60 62.0763
R334 minus.n27 minus.n3 54.7732
R335 minus.n17 minus.n16 54.7732
R336 minus.n52 minus.n51 54.7732
R337 minus.n64 minus.n63 54.7732
R338 minus.n35 minus.n34 47.4702
R339 minus.n10 minus.n8 47.4702
R340 minus.n44 minus.n43 47.4702
R341 minus.n72 minus.n71 47.4702
R342 minus.n27 minus.n26 40.1672
R343 minus.n18 minus.n17 40.1672
R344 minus.n53 minus.n52 40.1672
R345 minus.n64 minus.n62 40.1672
R346 minus.n74 minus.n36 35.9853
R347 minus.n26 minus.n25 32.8641
R348 minus.n19 minus.n18 32.8641
R349 minus.n55 minus.n53 32.8641
R350 minus.n62 minus.n61 32.8641
R351 minus.n34 minus.n33 25.5611
R352 minus.n11 minus.n10 25.5611
R353 minus.n46 minus.n44 25.5611
R354 minus.n71 minus.n70 25.5611
R355 minus.n3 minus.n1 18.2581
R356 minus.n16 minus.n15 18.2581
R357 minus.n51 minus.n50 18.2581
R358 minus.n63 minus.n38 18.2581
R359 minus.n24 minus.n23 10.955
R360 minus.n6 minus.n4 10.955
R361 minus.n54 minus.n40 10.955
R362 minus.n60 minus.n59 10.955
R363 minus.n74 minus.n73 6.52323
R364 minus.n32 minus.n31 3.65202
R365 minus.n9 minus.n7 3.65202
R366 minus.n45 minus.n42 3.65202
R367 minus.n69 minus.n68 3.65202
R368 minus.n36 minus.n0 0.189894
R369 minus.n30 minus.n0 0.189894
R370 minus.n30 minus.n29 0.189894
R371 minus.n29 minus.n28 0.189894
R372 minus.n28 minus.n2 0.189894
R373 minus.n22 minus.n2 0.189894
R374 minus.n22 minus.n21 0.189894
R375 minus.n21 minus.n20 0.189894
R376 minus.n20 minus.n5 0.189894
R377 minus.n14 minus.n5 0.189894
R378 minus.n14 minus.n13 0.189894
R379 minus.n13 minus.n12 0.189894
R380 minus.n48 minus.n47 0.189894
R381 minus.n49 minus.n48 0.189894
R382 minus.n49 minus.n41 0.189894
R383 minus.n56 minus.n41 0.189894
R384 minus.n57 minus.n56 0.189894
R385 minus.n58 minus.n57 0.189894
R386 minus.n58 minus.n39 0.189894
R387 minus.n65 minus.n39 0.189894
R388 minus.n66 minus.n65 0.189894
R389 minus.n67 minus.n66 0.189894
R390 minus.n67 minus.n37 0.189894
R391 minus.n73 minus.n37 0.189894
R392 minus minus.n74 0.188
R393 drain_right.n13 drain_right.n11 66.0978
R394 drain_right.n7 drain_right.n5 66.0977
R395 drain_right.n2 drain_right.n0 66.0977
R396 drain_right.n13 drain_right.n12 65.5376
R397 drain_right.n15 drain_right.n14 65.5376
R398 drain_right.n17 drain_right.n16 65.5376
R399 drain_right.n19 drain_right.n18 65.5376
R400 drain_right.n21 drain_right.n20 65.5376
R401 drain_right.n7 drain_right.n6 65.5373
R402 drain_right.n9 drain_right.n8 65.5373
R403 drain_right.n4 drain_right.n3 65.5373
R404 drain_right.n2 drain_right.n1 65.5373
R405 drain_right drain_right.n10 29.8644
R406 drain_right drain_right.n21 6.21356
R407 drain_right.n5 drain_right.t8 3.33383
R408 drain_right.n5 drain_right.t23 3.33383
R409 drain_right.n6 drain_right.t21 3.33383
R410 drain_right.n6 drain_right.t17 3.33383
R411 drain_right.n8 drain_right.t11 3.33383
R412 drain_right.n8 drain_right.t2 3.33383
R413 drain_right.n3 drain_right.t22 3.33383
R414 drain_right.n3 drain_right.t19 3.33383
R415 drain_right.n1 drain_right.t14 3.33383
R416 drain_right.n1 drain_right.t3 3.33383
R417 drain_right.n0 drain_right.t0 3.33383
R418 drain_right.n0 drain_right.t20 3.33383
R419 drain_right.n11 drain_right.t18 3.33383
R420 drain_right.n11 drain_right.t16 3.33383
R421 drain_right.n12 drain_right.t13 3.33383
R422 drain_right.n12 drain_right.t10 3.33383
R423 drain_right.n14 drain_right.t5 3.33383
R424 drain_right.n14 drain_right.t15 3.33383
R425 drain_right.n16 drain_right.t7 3.33383
R426 drain_right.n16 drain_right.t9 3.33383
R427 drain_right.n18 drain_right.t1 3.33383
R428 drain_right.n18 drain_right.t12 3.33383
R429 drain_right.n20 drain_right.t6 3.33383
R430 drain_right.n20 drain_right.t4 3.33383
R431 drain_right.n9 drain_right.n7 0.560845
R432 drain_right.n4 drain_right.n2 0.560845
R433 drain_right.n21 drain_right.n19 0.560845
R434 drain_right.n19 drain_right.n17 0.560845
R435 drain_right.n17 drain_right.n15 0.560845
R436 drain_right.n15 drain_right.n13 0.560845
R437 drain_right.n10 drain_right.n9 0.225326
R438 drain_right.n10 drain_right.n4 0.225326
C0 plus source 3.57326f
C1 drain_left source 35.0195f
C2 drain_right source 35.0202f
C3 minus source 3.55922f
C4 drain_left plus 4.08981f
C5 plus drain_right 0.392113f
C6 drain_left drain_right 1.29455f
C7 plus minus 5.58595f
C8 drain_left minus 0.171476f
C9 drain_right minus 3.85203f
C10 drain_right a_n2406_n2688# 6.27758f
C11 drain_left a_n2406_n2688# 6.62512f
C12 source a_n2406_n2688# 7.439424f
C13 minus a_n2406_n2688# 8.711829f
C14 plus a_n2406_n2688# 10.721651f
C15 drain_right.t0 a_n2406_n2688# 0.304526f
C16 drain_right.t20 a_n2406_n2688# 0.304526f
C17 drain_right.n0 a_n2406_n2688# 1.96793f
C18 drain_right.t14 a_n2406_n2688# 0.304526f
C19 drain_right.t3 a_n2406_n2688# 0.304526f
C20 drain_right.n1 a_n2406_n2688# 1.96505f
C21 drain_right.n2 a_n2406_n2688# 0.665334f
C22 drain_right.t22 a_n2406_n2688# 0.304526f
C23 drain_right.t19 a_n2406_n2688# 0.304526f
C24 drain_right.n3 a_n2406_n2688# 1.96505f
C25 drain_right.n4 a_n2406_n2688# 0.300778f
C26 drain_right.t8 a_n2406_n2688# 0.304526f
C27 drain_right.t23 a_n2406_n2688# 0.304526f
C28 drain_right.n5 a_n2406_n2688# 1.96793f
C29 drain_right.t21 a_n2406_n2688# 0.304526f
C30 drain_right.t17 a_n2406_n2688# 0.304526f
C31 drain_right.n6 a_n2406_n2688# 1.96505f
C32 drain_right.n7 a_n2406_n2688# 0.665334f
C33 drain_right.t11 a_n2406_n2688# 0.304526f
C34 drain_right.t2 a_n2406_n2688# 0.304526f
C35 drain_right.n8 a_n2406_n2688# 1.96505f
C36 drain_right.n9 a_n2406_n2688# 0.300778f
C37 drain_right.n10 a_n2406_n2688# 1.30041f
C38 drain_right.t18 a_n2406_n2688# 0.304526f
C39 drain_right.t16 a_n2406_n2688# 0.304526f
C40 drain_right.n11 a_n2406_n2688# 1.96792f
C41 drain_right.t13 a_n2406_n2688# 0.304526f
C42 drain_right.t10 a_n2406_n2688# 0.304526f
C43 drain_right.n12 a_n2406_n2688# 1.96505f
C44 drain_right.n13 a_n2406_n2688# 0.665334f
C45 drain_right.t5 a_n2406_n2688# 0.304526f
C46 drain_right.t15 a_n2406_n2688# 0.304526f
C47 drain_right.n14 a_n2406_n2688# 1.96505f
C48 drain_right.n15 a_n2406_n2688# 0.328413f
C49 drain_right.t7 a_n2406_n2688# 0.304526f
C50 drain_right.t9 a_n2406_n2688# 0.304526f
C51 drain_right.n16 a_n2406_n2688# 1.96505f
C52 drain_right.n17 a_n2406_n2688# 0.328413f
C53 drain_right.t1 a_n2406_n2688# 0.304526f
C54 drain_right.t12 a_n2406_n2688# 0.304526f
C55 drain_right.n18 a_n2406_n2688# 1.96505f
C56 drain_right.n19 a_n2406_n2688# 0.328413f
C57 drain_right.t6 a_n2406_n2688# 0.304526f
C58 drain_right.t4 a_n2406_n2688# 0.304526f
C59 drain_right.n20 a_n2406_n2688# 1.96505f
C60 drain_right.n21 a_n2406_n2688# 0.564414f
C61 minus.n0 a_n2406_n2688# 0.051104f
C62 minus.t17 a_n2406_n2688# 0.197966f
C63 minus.t19 a_n2406_n2688# 0.195492f
C64 minus.t22 a_n2406_n2688# 0.195492f
C65 minus.n1 a_n2406_n2688# 0.020891f
C66 minus.n2 a_n2406_n2688# 0.051104f
C67 minus.t11 a_n2406_n2688# 0.195492f
C68 minus.n3 a_n2406_n2688# 0.089511f
C69 minus.t16 a_n2406_n2688# 0.195492f
C70 minus.t14 a_n2406_n2688# 0.195492f
C71 minus.n4 a_n2406_n2688# 0.019316f
C72 minus.n5 a_n2406_n2688# 0.051104f
C73 minus.t18 a_n2406_n2688# 0.195492f
C74 minus.n6 a_n2406_n2688# 0.089511f
C75 minus.t8 a_n2406_n2688# 0.195492f
C76 minus.t10 a_n2406_n2688# 0.195492f
C77 minus.n7 a_n2406_n2688# 0.017741f
C78 minus.t7 a_n2406_n2688# 0.197966f
C79 minus.n8 a_n2406_n2688# 0.108f
C80 minus.t13 a_n2406_n2688# 0.195492f
C81 minus.n9 a_n2406_n2688# 0.089511f
C82 minus.t5 a_n2406_n2688# 0.195492f
C83 minus.n10 a_n2406_n2688# 0.089511f
C84 minus.n11 a_n2406_n2688# 0.021679f
C85 minus.n12 a_n2406_n2688# 0.11159f
C86 minus.n13 a_n2406_n2688# 0.051104f
C87 minus.n14 a_n2406_n2688# 0.051104f
C88 minus.n15 a_n2406_n2688# 0.020891f
C89 minus.n16 a_n2406_n2688# 0.089511f
C90 minus.n17 a_n2406_n2688# 0.021679f
C91 minus.n18 a_n2406_n2688# 0.089511f
C92 minus.n19 a_n2406_n2688# 0.021679f
C93 minus.n20 a_n2406_n2688# 0.051104f
C94 minus.n21 a_n2406_n2688# 0.051104f
C95 minus.n22 a_n2406_n2688# 0.051104f
C96 minus.n23 a_n2406_n2688# 0.019316f
C97 minus.n24 a_n2406_n2688# 0.089511f
C98 minus.n25 a_n2406_n2688# 0.021679f
C99 minus.n26 a_n2406_n2688# 0.089511f
C100 minus.n27 a_n2406_n2688# 0.021679f
C101 minus.n28 a_n2406_n2688# 0.051104f
C102 minus.n29 a_n2406_n2688# 0.051104f
C103 minus.n30 a_n2406_n2688# 0.051104f
C104 minus.n31 a_n2406_n2688# 0.017741f
C105 minus.n32 a_n2406_n2688# 0.089511f
C106 minus.n33 a_n2406_n2688# 0.021679f
C107 minus.n34 a_n2406_n2688# 0.089511f
C108 minus.n35 a_n2406_n2688# 0.107928f
C109 minus.n36 a_n2406_n2688# 1.79074f
C110 minus.n37 a_n2406_n2688# 0.051104f
C111 minus.t15 a_n2406_n2688# 0.195492f
C112 minus.t6 a_n2406_n2688# 0.195492f
C113 minus.n38 a_n2406_n2688# 0.020891f
C114 minus.n39 a_n2406_n2688# 0.051104f
C115 minus.t21 a_n2406_n2688# 0.195492f
C116 minus.t12 a_n2406_n2688# 0.195492f
C117 minus.n40 a_n2406_n2688# 0.019316f
C118 minus.n41 a_n2406_n2688# 0.051104f
C119 minus.t1 a_n2406_n2688# 0.195492f
C120 minus.t20 a_n2406_n2688# 0.195492f
C121 minus.n42 a_n2406_n2688# 0.017741f
C122 minus.t23 a_n2406_n2688# 0.197966f
C123 minus.n43 a_n2406_n2688# 0.108f
C124 minus.t3 a_n2406_n2688# 0.195492f
C125 minus.n44 a_n2406_n2688# 0.089511f
C126 minus.t9 a_n2406_n2688# 0.195492f
C127 minus.n45 a_n2406_n2688# 0.089511f
C128 minus.n46 a_n2406_n2688# 0.021679f
C129 minus.n47 a_n2406_n2688# 0.11159f
C130 minus.n48 a_n2406_n2688# 0.051104f
C131 minus.n49 a_n2406_n2688# 0.051104f
C132 minus.n50 a_n2406_n2688# 0.020891f
C133 minus.n51 a_n2406_n2688# 0.089511f
C134 minus.n52 a_n2406_n2688# 0.021679f
C135 minus.n53 a_n2406_n2688# 0.089511f
C136 minus.t4 a_n2406_n2688# 0.195492f
C137 minus.n54 a_n2406_n2688# 0.089511f
C138 minus.n55 a_n2406_n2688# 0.021679f
C139 minus.n56 a_n2406_n2688# 0.051104f
C140 minus.n57 a_n2406_n2688# 0.051104f
C141 minus.n58 a_n2406_n2688# 0.051104f
C142 minus.n59 a_n2406_n2688# 0.019316f
C143 minus.n60 a_n2406_n2688# 0.089511f
C144 minus.n61 a_n2406_n2688# 0.021679f
C145 minus.n62 a_n2406_n2688# 0.089511f
C146 minus.t2 a_n2406_n2688# 0.195492f
C147 minus.n63 a_n2406_n2688# 0.089511f
C148 minus.n64 a_n2406_n2688# 0.021679f
C149 minus.n65 a_n2406_n2688# 0.051104f
C150 minus.n66 a_n2406_n2688# 0.051104f
C151 minus.n67 a_n2406_n2688# 0.051104f
C152 minus.n68 a_n2406_n2688# 0.017741f
C153 minus.n69 a_n2406_n2688# 0.089511f
C154 minus.n70 a_n2406_n2688# 0.021679f
C155 minus.n71 a_n2406_n2688# 0.089511f
C156 minus.t0 a_n2406_n2688# 0.197966f
C157 minus.n72 a_n2406_n2688# 0.107928f
C158 minus.n73 a_n2406_n2688# 0.336899f
C159 minus.n74 a_n2406_n2688# 2.1756f
C160 drain_left.t19 a_n2406_n2688# 0.305225f
C161 drain_left.t23 a_n2406_n2688# 0.305225f
C162 drain_left.n0 a_n2406_n2688# 1.97244f
C163 drain_left.t9 a_n2406_n2688# 0.305225f
C164 drain_left.t17 a_n2406_n2688# 0.305225f
C165 drain_left.n1 a_n2406_n2688# 1.96955f
C166 drain_left.n2 a_n2406_n2688# 0.666859f
C167 drain_left.t20 a_n2406_n2688# 0.305225f
C168 drain_left.t21 a_n2406_n2688# 0.305225f
C169 drain_left.n3 a_n2406_n2688# 1.96955f
C170 drain_left.n4 a_n2406_n2688# 0.301467f
C171 drain_left.t14 a_n2406_n2688# 0.305225f
C172 drain_left.t16 a_n2406_n2688# 0.305225f
C173 drain_left.n5 a_n2406_n2688# 1.97244f
C174 drain_left.t18 a_n2406_n2688# 0.305225f
C175 drain_left.t22 a_n2406_n2688# 0.305225f
C176 drain_left.n6 a_n2406_n2688# 1.96955f
C177 drain_left.n7 a_n2406_n2688# 0.666859f
C178 drain_left.t2 a_n2406_n2688# 0.305225f
C179 drain_left.t15 a_n2406_n2688# 0.305225f
C180 drain_left.n8 a_n2406_n2688# 1.96955f
C181 drain_left.n9 a_n2406_n2688# 0.301467f
C182 drain_left.n10 a_n2406_n2688# 1.36113f
C183 drain_left.t12 a_n2406_n2688# 0.305225f
C184 drain_left.t3 a_n2406_n2688# 0.305225f
C185 drain_left.n11 a_n2406_n2688# 1.97244f
C186 drain_left.t6 a_n2406_n2688# 0.305225f
C187 drain_left.t10 a_n2406_n2688# 0.305225f
C188 drain_left.n12 a_n2406_n2688# 1.96956f
C189 drain_left.n13 a_n2406_n2688# 0.666853f
C190 drain_left.t0 a_n2406_n2688# 0.305225f
C191 drain_left.t4 a_n2406_n2688# 0.305225f
C192 drain_left.n14 a_n2406_n2688# 1.96956f
C193 drain_left.n15 a_n2406_n2688# 0.329166f
C194 drain_left.t7 a_n2406_n2688# 0.305225f
C195 drain_left.t13 a_n2406_n2688# 0.305225f
C196 drain_left.n16 a_n2406_n2688# 1.96956f
C197 drain_left.n17 a_n2406_n2688# 0.329166f
C198 drain_left.t5 a_n2406_n2688# 0.305225f
C199 drain_left.t8 a_n2406_n2688# 0.305225f
C200 drain_left.n18 a_n2406_n2688# 1.96956f
C201 drain_left.n19 a_n2406_n2688# 0.329166f
C202 drain_left.t11 a_n2406_n2688# 0.305225f
C203 drain_left.t1 a_n2406_n2688# 0.305225f
C204 drain_left.n20 a_n2406_n2688# 1.96955f
C205 drain_left.n21 a_n2406_n2688# 0.565715f
C206 source.t45 a_n2406_n2688# 2.1023f
C207 source.n0 a_n2406_n2688# 1.1727f
C208 source.t26 a_n2406_n2688# 0.278167f
C209 source.t30 a_n2406_n2688# 0.278167f
C210 source.n1 a_n2406_n2688# 1.72605f
C211 source.n2 a_n2406_n2688# 0.333807f
C212 source.t35 a_n2406_n2688# 0.278167f
C213 source.t39 a_n2406_n2688# 0.278167f
C214 source.n3 a_n2406_n2688# 1.72605f
C215 source.n4 a_n2406_n2688# 0.333807f
C216 source.t42 a_n2406_n2688# 0.278167f
C217 source.t47 a_n2406_n2688# 0.278167f
C218 source.n5 a_n2406_n2688# 1.72605f
C219 source.n6 a_n2406_n2688# 0.333807f
C220 source.t44 a_n2406_n2688# 0.278167f
C221 source.t24 a_n2406_n2688# 0.278167f
C222 source.n7 a_n2406_n2688# 1.72605f
C223 source.n8 a_n2406_n2688# 0.333807f
C224 source.t37 a_n2406_n2688# 0.278167f
C225 source.t28 a_n2406_n2688# 0.278167f
C226 source.n9 a_n2406_n2688# 1.72605f
C227 source.n10 a_n2406_n2688# 0.333807f
C228 source.t33 a_n2406_n2688# 2.1023f
C229 source.n11 a_n2406_n2688# 0.450729f
C230 source.t6 a_n2406_n2688# 2.1023f
C231 source.n12 a_n2406_n2688# 0.450729f
C232 source.t18 a_n2406_n2688# 0.278167f
C233 source.t1 a_n2406_n2688# 0.278167f
C234 source.n13 a_n2406_n2688# 1.72605f
C235 source.n14 a_n2406_n2688# 0.333807f
C236 source.t11 a_n2406_n2688# 0.278167f
C237 source.t2 a_n2406_n2688# 0.278167f
C238 source.n15 a_n2406_n2688# 1.72605f
C239 source.n16 a_n2406_n2688# 0.333807f
C240 source.t20 a_n2406_n2688# 0.278167f
C241 source.t22 a_n2406_n2688# 0.278167f
C242 source.n17 a_n2406_n2688# 1.72605f
C243 source.n18 a_n2406_n2688# 0.333807f
C244 source.t10 a_n2406_n2688# 0.278167f
C245 source.t17 a_n2406_n2688# 0.278167f
C246 source.n19 a_n2406_n2688# 1.72605f
C247 source.n20 a_n2406_n2688# 0.333807f
C248 source.t4 a_n2406_n2688# 0.278167f
C249 source.t7 a_n2406_n2688# 0.278167f
C250 source.n21 a_n2406_n2688# 1.72605f
C251 source.n22 a_n2406_n2688# 0.333807f
C252 source.t21 a_n2406_n2688# 2.1023f
C253 source.n23 a_n2406_n2688# 1.54824f
C254 source.t43 a_n2406_n2688# 2.1023f
C255 source.n24 a_n2406_n2688# 1.54825f
C256 source.t40 a_n2406_n2688# 0.278167f
C257 source.t36 a_n2406_n2688# 0.278167f
C258 source.n25 a_n2406_n2688# 1.72605f
C259 source.n26 a_n2406_n2688# 0.333812f
C260 source.t46 a_n2406_n2688# 0.278167f
C261 source.t29 a_n2406_n2688# 0.278167f
C262 source.n27 a_n2406_n2688# 1.72605f
C263 source.n28 a_n2406_n2688# 0.333812f
C264 source.t32 a_n2406_n2688# 0.278167f
C265 source.t31 a_n2406_n2688# 0.278167f
C266 source.n29 a_n2406_n2688# 1.72605f
C267 source.n30 a_n2406_n2688# 0.333812f
C268 source.t38 a_n2406_n2688# 0.278167f
C269 source.t25 a_n2406_n2688# 0.278167f
C270 source.n31 a_n2406_n2688# 1.72605f
C271 source.n32 a_n2406_n2688# 0.333812f
C272 source.t34 a_n2406_n2688# 0.278167f
C273 source.t41 a_n2406_n2688# 0.278167f
C274 source.n33 a_n2406_n2688# 1.72605f
C275 source.n34 a_n2406_n2688# 0.333812f
C276 source.t27 a_n2406_n2688# 2.1023f
C277 source.n35 a_n2406_n2688# 0.450734f
C278 source.t14 a_n2406_n2688# 2.1023f
C279 source.n36 a_n2406_n2688# 0.450734f
C280 source.t23 a_n2406_n2688# 0.278167f
C281 source.t8 a_n2406_n2688# 0.278167f
C282 source.n37 a_n2406_n2688# 1.72605f
C283 source.n38 a_n2406_n2688# 0.333812f
C284 source.t9 a_n2406_n2688# 0.278167f
C285 source.t15 a_n2406_n2688# 0.278167f
C286 source.n39 a_n2406_n2688# 1.72605f
C287 source.n40 a_n2406_n2688# 0.333812f
C288 source.t16 a_n2406_n2688# 0.278167f
C289 source.t13 a_n2406_n2688# 0.278167f
C290 source.n41 a_n2406_n2688# 1.72605f
C291 source.n42 a_n2406_n2688# 0.333812f
C292 source.t3 a_n2406_n2688# 0.278167f
C293 source.t19 a_n2406_n2688# 0.278167f
C294 source.n43 a_n2406_n2688# 1.72605f
C295 source.n44 a_n2406_n2688# 0.333812f
C296 source.t5 a_n2406_n2688# 0.278167f
C297 source.t12 a_n2406_n2688# 0.278167f
C298 source.n45 a_n2406_n2688# 1.72605f
C299 source.n46 a_n2406_n2688# 0.333812f
C300 source.t0 a_n2406_n2688# 2.1023f
C301 source.n47 a_n2406_n2688# 0.597598f
C302 source.n48 a_n2406_n2688# 1.34455f
C303 plus.n0 a_n2406_n2688# 0.052297f
C304 plus.t12 a_n2406_n2688# 0.200055f
C305 plus.t15 a_n2406_n2688# 0.200055f
C306 plus.n1 a_n2406_n2688# 0.021379f
C307 plus.n2 a_n2406_n2688# 0.052297f
C308 plus.t10 a_n2406_n2688# 0.200055f
C309 plus.t16 a_n2406_n2688# 0.200055f
C310 plus.n3 a_n2406_n2688# 0.019767f
C311 plus.n4 a_n2406_n2688# 0.052297f
C312 plus.t23 a_n2406_n2688# 0.200055f
C313 plus.t13 a_n2406_n2688# 0.200055f
C314 plus.n5 a_n2406_n2688# 0.018155f
C315 plus.t11 a_n2406_n2688# 0.202587f
C316 plus.n6 a_n2406_n2688# 0.11052f
C317 plus.t20 a_n2406_n2688# 0.200055f
C318 plus.n7 a_n2406_n2688# 0.0916f
C319 plus.t17 a_n2406_n2688# 0.200055f
C320 plus.n8 a_n2406_n2688# 0.0916f
C321 plus.n9 a_n2406_n2688# 0.022185f
C322 plus.n10 a_n2406_n2688# 0.114194f
C323 plus.n11 a_n2406_n2688# 0.052297f
C324 plus.n12 a_n2406_n2688# 0.052297f
C325 plus.n13 a_n2406_n2688# 0.021379f
C326 plus.n14 a_n2406_n2688# 0.0916f
C327 plus.n15 a_n2406_n2688# 0.022185f
C328 plus.n16 a_n2406_n2688# 0.0916f
C329 plus.t19 a_n2406_n2688# 0.200055f
C330 plus.n17 a_n2406_n2688# 0.0916f
C331 plus.n18 a_n2406_n2688# 0.022185f
C332 plus.n19 a_n2406_n2688# 0.052297f
C333 plus.n20 a_n2406_n2688# 0.052297f
C334 plus.n21 a_n2406_n2688# 0.052297f
C335 plus.n22 a_n2406_n2688# 0.019767f
C336 plus.n23 a_n2406_n2688# 0.0916f
C337 plus.n24 a_n2406_n2688# 0.022185f
C338 plus.n25 a_n2406_n2688# 0.0916f
C339 plus.t18 a_n2406_n2688# 0.200055f
C340 plus.n26 a_n2406_n2688# 0.0916f
C341 plus.n27 a_n2406_n2688# 0.022185f
C342 plus.n28 a_n2406_n2688# 0.052297f
C343 plus.n29 a_n2406_n2688# 0.052297f
C344 plus.n30 a_n2406_n2688# 0.052297f
C345 plus.n31 a_n2406_n2688# 0.018155f
C346 plus.n32 a_n2406_n2688# 0.0916f
C347 plus.n33 a_n2406_n2688# 0.022185f
C348 plus.n34 a_n2406_n2688# 0.0916f
C349 plus.t22 a_n2406_n2688# 0.202587f
C350 plus.n35 a_n2406_n2688# 0.110448f
C351 plus.n36 a_n2406_n2688# 0.516656f
C352 plus.n37 a_n2406_n2688# 0.052297f
C353 plus.t4 a_n2406_n2688# 0.202587f
C354 plus.t0 a_n2406_n2688# 0.200055f
C355 plus.t14 a_n2406_n2688# 0.200055f
C356 plus.n38 a_n2406_n2688# 0.021379f
C357 plus.n39 a_n2406_n2688# 0.052297f
C358 plus.t6 a_n2406_n2688# 0.200055f
C359 plus.n40 a_n2406_n2688# 0.0916f
C360 plus.t3 a_n2406_n2688# 0.200055f
C361 plus.t2 a_n2406_n2688# 0.200055f
C362 plus.n41 a_n2406_n2688# 0.019767f
C363 plus.n42 a_n2406_n2688# 0.052297f
C364 plus.t21 a_n2406_n2688# 0.200055f
C365 plus.n43 a_n2406_n2688# 0.0916f
C366 plus.t8 a_n2406_n2688# 0.200055f
C367 plus.t5 a_n2406_n2688# 0.200055f
C368 plus.n44 a_n2406_n2688# 0.018155f
C369 plus.t7 a_n2406_n2688# 0.202587f
C370 plus.n45 a_n2406_n2688# 0.11052f
C371 plus.t1 a_n2406_n2688# 0.200055f
C372 plus.n46 a_n2406_n2688# 0.0916f
C373 plus.t9 a_n2406_n2688# 0.200055f
C374 plus.n47 a_n2406_n2688# 0.0916f
C375 plus.n48 a_n2406_n2688# 0.022185f
C376 plus.n49 a_n2406_n2688# 0.114194f
C377 plus.n50 a_n2406_n2688# 0.052297f
C378 plus.n51 a_n2406_n2688# 0.052297f
C379 plus.n52 a_n2406_n2688# 0.021379f
C380 plus.n53 a_n2406_n2688# 0.0916f
C381 plus.n54 a_n2406_n2688# 0.022185f
C382 plus.n55 a_n2406_n2688# 0.0916f
C383 plus.n56 a_n2406_n2688# 0.022185f
C384 plus.n57 a_n2406_n2688# 0.052297f
C385 plus.n58 a_n2406_n2688# 0.052297f
C386 plus.n59 a_n2406_n2688# 0.052297f
C387 plus.n60 a_n2406_n2688# 0.019767f
C388 plus.n61 a_n2406_n2688# 0.0916f
C389 plus.n62 a_n2406_n2688# 0.022185f
C390 plus.n63 a_n2406_n2688# 0.0916f
C391 plus.n64 a_n2406_n2688# 0.022185f
C392 plus.n65 a_n2406_n2688# 0.052297f
C393 plus.n66 a_n2406_n2688# 0.052297f
C394 plus.n67 a_n2406_n2688# 0.052297f
C395 plus.n68 a_n2406_n2688# 0.018155f
C396 plus.n69 a_n2406_n2688# 0.0916f
C397 plus.n70 a_n2406_n2688# 0.022185f
C398 plus.n71 a_n2406_n2688# 0.0916f
C399 plus.n72 a_n2406_n2688# 0.110448f
C400 plus.n73 a_n2406_n2688# 1.60364f
.ends

