* NGSPICE file created from diffpair131.ext - technology: sky130A

.subckt diffpair131 minus drain_right drain_left source plus
X0 a_n1274_n1288# a_n1274_n1288# a_n1274_n1288# a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.6
X1 a_n1274_n1288# a_n1274_n1288# a_n1274_n1288# a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X2 a_n1274_n1288# a_n1274_n1288# a_n1274_n1288# a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X3 source minus drain_right a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X4 source plus drain_left a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X5 source minus drain_right a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X6 drain_right minus source a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X7 drain_left plus source a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X8 source plus drain_left a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.6
X9 a_n1274_n1288# a_n1274_n1288# a_n1274_n1288# a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.6
X10 drain_right minus source a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
X11 drain_left plus source a_n1274_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.6
.ends

