* NGSPICE file created from diffpair636.ext - technology: sky130A

.subckt diffpair636 minus drain_right drain_left source plus
X0 drain_left.t13 plus.t0 source.t16 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X1 drain_right.t13 minus.t0 source.t7 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X2 drain_right.t12 minus.t1 source.t9 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X3 source.t19 plus.t1 drain_left.t12 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X4 a_n2524_n4888# a_n2524_n4888# a_n2524_n4888# a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.8
X5 a_n2524_n4888# a_n2524_n4888# a_n2524_n4888# a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X6 a_n2524_n4888# a_n2524_n4888# a_n2524_n4888# a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X7 a_n2524_n4888# a_n2524_n4888# a_n2524_n4888# a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X8 source.t27 minus.t2 drain_right.t11 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X9 source.t5 minus.t3 drain_right.t10 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X10 source.t22 plus.t2 drain_left.t11 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X11 drain_right.t9 minus.t4 source.t3 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X12 source.t25 minus.t5 drain_right.t8 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X13 source.t11 plus.t3 drain_left.t10 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X14 drain_right.t7 minus.t6 source.t1 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X15 drain_right.t6 minus.t7 source.t8 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X16 source.t10 minus.t8 drain_right.t5 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X17 drain_left.t9 plus.t4 source.t14 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X18 source.t26 minus.t9 drain_right.t4 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X19 source.t4 minus.t10 drain_right.t3 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X20 drain_right.t2 minus.t11 source.t2 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X21 drain_left.t8 plus.t5 source.t17 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X22 source.t21 plus.t6 drain_left.t7 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X23 source.t15 plus.t7 drain_left.t6 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X24 drain_left.t5 plus.t8 source.t23 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X25 drain_left.t4 plus.t9 source.t13 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X26 drain_left.t3 plus.t10 source.t20 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X27 drain_left.t2 plus.t11 source.t24 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X28 source.t12 plus.t12 drain_left.t1 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X29 drain_right.t1 minus.t12 source.t6 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X30 drain_right.t0 minus.t13 source.t0 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X31 drain_left.t0 plus.t13 source.t18 a_n2524_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
R0 plus.n5 plus.t13 675.451
R1 plus.n23 plus.t0 675.451
R2 plus.n16 plus.t5 651.605
R3 plus.n14 plus.t6 651.605
R4 plus.n2 plus.t11 651.605
R5 plus.n9 plus.t7 651.605
R6 plus.n8 plus.t8 651.605
R7 plus.n4 plus.t12 651.605
R8 plus.n34 plus.t4 651.605
R9 plus.n32 plus.t1 651.605
R10 plus.n20 plus.t9 651.605
R11 plus.n27 plus.t2 651.605
R12 plus.n26 plus.t10 651.605
R13 plus.n22 plus.t3 651.605
R14 plus.n7 plus.n6 161.3
R15 plus.n13 plus.n12 161.3
R16 plus.n14 plus.n1 161.3
R17 plus.n15 plus.n0 161.3
R18 plus.n17 plus.n16 161.3
R19 plus.n25 plus.n24 161.3
R20 plus.n31 plus.n30 161.3
R21 plus.n32 plus.n19 161.3
R22 plus.n33 plus.n18 161.3
R23 plus.n35 plus.n34 161.3
R24 plus.n8 plus.n3 80.6037
R25 plus.n10 plus.n9 80.6037
R26 plus.n11 plus.n2 80.6037
R27 plus.n26 plus.n21 80.6037
R28 plus.n28 plus.n27 80.6037
R29 plus.n29 plus.n20 80.6037
R30 plus.n9 plus.n2 48.2005
R31 plus.n9 plus.n8 48.2005
R32 plus.n27 plus.n20 48.2005
R33 plus.n27 plus.n26 48.2005
R34 plus.n24 plus.n23 44.9119
R35 plus.n6 plus.n5 44.9119
R36 plus plus.n35 35.8191
R37 plus.n16 plus.n15 35.055
R38 plus.n34 plus.n33 35.055
R39 plus.n13 plus.n2 32.1338
R40 plus.n8 plus.n7 32.1338
R41 plus.n31 plus.n20 32.1338
R42 plus.n26 plus.n25 32.1338
R43 plus.n23 plus.n22 17.739
R44 plus.n5 plus.n4 17.739
R45 plus.n14 plus.n13 16.0672
R46 plus.n7 plus.n4 16.0672
R47 plus.n32 plus.n31 16.0672
R48 plus.n25 plus.n22 16.0672
R49 plus plus.n17 15.4001
R50 plus.n15 plus.n14 13.146
R51 plus.n33 plus.n32 13.146
R52 plus.n10 plus.n3 0.380177
R53 plus.n11 plus.n10 0.380177
R54 plus.n29 plus.n28 0.380177
R55 plus.n28 plus.n21 0.380177
R56 plus.n6 plus.n3 0.285035
R57 plus.n12 plus.n11 0.285035
R58 plus.n30 plus.n29 0.285035
R59 plus.n24 plus.n21 0.285035
R60 plus.n12 plus.n1 0.189894
R61 plus.n1 plus.n0 0.189894
R62 plus.n17 plus.n0 0.189894
R63 plus.n35 plus.n18 0.189894
R64 plus.n19 plus.n18 0.189894
R65 plus.n30 plus.n19 0.189894
R66 source.n0 source.t17 44.1297
R67 source.n7 source.t8 44.1296
R68 source.n27 source.t6 44.1295
R69 source.n20 source.t16 44.1295
R70 source.n2 source.n1 43.1397
R71 source.n4 source.n3 43.1397
R72 source.n6 source.n5 43.1397
R73 source.n9 source.n8 43.1397
R74 source.n11 source.n10 43.1397
R75 source.n13 source.n12 43.1397
R76 source.n26 source.n25 43.1396
R77 source.n24 source.n23 43.1396
R78 source.n22 source.n21 43.1396
R79 source.n19 source.n18 43.1396
R80 source.n17 source.n16 43.1396
R81 source.n15 source.n14 43.1396
R82 source.n15 source.n13 29.2966
R83 source.n28 source.n0 22.5725
R84 source.n28 source.n27 5.7505
R85 source.n25 source.t7 0.9905
R86 source.n25 source.t27 0.9905
R87 source.n23 source.t0 0.9905
R88 source.n23 source.t5 0.9905
R89 source.n21 source.t9 0.9905
R90 source.n21 source.t10 0.9905
R91 source.n18 source.t20 0.9905
R92 source.n18 source.t11 0.9905
R93 source.n16 source.t13 0.9905
R94 source.n16 source.t22 0.9905
R95 source.n14 source.t14 0.9905
R96 source.n14 source.t19 0.9905
R97 source.n1 source.t24 0.9905
R98 source.n1 source.t21 0.9905
R99 source.n3 source.t23 0.9905
R100 source.n3 source.t15 0.9905
R101 source.n5 source.t18 0.9905
R102 source.n5 source.t12 0.9905
R103 source.n8 source.t3 0.9905
R104 source.n8 source.t25 0.9905
R105 source.n10 source.t2 0.9905
R106 source.n10 source.t4 0.9905
R107 source.n12 source.t1 0.9905
R108 source.n12 source.t26 0.9905
R109 source.n13 source.n11 0.974638
R110 source.n11 source.n9 0.974638
R111 source.n9 source.n7 0.974638
R112 source.n6 source.n4 0.974638
R113 source.n4 source.n2 0.974638
R114 source.n2 source.n0 0.974638
R115 source.n17 source.n15 0.974638
R116 source.n19 source.n17 0.974638
R117 source.n20 source.n19 0.974638
R118 source.n24 source.n22 0.974638
R119 source.n26 source.n24 0.974638
R120 source.n27 source.n26 0.974638
R121 source.n7 source.n6 0.957397
R122 source.n22 source.n20 0.957397
R123 source source.n28 0.188
R124 drain_left.n7 drain_left.t0 61.7825
R125 drain_left.n1 drain_left.t9 61.7824
R126 drain_left.n4 drain_left.n2 60.7925
R127 drain_left.n11 drain_left.n10 59.8185
R128 drain_left.n9 drain_left.n8 59.8185
R129 drain_left.n7 drain_left.n6 59.8185
R130 drain_left.n4 drain_left.n3 59.8184
R131 drain_left.n1 drain_left.n0 59.8184
R132 drain_left drain_left.n5 39.029
R133 drain_left drain_left.n11 6.62735
R134 drain_left.n2 drain_left.t10 0.9905
R135 drain_left.n2 drain_left.t13 0.9905
R136 drain_left.n3 drain_left.t11 0.9905
R137 drain_left.n3 drain_left.t3 0.9905
R138 drain_left.n0 drain_left.t12 0.9905
R139 drain_left.n0 drain_left.t4 0.9905
R140 drain_left.n10 drain_left.t7 0.9905
R141 drain_left.n10 drain_left.t8 0.9905
R142 drain_left.n8 drain_left.t6 0.9905
R143 drain_left.n8 drain_left.t2 0.9905
R144 drain_left.n6 drain_left.t1 0.9905
R145 drain_left.n6 drain_left.t5 0.9905
R146 drain_left.n9 drain_left.n7 0.974638
R147 drain_left.n11 drain_left.n9 0.974638
R148 drain_left.n5 drain_left.n1 0.675757
R149 drain_left.n5 drain_left.n4 0.188688
R150 minus.n5 minus.t7 675.451
R151 minus.n23 minus.t1 675.451
R152 minus.n4 minus.t5 651.605
R153 minus.n8 minus.t4 651.605
R154 minus.n9 minus.t10 651.605
R155 minus.n10 minus.t11 651.605
R156 minus.n14 minus.t9 651.605
R157 minus.n16 minus.t6 651.605
R158 minus.n22 minus.t8 651.605
R159 minus.n26 minus.t13 651.605
R160 minus.n27 minus.t3 651.605
R161 minus.n28 minus.t0 651.605
R162 minus.n32 minus.t2 651.605
R163 minus.n34 minus.t12 651.605
R164 minus.n17 minus.n16 161.3
R165 minus.n15 minus.n0 161.3
R166 minus.n14 minus.n13 161.3
R167 minus.n12 minus.n1 161.3
R168 minus.n6 minus.n3 161.3
R169 minus.n35 minus.n34 161.3
R170 minus.n33 minus.n18 161.3
R171 minus.n32 minus.n31 161.3
R172 minus.n30 minus.n19 161.3
R173 minus.n24 minus.n21 161.3
R174 minus.n11 minus.n10 80.6037
R175 minus.n9 minus.n2 80.6037
R176 minus.n8 minus.n7 80.6037
R177 minus.n29 minus.n28 80.6037
R178 minus.n27 minus.n20 80.6037
R179 minus.n26 minus.n25 80.6037
R180 minus.n9 minus.n8 48.2005
R181 minus.n10 minus.n9 48.2005
R182 minus.n27 minus.n26 48.2005
R183 minus.n28 minus.n27 48.2005
R184 minus.n36 minus.n17 44.9683
R185 minus.n6 minus.n5 44.9119
R186 minus.n24 minus.n23 44.9119
R187 minus.n16 minus.n15 35.055
R188 minus.n34 minus.n33 35.055
R189 minus.n8 minus.n3 32.1338
R190 minus.n10 minus.n1 32.1338
R191 minus.n26 minus.n21 32.1338
R192 minus.n28 minus.n19 32.1338
R193 minus.n5 minus.n4 17.739
R194 minus.n23 minus.n22 17.739
R195 minus.n4 minus.n3 16.0672
R196 minus.n14 minus.n1 16.0672
R197 minus.n22 minus.n21 16.0672
R198 minus.n32 minus.n19 16.0672
R199 minus.n15 minus.n14 13.146
R200 minus.n33 minus.n32 13.146
R201 minus.n36 minus.n35 6.72588
R202 minus.n11 minus.n2 0.380177
R203 minus.n7 minus.n2 0.380177
R204 minus.n25 minus.n20 0.380177
R205 minus.n29 minus.n20 0.380177
R206 minus.n12 minus.n11 0.285035
R207 minus.n7 minus.n6 0.285035
R208 minus.n25 minus.n24 0.285035
R209 minus.n30 minus.n29 0.285035
R210 minus.n17 minus.n0 0.189894
R211 minus.n13 minus.n0 0.189894
R212 minus.n13 minus.n12 0.189894
R213 minus.n31 minus.n30 0.189894
R214 minus.n31 minus.n18 0.189894
R215 minus.n35 minus.n18 0.189894
R216 minus minus.n36 0.188
R217 drain_right.n1 drain_right.t12 61.7824
R218 drain_right.n11 drain_right.t7 60.8084
R219 drain_right.n8 drain_right.n6 60.7926
R220 drain_right.n4 drain_right.n2 60.7925
R221 drain_right.n8 drain_right.n7 59.8185
R222 drain_right.n10 drain_right.n9 59.8185
R223 drain_right.n4 drain_right.n3 59.8184
R224 drain_right.n1 drain_right.n0 59.8184
R225 drain_right drain_right.n5 38.4757
R226 drain_right drain_right.n11 6.14028
R227 drain_right.n2 drain_right.t11 0.9905
R228 drain_right.n2 drain_right.t1 0.9905
R229 drain_right.n3 drain_right.t10 0.9905
R230 drain_right.n3 drain_right.t13 0.9905
R231 drain_right.n0 drain_right.t5 0.9905
R232 drain_right.n0 drain_right.t0 0.9905
R233 drain_right.n6 drain_right.t8 0.9905
R234 drain_right.n6 drain_right.t6 0.9905
R235 drain_right.n7 drain_right.t3 0.9905
R236 drain_right.n7 drain_right.t9 0.9905
R237 drain_right.n9 drain_right.t4 0.9905
R238 drain_right.n9 drain_right.t2 0.9905
R239 drain_right.n11 drain_right.n10 0.974638
R240 drain_right.n10 drain_right.n8 0.974638
R241 drain_right.n5 drain_right.n1 0.675757
R242 drain_right.n5 drain_right.n4 0.188688
C0 plus source 15.572701f
C1 minus source 15.557799f
C2 drain_left source 26.9903f
C3 source drain_right 26.9801f
C4 plus minus 7.76813f
C5 plus drain_left 16.0872f
C6 plus drain_right 0.409473f
C7 minus drain_left 0.173289f
C8 minus drain_right 15.8411f
C9 drain_left drain_right 1.31943f
C10 drain_right a_n2524_n4888# 9.86671f
C11 drain_left a_n2524_n4888# 10.24104f
C12 source a_n2524_n4888# 9.74464f
C13 minus a_n2524_n4888# 10.573273f
C14 plus a_n2524_n4888# 12.6287f
C15 drain_right.t12 a_n2524_n4888# 4.49979f
C16 drain_right.t5 a_n2524_n4888# 0.384359f
C17 drain_right.t0 a_n2524_n4888# 0.384359f
C18 drain_right.n0 a_n2524_n4888# 3.5139f
C19 drain_right.n1 a_n2524_n4888# 0.689027f
C20 drain_right.t11 a_n2524_n4888# 0.384359f
C21 drain_right.t1 a_n2524_n4888# 0.384359f
C22 drain_right.n2 a_n2524_n4888# 3.51979f
C23 drain_right.t10 a_n2524_n4888# 0.384359f
C24 drain_right.t13 a_n2524_n4888# 0.384359f
C25 drain_right.n3 a_n2524_n4888# 3.5139f
C26 drain_right.n4 a_n2524_n4888# 0.661097f
C27 drain_right.n5 a_n2524_n4888# 1.81677f
C28 drain_right.t8 a_n2524_n4888# 0.384359f
C29 drain_right.t6 a_n2524_n4888# 0.384359f
C30 drain_right.n6 a_n2524_n4888# 3.51979f
C31 drain_right.t3 a_n2524_n4888# 0.384359f
C32 drain_right.t9 a_n2524_n4888# 0.384359f
C33 drain_right.n7 a_n2524_n4888# 3.51389f
C34 drain_right.n8 a_n2524_n4888# 0.719701f
C35 drain_right.t4 a_n2524_n4888# 0.384359f
C36 drain_right.t2 a_n2524_n4888# 0.384359f
C37 drain_right.n9 a_n2524_n4888# 3.51389f
C38 drain_right.n10 a_n2524_n4888# 0.357899f
C39 drain_right.t7 a_n2524_n4888# 4.49414f
C40 drain_right.n11 a_n2524_n4888# 0.587972f
C41 minus.n0 a_n2524_n4888# 0.038637f
C42 minus.n1 a_n2524_n4888# 0.008768f
C43 minus.t9 a_n2524_n4888# 1.75065f
C44 minus.n2 a_n2524_n4888# 0.077274f
C45 minus.n3 a_n2524_n4888# 0.008768f
C46 minus.t4 a_n2524_n4888# 1.75065f
C47 minus.t7 a_n2524_n4888# 1.77366f
C48 minus.t5 a_n2524_n4888# 1.75065f
C49 minus.n4 a_n2524_n4888# 0.654065f
C50 minus.n5 a_n2524_n4888# 0.632049f
C51 minus.n6 a_n2524_n4888# 0.18044f
C52 minus.n7 a_n2524_n4888# 0.064355f
C53 minus.n8 a_n2524_n4888# 0.658523f
C54 minus.t10 a_n2524_n4888# 1.75065f
C55 minus.n9 a_n2524_n4888# 0.661144f
C56 minus.t11 a_n2524_n4888# 1.75065f
C57 minus.n10 a_n2524_n4888# 0.658523f
C58 minus.n11 a_n2524_n4888# 0.064355f
C59 minus.n12 a_n2524_n4888# 0.051556f
C60 minus.n13 a_n2524_n4888# 0.038637f
C61 minus.n14 a_n2524_n4888# 0.649279f
C62 minus.n15 a_n2524_n4888# 0.008768f
C63 minus.t6 a_n2524_n4888# 1.75065f
C64 minus.n16 a_n2524_n4888# 0.650232f
C65 minus.n17 a_n2524_n4888# 1.89515f
C66 minus.n18 a_n2524_n4888# 0.038637f
C67 minus.n19 a_n2524_n4888# 0.008768f
C68 minus.n20 a_n2524_n4888# 0.077274f
C69 minus.n21 a_n2524_n4888# 0.008768f
C70 minus.t1 a_n2524_n4888# 1.77366f
C71 minus.t8 a_n2524_n4888# 1.75065f
C72 minus.n22 a_n2524_n4888# 0.654065f
C73 minus.n23 a_n2524_n4888# 0.632049f
C74 minus.n24 a_n2524_n4888# 0.18044f
C75 minus.n25 a_n2524_n4888# 0.064355f
C76 minus.t13 a_n2524_n4888# 1.75065f
C77 minus.n26 a_n2524_n4888# 0.658523f
C78 minus.t3 a_n2524_n4888# 1.75065f
C79 minus.n27 a_n2524_n4888# 0.661144f
C80 minus.t0 a_n2524_n4888# 1.75065f
C81 minus.n28 a_n2524_n4888# 0.658523f
C82 minus.n29 a_n2524_n4888# 0.064355f
C83 minus.n30 a_n2524_n4888# 0.051556f
C84 minus.n31 a_n2524_n4888# 0.038637f
C85 minus.t2 a_n2524_n4888# 1.75065f
C86 minus.n32 a_n2524_n4888# 0.649279f
C87 minus.n33 a_n2524_n4888# 0.008768f
C88 minus.t12 a_n2524_n4888# 1.75065f
C89 minus.n34 a_n2524_n4888# 0.650232f
C90 minus.n35 a_n2524_n4888# 0.272945f
C91 minus.n36 a_n2524_n4888# 2.24067f
C92 drain_left.t9 a_n2524_n4888# 4.52128f
C93 drain_left.t12 a_n2524_n4888# 0.386195f
C94 drain_left.t4 a_n2524_n4888# 0.386195f
C95 drain_left.n0 a_n2524_n4888# 3.53068f
C96 drain_left.n1 a_n2524_n4888# 0.692317f
C97 drain_left.t10 a_n2524_n4888# 0.386195f
C98 drain_left.t13 a_n2524_n4888# 0.386195f
C99 drain_left.n2 a_n2524_n4888# 3.5366f
C100 drain_left.t11 a_n2524_n4888# 0.386195f
C101 drain_left.t3 a_n2524_n4888# 0.386195f
C102 drain_left.n3 a_n2524_n4888# 3.53068f
C103 drain_left.n4 a_n2524_n4888# 0.664255f
C104 drain_left.n5 a_n2524_n4888# 1.87583f
C105 drain_left.t0 a_n2524_n4888# 4.52129f
C106 drain_left.t1 a_n2524_n4888# 0.386195f
C107 drain_left.t5 a_n2524_n4888# 0.386195f
C108 drain_left.n6 a_n2524_n4888# 3.53068f
C109 drain_left.n7 a_n2524_n4888# 0.714999f
C110 drain_left.t6 a_n2524_n4888# 0.386195f
C111 drain_left.t2 a_n2524_n4888# 0.386195f
C112 drain_left.n8 a_n2524_n4888# 3.53068f
C113 drain_left.n9 a_n2524_n4888# 0.359608f
C114 drain_left.t7 a_n2524_n4888# 0.386195f
C115 drain_left.t8 a_n2524_n4888# 0.386195f
C116 drain_left.n10 a_n2524_n4888# 3.53068f
C117 drain_left.n11 a_n2524_n4888# 0.578721f
C118 source.t17 a_n2524_n4888# 4.53456f
C119 source.n0 a_n2524_n4888# 1.98364f
C120 source.t24 a_n2524_n4888# 0.396781f
C121 source.t21 a_n2524_n4888# 0.396781f
C122 source.n1 a_n2524_n4888# 3.54739f
C123 source.n2 a_n2524_n4888# 0.415404f
C124 source.t23 a_n2524_n4888# 0.396781f
C125 source.t15 a_n2524_n4888# 0.396781f
C126 source.n3 a_n2524_n4888# 3.54739f
C127 source.n4 a_n2524_n4888# 0.415404f
C128 source.t18 a_n2524_n4888# 0.396781f
C129 source.t12 a_n2524_n4888# 0.396781f
C130 source.n5 a_n2524_n4888# 3.54739f
C131 source.n6 a_n2524_n4888# 0.414009f
C132 source.t8 a_n2524_n4888# 4.53457f
C133 source.n7 a_n2524_n4888# 0.508957f
C134 source.t3 a_n2524_n4888# 0.396781f
C135 source.t25 a_n2524_n4888# 0.396781f
C136 source.n8 a_n2524_n4888# 3.54739f
C137 source.n9 a_n2524_n4888# 0.415404f
C138 source.t2 a_n2524_n4888# 0.396781f
C139 source.t4 a_n2524_n4888# 0.396781f
C140 source.n10 a_n2524_n4888# 3.54739f
C141 source.n11 a_n2524_n4888# 0.415404f
C142 source.t1 a_n2524_n4888# 0.396781f
C143 source.t26 a_n2524_n4888# 0.396781f
C144 source.n12 a_n2524_n4888# 3.54739f
C145 source.n13 a_n2524_n4888# 2.42719f
C146 source.t14 a_n2524_n4888# 0.396781f
C147 source.t19 a_n2524_n4888# 0.396781f
C148 source.n14 a_n2524_n4888# 3.54739f
C149 source.n15 a_n2524_n4888# 2.42718f
C150 source.t13 a_n2524_n4888# 0.396781f
C151 source.t22 a_n2524_n4888# 0.396781f
C152 source.n16 a_n2524_n4888# 3.54739f
C153 source.n17 a_n2524_n4888# 0.415397f
C154 source.t20 a_n2524_n4888# 0.396781f
C155 source.t11 a_n2524_n4888# 0.396781f
C156 source.n18 a_n2524_n4888# 3.54739f
C157 source.n19 a_n2524_n4888# 0.415397f
C158 source.t16 a_n2524_n4888# 4.53454f
C159 source.n20 a_n2524_n4888# 0.508982f
C160 source.t9 a_n2524_n4888# 0.396781f
C161 source.t10 a_n2524_n4888# 0.396781f
C162 source.n21 a_n2524_n4888# 3.54739f
C163 source.n22 a_n2524_n4888# 0.414002f
C164 source.t0 a_n2524_n4888# 0.396781f
C165 source.t5 a_n2524_n4888# 0.396781f
C166 source.n23 a_n2524_n4888# 3.54739f
C167 source.n24 a_n2524_n4888# 0.415397f
C168 source.t7 a_n2524_n4888# 0.396781f
C169 source.t27 a_n2524_n4888# 0.396781f
C170 source.n25 a_n2524_n4888# 3.54739f
C171 source.n26 a_n2524_n4888# 0.415397f
C172 source.t6 a_n2524_n4888# 4.53454f
C173 source.n27 a_n2524_n4888# 0.638779f
C174 source.n28 a_n2524_n4888# 2.28214f
C175 plus.n0 a_n2524_n4888# 0.03901f
C176 plus.t5 a_n2524_n4888# 1.76757f
C177 plus.t6 a_n2524_n4888# 1.76757f
C178 plus.n1 a_n2524_n4888# 0.03901f
C179 plus.t11 a_n2524_n4888# 1.76757f
C180 plus.n2 a_n2524_n4888# 0.664888f
C181 plus.n3 a_n2524_n4888# 0.064977f
C182 plus.t7 a_n2524_n4888# 1.76757f
C183 plus.t8 a_n2524_n4888# 1.76757f
C184 plus.t12 a_n2524_n4888# 1.76757f
C185 plus.n4 a_n2524_n4888# 0.660387f
C186 plus.t13 a_n2524_n4888# 1.7908f
C187 plus.n5 a_n2524_n4888# 0.638158f
C188 plus.n6 a_n2524_n4888# 0.182184f
C189 plus.n7 a_n2524_n4888# 0.008852f
C190 plus.n8 a_n2524_n4888# 0.664888f
C191 plus.n9 a_n2524_n4888# 0.667534f
C192 plus.n10 a_n2524_n4888# 0.078021f
C193 plus.n11 a_n2524_n4888# 0.064977f
C194 plus.n12 a_n2524_n4888# 0.052054f
C195 plus.n13 a_n2524_n4888# 0.008852f
C196 plus.n14 a_n2524_n4888# 0.655555f
C197 plus.n15 a_n2524_n4888# 0.008852f
C198 plus.n16 a_n2524_n4888# 0.656517f
C199 plus.n17 a_n2524_n4888# 0.612528f
C200 plus.n18 a_n2524_n4888# 0.03901f
C201 plus.t4 a_n2524_n4888# 1.76757f
C202 plus.n19 a_n2524_n4888# 0.03901f
C203 plus.t1 a_n2524_n4888# 1.76757f
C204 plus.t9 a_n2524_n4888# 1.76757f
C205 plus.n20 a_n2524_n4888# 0.664888f
C206 plus.n21 a_n2524_n4888# 0.064977f
C207 plus.t2 a_n2524_n4888# 1.76757f
C208 plus.t10 a_n2524_n4888# 1.76757f
C209 plus.t3 a_n2524_n4888# 1.76757f
C210 plus.n22 a_n2524_n4888# 0.660387f
C211 plus.t0 a_n2524_n4888# 1.7908f
C212 plus.n23 a_n2524_n4888# 0.638158f
C213 plus.n24 a_n2524_n4888# 0.182184f
C214 plus.n25 a_n2524_n4888# 0.008852f
C215 plus.n26 a_n2524_n4888# 0.664888f
C216 plus.n27 a_n2524_n4888# 0.667534f
C217 plus.n28 a_n2524_n4888# 0.078021f
C218 plus.n29 a_n2524_n4888# 0.064977f
C219 plus.n30 a_n2524_n4888# 0.052054f
C220 plus.n31 a_n2524_n4888# 0.008852f
C221 plus.n32 a_n2524_n4888# 0.655555f
C222 plus.n33 a_n2524_n4888# 0.008852f
C223 plus.n34 a_n2524_n4888# 0.656517f
C224 plus.n35 a_n2524_n4888# 1.53258f
.ends

