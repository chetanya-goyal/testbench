* NGSPICE file created from diffpair101.ext - technology: sky130A

.subckt diffpair101 minus drain_right drain_left source plus
X0 source minus drain_right a_n1064_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X1 drain_right minus source a_n1064_n1292# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X2 source plus drain_left a_n1064_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X3 a_n1064_n1292# a_n1064_n1292# a_n1064_n1292# a_n1064_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.25
X4 drain_left plus source a_n1064_n1292# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X5 a_n1064_n1292# a_n1064_n1292# a_n1064_n1292# a_n1064_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X6 drain_left plus source a_n1064_n1292# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X7 source minus drain_right a_n1064_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X8 a_n1064_n1292# a_n1064_n1292# a_n1064_n1292# a_n1064_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X9 source plus drain_left a_n1064_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X10 drain_right minus source a_n1064_n1292# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X11 a_n1064_n1292# a_n1064_n1292# a_n1064_n1292# a_n1064_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
.ends

