* NGSPICE file created from diffpair451.ext - technology: sky130A

.subckt diffpair451 minus drain_right drain_left source plus
X0 a_n1274_n3288# a_n1274_n3288# a_n1274_n3288# a_n1274_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.6
X1 drain_right minus source a_n1274_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.6
X2 a_n1274_n3288# a_n1274_n3288# a_n1274_n3288# a_n1274_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.6
X3 a_n1274_n3288# a_n1274_n3288# a_n1274_n3288# a_n1274_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.6
X4 source plus drain_left a_n1274_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.6
X5 source minus drain_right a_n1274_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.6
X6 a_n1274_n3288# a_n1274_n3288# a_n1274_n3288# a_n1274_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.6
X7 source minus drain_right a_n1274_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.6
X8 drain_right minus source a_n1274_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.6
X9 drain_left plus source a_n1274_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.6
X10 source plus drain_left a_n1274_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.6
X11 drain_left plus source a_n1274_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.6
.ends

