* NGSPICE file created from diffpair213.ext - technology: sky130A

.subckt diffpair213 minus drain_right drain_left source plus
X0 a_n1646_n1488# a_n1646_n1488# a_n1646_n1488# a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.6
X1 source.t15 minus.t0 drain_right.t2 a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X2 a_n1646_n1488# a_n1646_n1488# a_n1646_n1488# a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X3 drain_right.t3 minus.t1 source.t14 a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X4 drain_left.t7 plus.t0 source.t4 a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X5 source.t13 minus.t2 drain_right.t0 a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X6 drain_right.t4 minus.t3 source.t12 a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X7 source.t5 plus.t1 drain_left.t6 a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X8 a_n1646_n1488# a_n1646_n1488# a_n1646_n1488# a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X9 drain_left.t5 plus.t2 source.t2 a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X10 source.t11 minus.t4 drain_right.t5 a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X11 drain_right.t1 minus.t5 source.t10 a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X12 source.t3 plus.t3 drain_left.t4 a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X13 drain_right.t6 minus.t6 source.t9 a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X14 source.t8 minus.t7 drain_right.t7 a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X15 drain_left.t3 plus.t4 source.t1 a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X16 source.t0 plus.t5 drain_left.t2 a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X17 drain_left.t1 plus.t6 source.t7 a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X18 source.t6 plus.t7 drain_left.t0 a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X19 a_n1646_n1488# a_n1646_n1488# a_n1646_n1488# a_n1646_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
R0 minus.n1 minus.t6 212.793
R1 minus.n7 minus.t7 212.793
R2 minus.n2 minus.t4 185.972
R3 minus.n3 minus.t3 185.972
R4 minus.n4 minus.t2 185.972
R5 minus.n8 minus.t1 185.972
R6 minus.n9 minus.t0 185.972
R7 minus.n10 minus.t5 185.972
R8 minus.n5 minus.n4 161.3
R9 minus.n11 minus.n10 161.3
R10 minus.n3 minus.n0 80.6037
R11 minus.n9 minus.n6 80.6037
R12 minus.n3 minus.n2 48.2005
R13 minus.n4 minus.n3 48.2005
R14 minus.n9 minus.n8 48.2005
R15 minus.n10 minus.n9 48.2005
R16 minus.n1 minus.n0 45.2318
R17 minus.n7 minus.n6 45.2318
R18 minus.n12 minus.n5 28.652
R19 minus.n2 minus.n1 13.3799
R20 minus.n8 minus.n7 13.3799
R21 minus.n12 minus.n11 6.61414
R22 minus.n5 minus.n0 0.285035
R23 minus.n11 minus.n6 0.285035
R24 minus minus.n12 0.188
R25 drain_right.n5 drain_right.n3 80.5748
R26 drain_right.n2 drain_right.n1 80.1185
R27 drain_right.n2 drain_right.n0 80.1185
R28 drain_right.n5 drain_right.n4 79.7731
R29 drain_right drain_right.n2 22.8017
R30 drain_right.n1 drain_right.t2 6.6005
R31 drain_right.n1 drain_right.t1 6.6005
R32 drain_right.n0 drain_right.t7 6.6005
R33 drain_right.n0 drain_right.t3 6.6005
R34 drain_right.n3 drain_right.t5 6.6005
R35 drain_right.n3 drain_right.t6 6.6005
R36 drain_right.n4 drain_right.t0 6.6005
R37 drain_right.n4 drain_right.t4 6.6005
R38 drain_right drain_right.n5 6.45494
R39 source.n0 source.t2 69.6943
R40 source.n3 source.t0 69.6943
R41 source.n4 source.t9 69.6943
R42 source.n7 source.t13 69.6943
R43 source.n15 source.t10 69.6942
R44 source.n12 source.t8 69.6942
R45 source.n11 source.t4 69.6942
R46 source.n8 source.t5 69.6942
R47 source.n2 source.n1 63.0943
R48 source.n6 source.n5 63.0943
R49 source.n14 source.n13 63.0942
R50 source.n10 source.n9 63.0942
R51 source.n8 source.n7 15.2713
R52 source.n16 source.n0 9.60747
R53 source.n13 source.t14 6.6005
R54 source.n13 source.t15 6.6005
R55 source.n9 source.t7 6.6005
R56 source.n9 source.t6 6.6005
R57 source.n1 source.t1 6.6005
R58 source.n1 source.t3 6.6005
R59 source.n5 source.t12 6.6005
R60 source.n5 source.t11 6.6005
R61 source.n16 source.n15 5.66429
R62 source.n7 source.n6 0.802224
R63 source.n6 source.n4 0.802224
R64 source.n3 source.n2 0.802224
R65 source.n2 source.n0 0.802224
R66 source.n10 source.n8 0.802224
R67 source.n11 source.n10 0.802224
R68 source.n14 source.n12 0.802224
R69 source.n15 source.n14 0.802224
R70 source.n4 source.n3 0.470328
R71 source.n12 source.n11 0.470328
R72 source source.n16 0.188
R73 plus.n1 plus.t5 212.793
R74 plus.n7 plus.t0 212.793
R75 plus.n4 plus.t2 185.972
R76 plus.n3 plus.t3 185.972
R77 plus.n2 plus.t4 185.972
R78 plus.n10 plus.t1 185.972
R79 plus.n9 plus.t6 185.972
R80 plus.n8 plus.t7 185.972
R81 plus.n5 plus.n4 161.3
R82 plus.n11 plus.n10 161.3
R83 plus.n3 plus.n0 80.6037
R84 plus.n9 plus.n6 80.6037
R85 plus.n4 plus.n3 48.2005
R86 plus.n3 plus.n2 48.2005
R87 plus.n10 plus.n9 48.2005
R88 plus.n9 plus.n8 48.2005
R89 plus.n1 plus.n0 45.2318
R90 plus.n7 plus.n6 45.2318
R91 plus plus.n11 25.9422
R92 plus.n2 plus.n1 13.3799
R93 plus.n8 plus.n7 13.3799
R94 plus plus.n5 8.84898
R95 plus.n5 plus.n0 0.285035
R96 plus.n11 plus.n6 0.285035
R97 drain_left.n5 drain_left.n3 80.5748
R98 drain_left.n2 drain_left.n1 80.1185
R99 drain_left.n2 drain_left.n0 80.1185
R100 drain_left.n5 drain_left.n4 79.7731
R101 drain_left drain_left.n2 23.3549
R102 drain_left.n1 drain_left.t0 6.6005
R103 drain_left.n1 drain_left.t7 6.6005
R104 drain_left.n0 drain_left.t6 6.6005
R105 drain_left.n0 drain_left.t1 6.6005
R106 drain_left.n4 drain_left.t4 6.6005
R107 drain_left.n4 drain_left.t5 6.6005
R108 drain_left.n3 drain_left.t2 6.6005
R109 drain_left.n3 drain_left.t3 6.6005
R110 drain_left drain_left.n5 6.45494
C0 drain_right minus 1.55428f
C1 minus plus 3.53537f
C2 drain_right drain_left 0.775958f
C3 plus drain_left 1.71268f
C4 source minus 1.71759f
C5 drain_right plus 0.318271f
C6 source drain_left 4.5659f
C7 drain_right source 4.56704f
C8 source plus 1.73158f
C9 minus drain_left 0.17632f
C10 drain_right a_n1646_n1488# 3.40555f
C11 drain_left a_n1646_n1488# 3.61271f
C12 source a_n1646_n1488# 3.61498f
C13 minus a_n1646_n1488# 5.629075f
C14 plus a_n1646_n1488# 6.176324f
C15 drain_left.t6 a_n1646_n1488# 0.046486f
C16 drain_left.t1 a_n1646_n1488# 0.046486f
C17 drain_left.n0 a_n1646_n1488# 0.336282f
C18 drain_left.t0 a_n1646_n1488# 0.046486f
C19 drain_left.t7 a_n1646_n1488# 0.046486f
C20 drain_left.n1 a_n1646_n1488# 0.336282f
C21 drain_left.n2 a_n1646_n1488# 1.0437f
C22 drain_left.t2 a_n1646_n1488# 0.046486f
C23 drain_left.t3 a_n1646_n1488# 0.046486f
C24 drain_left.n3 a_n1646_n1488# 0.337903f
C25 drain_left.t4 a_n1646_n1488# 0.046486f
C26 drain_left.t5 a_n1646_n1488# 0.046486f
C27 drain_left.n4 a_n1646_n1488# 0.335254f
C28 drain_left.n5 a_n1646_n1488# 0.692784f
C29 plus.n0 a_n1646_n1488# 0.122456f
C30 plus.t2 a_n1646_n1488# 0.135551f
C31 plus.t3 a_n1646_n1488# 0.135551f
C32 plus.t4 a_n1646_n1488# 0.135551f
C33 plus.t5 a_n1646_n1488# 0.145664f
C34 plus.n1 a_n1646_n1488# 0.0708f
C35 plus.n2 a_n1646_n1488# 0.085859f
C36 plus.n3 a_n1646_n1488# 0.085859f
C37 plus.n4 a_n1646_n1488# 0.08016f
C38 plus.n5 a_n1646_n1488# 0.203067f
C39 plus.n6 a_n1646_n1488# 0.122456f
C40 plus.t1 a_n1646_n1488# 0.135551f
C41 plus.t6 a_n1646_n1488# 0.135551f
C42 plus.t0 a_n1646_n1488# 0.145664f
C43 plus.n7 a_n1646_n1488# 0.0708f
C44 plus.t7 a_n1646_n1488# 0.135551f
C45 plus.n8 a_n1646_n1488# 0.085859f
C46 plus.n9 a_n1646_n1488# 0.085859f
C47 plus.n10 a_n1646_n1488# 0.08016f
C48 plus.n11 a_n1646_n1488# 0.579752f
C49 source.t2 a_n1646_n1488# 0.355984f
C50 source.n0 a_n1646_n1488# 0.512169f
C51 source.t1 a_n1646_n1488# 0.04287f
C52 source.t3 a_n1646_n1488# 0.04287f
C53 source.n1 a_n1646_n1488# 0.27182f
C54 source.n2 a_n1646_n1488# 0.250959f
C55 source.t0 a_n1646_n1488# 0.355984f
C56 source.n3 a_n1646_n1488# 0.264374f
C57 source.t9 a_n1646_n1488# 0.355984f
C58 source.n4 a_n1646_n1488# 0.264374f
C59 source.t12 a_n1646_n1488# 0.04287f
C60 source.t11 a_n1646_n1488# 0.04287f
C61 source.n5 a_n1646_n1488# 0.27182f
C62 source.n6 a_n1646_n1488# 0.250959f
C63 source.t13 a_n1646_n1488# 0.355984f
C64 source.n7 a_n1646_n1488# 0.704314f
C65 source.t5 a_n1646_n1488# 0.355982f
C66 source.n8 a_n1646_n1488# 0.704316f
C67 source.t7 a_n1646_n1488# 0.04287f
C68 source.t6 a_n1646_n1488# 0.04287f
C69 source.n9 a_n1646_n1488# 0.271818f
C70 source.n10 a_n1646_n1488# 0.250961f
C71 source.t4 a_n1646_n1488# 0.355982f
C72 source.n11 a_n1646_n1488# 0.264375f
C73 source.t8 a_n1646_n1488# 0.355982f
C74 source.n12 a_n1646_n1488# 0.264375f
C75 source.t14 a_n1646_n1488# 0.04287f
C76 source.t15 a_n1646_n1488# 0.04287f
C77 source.n13 a_n1646_n1488# 0.271818f
C78 source.n14 a_n1646_n1488# 0.250961f
C79 source.t10 a_n1646_n1488# 0.355982f
C80 source.n15 a_n1646_n1488# 0.378397f
C81 source.n16 a_n1646_n1488# 0.530926f
C82 drain_right.t7 a_n1646_n1488# 0.047274f
C83 drain_right.t3 a_n1646_n1488# 0.047274f
C84 drain_right.n0 a_n1646_n1488# 0.341985f
C85 drain_right.t2 a_n1646_n1488# 0.047274f
C86 drain_right.t1 a_n1646_n1488# 0.047274f
C87 drain_right.n1 a_n1646_n1488# 0.341985f
C88 drain_right.n2 a_n1646_n1488# 1.02178f
C89 drain_right.t5 a_n1646_n1488# 0.047274f
C90 drain_right.t6 a_n1646_n1488# 0.047274f
C91 drain_right.n3 a_n1646_n1488# 0.343633f
C92 drain_right.t0 a_n1646_n1488# 0.047274f
C93 drain_right.t4 a_n1646_n1488# 0.047274f
C94 drain_right.n4 a_n1646_n1488# 0.34094f
C95 drain_right.n5 a_n1646_n1488# 0.704532f
C96 minus.n0 a_n1646_n1488# 0.120705f
C97 minus.t4 a_n1646_n1488# 0.133612f
C98 minus.t6 a_n1646_n1488# 0.14358f
C99 minus.n1 a_n1646_n1488# 0.069788f
C100 minus.n2 a_n1646_n1488# 0.084631f
C101 minus.t3 a_n1646_n1488# 0.133612f
C102 minus.n3 a_n1646_n1488# 0.084631f
C103 minus.t2 a_n1646_n1488# 0.133612f
C104 minus.n4 a_n1646_n1488# 0.079014f
C105 minus.n5 a_n1646_n1488# 0.605815f
C106 minus.n6 a_n1646_n1488# 0.120705f
C107 minus.t7 a_n1646_n1488# 0.14358f
C108 minus.n7 a_n1646_n1488# 0.069788f
C109 minus.t1 a_n1646_n1488# 0.133612f
C110 minus.n8 a_n1646_n1488# 0.084631f
C111 minus.t0 a_n1646_n1488# 0.133612f
C112 minus.n9 a_n1646_n1488# 0.084631f
C113 minus.t5 a_n1646_n1488# 0.133612f
C114 minus.n10 a_n1646_n1488# 0.079014f
C115 minus.n11 a_n1646_n1488# 0.176735f
C116 minus.n12 a_n1646_n1488# 0.734821f
.ends

