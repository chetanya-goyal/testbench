* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t9 plus.t0 source.t19 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X1 source.t0 minus.t0 drain_right.t9 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X2 a_n1952_n1088# a_n1952_n1088# a_n1952_n1088# a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.7
X3 drain_left.t8 plus.t1 source.t11 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X4 drain_left.t7 plus.t2 source.t17 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X5 source.t9 minus.t1 drain_right.t8 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X6 drain_right.t7 minus.t2 source.t1 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X7 drain_right.t6 minus.t3 source.t6 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X8 source.t8 minus.t4 drain_right.t5 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X9 a_n1952_n1088# a_n1952_n1088# a_n1952_n1088# a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X10 drain_right.t4 minus.t5 source.t3 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X11 drain_right.t3 minus.t6 source.t5 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X12 source.t16 plus.t3 drain_left.t6 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X13 drain_right.t2 minus.t7 source.t7 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X14 drain_left.t5 plus.t4 source.t13 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X15 source.t18 plus.t5 drain_left.t4 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X16 a_n1952_n1088# a_n1952_n1088# a_n1952_n1088# a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X17 drain_right.t1 minus.t8 source.t2 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X18 source.t14 plus.t6 drain_left.t3 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X19 drain_left.t2 plus.t7 source.t15 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X20 a_n1952_n1088# a_n1952_n1088# a_n1952_n1088# a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X21 source.t4 minus.t9 drain_right.t0 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X22 source.t12 plus.t8 drain_left.t1 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X23 drain_left.t0 plus.t9 source.t10 a_n1952_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
R0 plus.n6 plus.n5 161.3
R1 plus.n7 plus.n2 161.3
R2 plus.n9 plus.n8 161.3
R3 plus.n10 plus.n1 161.3
R4 plus.n11 plus.n0 161.3
R5 plus.n13 plus.n12 161.3
R6 plus.n20 plus.n19 161.3
R7 plus.n21 plus.n16 161.3
R8 plus.n23 plus.n22 161.3
R9 plus.n24 plus.n15 161.3
R10 plus.n25 plus.n14 161.3
R11 plus.n27 plus.n26 161.3
R12 plus.n3 plus.t2 113.296
R13 plus.n17 plus.t4 113.296
R14 plus.n12 plus.t1 90.5476
R15 plus.n10 plus.t5 90.5476
R16 plus.n2 plus.t0 90.5476
R17 plus.n4 plus.t6 90.5476
R18 plus.n26 plus.t9 90.5476
R19 plus.n24 plus.t8 90.5476
R20 plus.n16 plus.t7 90.5476
R21 plus.n18 plus.t3 90.5476
R22 plus.n6 plus.n3 44.8741
R23 plus.n20 plus.n17 44.8741
R24 plus.n12 plus.n11 30.6732
R25 plus.n26 plus.n25 30.6732
R26 plus plus.n27 26.3683
R27 plus.n10 plus.n9 26.2914
R28 plus.n5 plus.n4 26.2914
R29 plus.n24 plus.n23 26.2914
R30 plus.n19 plus.n18 26.2914
R31 plus.n9 plus.n2 21.9096
R32 plus.n5 plus.n2 21.9096
R33 plus.n23 plus.n16 21.9096
R34 plus.n19 plus.n16 21.9096
R35 plus.n4 plus.n3 19.0667
R36 plus.n18 plus.n17 19.0667
R37 plus.n11 plus.n10 17.5278
R38 plus.n25 plus.n24 17.5278
R39 plus plus.n13 8.11603
R40 plus.n7 plus.n6 0.189894
R41 plus.n8 plus.n7 0.189894
R42 plus.n8 plus.n1 0.189894
R43 plus.n1 plus.n0 0.189894
R44 plus.n13 plus.n0 0.189894
R45 plus.n27 plus.n14 0.189894
R46 plus.n15 plus.n14 0.189894
R47 plus.n22 plus.n15 0.189894
R48 plus.n22 plus.n21 0.189894
R49 plus.n21 plus.n20 0.189894
R50 source.n0 source.t11 243.255
R51 source.n5 source.t2 243.255
R52 source.n19 source.t5 243.254
R53 source.n14 source.t13 243.254
R54 source.n2 source.n1 223.454
R55 source.n4 source.n3 223.454
R56 source.n7 source.n6 223.454
R57 source.n9 source.n8 223.454
R58 source.n18 source.n17 223.453
R59 source.n16 source.n15 223.453
R60 source.n13 source.n12 223.453
R61 source.n11 source.n10 223.453
R62 source.n17 source.t3 19.8005
R63 source.n17 source.t8 19.8005
R64 source.n15 source.t1 19.8005
R65 source.n15 source.t9 19.8005
R66 source.n12 source.t15 19.8005
R67 source.n12 source.t16 19.8005
R68 source.n10 source.t10 19.8005
R69 source.n10 source.t12 19.8005
R70 source.n1 source.t19 19.8005
R71 source.n1 source.t18 19.8005
R72 source.n3 source.t17 19.8005
R73 source.n3 source.t14 19.8005
R74 source.n6 source.t7 19.8005
R75 source.n6 source.t0 19.8005
R76 source.n8 source.t6 19.8005
R77 source.n8 source.t4 19.8005
R78 source.n11 source.n9 14.7303
R79 source.n20 source.n0 8.13543
R80 source.n20 source.n19 5.7074
R81 source.n5 source.n4 0.914293
R82 source.n16 source.n14 0.914293
R83 source.n9 source.n7 0.888431
R84 source.n7 source.n5 0.888431
R85 source.n4 source.n2 0.888431
R86 source.n2 source.n0 0.888431
R87 source.n13 source.n11 0.888431
R88 source.n14 source.n13 0.888431
R89 source.n18 source.n16 0.888431
R90 source.n19 source.n18 0.888431
R91 source source.n20 0.188
R92 drain_left.n5 drain_left.t7 260.82
R93 drain_left.n1 drain_left.t0 260.82
R94 drain_left.n3 drain_left.n2 240.743
R95 drain_left.n7 drain_left.n6 240.132
R96 drain_left.n5 drain_left.n4 240.132
R97 drain_left.n1 drain_left.n0 240.131
R98 drain_left drain_left.n3 22.8074
R99 drain_left.n2 drain_left.t6 19.8005
R100 drain_left.n2 drain_left.t5 19.8005
R101 drain_left.n0 drain_left.t1 19.8005
R102 drain_left.n0 drain_left.t2 19.8005
R103 drain_left.n6 drain_left.t4 19.8005
R104 drain_left.n6 drain_left.t8 19.8005
R105 drain_left.n4 drain_left.t3 19.8005
R106 drain_left.n4 drain_left.t9 19.8005
R107 drain_left drain_left.n7 6.54115
R108 drain_left.n7 drain_left.n5 0.888431
R109 drain_left.n3 drain_left.n1 0.167137
R110 minus.n13 minus.n12 161.3
R111 minus.n11 minus.n0 161.3
R112 minus.n10 minus.n9 161.3
R113 minus.n8 minus.n1 161.3
R114 minus.n7 minus.n6 161.3
R115 minus.n5 minus.n2 161.3
R116 minus.n27 minus.n26 161.3
R117 minus.n25 minus.n14 161.3
R118 minus.n24 minus.n23 161.3
R119 minus.n22 minus.n15 161.3
R120 minus.n21 minus.n20 161.3
R121 minus.n19 minus.n16 161.3
R122 minus.n3 minus.t8 113.296
R123 minus.n17 minus.t2 113.296
R124 minus.n4 minus.t0 90.5476
R125 minus.n6 minus.t7 90.5476
R126 minus.n10 minus.t9 90.5476
R127 minus.n12 minus.t3 90.5476
R128 minus.n18 minus.t1 90.5476
R129 minus.n20 minus.t5 90.5476
R130 minus.n24 minus.t4 90.5476
R131 minus.n26 minus.t6 90.5476
R132 minus.n3 minus.n2 44.8741
R133 minus.n17 minus.n16 44.8741
R134 minus.n12 minus.n11 30.6732
R135 minus.n26 minus.n25 30.6732
R136 minus.n28 minus.n13 28.3206
R137 minus.n5 minus.n4 26.2914
R138 minus.n10 minus.n1 26.2914
R139 minus.n19 minus.n18 26.2914
R140 minus.n24 minus.n15 26.2914
R141 minus.n6 minus.n5 21.9096
R142 minus.n6 minus.n1 21.9096
R143 minus.n20 minus.n19 21.9096
R144 minus.n20 minus.n15 21.9096
R145 minus.n4 minus.n3 19.0667
R146 minus.n18 minus.n17 19.0667
R147 minus.n11 minus.n10 17.5278
R148 minus.n25 minus.n24 17.5278
R149 minus.n28 minus.n27 6.63876
R150 minus.n13 minus.n0 0.189894
R151 minus.n9 minus.n0 0.189894
R152 minus.n9 minus.n8 0.189894
R153 minus.n8 minus.n7 0.189894
R154 minus.n7 minus.n2 0.189894
R155 minus.n21 minus.n16 0.189894
R156 minus.n22 minus.n21 0.189894
R157 minus.n23 minus.n22 0.189894
R158 minus.n23 minus.n14 0.189894
R159 minus.n27 minus.n14 0.189894
R160 minus minus.n28 0.188
R161 drain_right.n1 drain_right.t7 260.82
R162 drain_right.n7 drain_right.t6 259.933
R163 drain_right.n6 drain_right.n4 241.02
R164 drain_right.n3 drain_right.n2 240.743
R165 drain_right.n6 drain_right.n5 240.132
R166 drain_right.n1 drain_right.n0 240.131
R167 drain_right drain_right.n3 22.2542
R168 drain_right.n2 drain_right.t5 19.8005
R169 drain_right.n2 drain_right.t3 19.8005
R170 drain_right.n0 drain_right.t8 19.8005
R171 drain_right.n0 drain_right.t4 19.8005
R172 drain_right.n4 drain_right.t9 19.8005
R173 drain_right.n4 drain_right.t1 19.8005
R174 drain_right.n5 drain_right.t0 19.8005
R175 drain_right.n5 drain_right.t2 19.8005
R176 drain_right drain_right.n7 6.09718
R177 drain_right.n7 drain_right.n6 0.888431
R178 drain_right.n3 drain_right.n1 0.167137
C0 source drain_right 3.55073f
C1 drain_right plus 0.354549f
C2 drain_right drain_left 0.965706f
C3 source minus 1.41895f
C4 minus plus 3.54935f
C5 drain_left minus 0.179761f
C6 source plus 1.43286f
C7 source drain_left 3.5503f
C8 drain_left plus 1.15792f
C9 drain_right minus 0.967941f
C10 drain_right a_n1952_n1088# 3.566106f
C11 drain_left a_n1952_n1088# 3.82321f
C12 source a_n1952_n1088# 2.189102f
C13 minus a_n1952_n1088# 6.715978f
C14 plus a_n1952_n1088# 7.319394f
C15 drain_right.t7 a_n1952_n1088# 0.096269f
C16 drain_right.t8 a_n1952_n1088# 0.01545f
C17 drain_right.t4 a_n1952_n1088# 0.01545f
C18 drain_right.n0 a_n1952_n1088# 0.060033f
C19 drain_right.n1 a_n1952_n1088# 0.412313f
C20 drain_right.t5 a_n1952_n1088# 0.01545f
C21 drain_right.t3 a_n1952_n1088# 0.01545f
C22 drain_right.n2 a_n1952_n1088# 0.060641f
C23 drain_right.n3 a_n1952_n1088# 0.764795f
C24 drain_right.t9 a_n1952_n1088# 0.01545f
C25 drain_right.t1 a_n1952_n1088# 0.01545f
C26 drain_right.n4 a_n1952_n1088# 0.060978f
C27 drain_right.t0 a_n1952_n1088# 0.01545f
C28 drain_right.t2 a_n1952_n1088# 0.01545f
C29 drain_right.n5 a_n1952_n1088# 0.060033f
C30 drain_right.n6 a_n1952_n1088# 0.504125f
C31 drain_right.t6 a_n1952_n1088# 0.095564f
C32 drain_right.n7 a_n1952_n1088# 0.386825f
C33 minus.n0 a_n1952_n1088# 0.027864f
C34 minus.n1 a_n1952_n1088# 0.006323f
C35 minus.t9 a_n1952_n1088# 0.066141f
C36 minus.n2 a_n1952_n1088# 0.116383f
C37 minus.t8 a_n1952_n1088# 0.079324f
C38 minus.n3 a_n1952_n1088# 0.055111f
C39 minus.t0 a_n1952_n1088# 0.066141f
C40 minus.n4 a_n1952_n1088# 0.068561f
C41 minus.n5 a_n1952_n1088# 0.006323f
C42 minus.t7 a_n1952_n1088# 0.066141f
C43 minus.n6 a_n1952_n1088# 0.065753f
C44 minus.n7 a_n1952_n1088# 0.027864f
C45 minus.n8 a_n1952_n1088# 0.027864f
C46 minus.n9 a_n1952_n1088# 0.027864f
C47 minus.n10 a_n1952_n1088# 0.065753f
C48 minus.n11 a_n1952_n1088# 0.006323f
C49 minus.t3 a_n1952_n1088# 0.066141f
C50 minus.n12 a_n1952_n1088# 0.064207f
C51 minus.n13 a_n1952_n1088# 0.659794f
C52 minus.n14 a_n1952_n1088# 0.027864f
C53 minus.n15 a_n1952_n1088# 0.006323f
C54 minus.n16 a_n1952_n1088# 0.116383f
C55 minus.t2 a_n1952_n1088# 0.079324f
C56 minus.n17 a_n1952_n1088# 0.055111f
C57 minus.t1 a_n1952_n1088# 0.066141f
C58 minus.n18 a_n1952_n1088# 0.068561f
C59 minus.n19 a_n1952_n1088# 0.006323f
C60 minus.t5 a_n1952_n1088# 0.066141f
C61 minus.n20 a_n1952_n1088# 0.065753f
C62 minus.n21 a_n1952_n1088# 0.027864f
C63 minus.n22 a_n1952_n1088# 0.027864f
C64 minus.n23 a_n1952_n1088# 0.027864f
C65 minus.t4 a_n1952_n1088# 0.066141f
C66 minus.n24 a_n1952_n1088# 0.065753f
C67 minus.n25 a_n1952_n1088# 0.006323f
C68 minus.t6 a_n1952_n1088# 0.066141f
C69 minus.n26 a_n1952_n1088# 0.064207f
C70 minus.n27 a_n1952_n1088# 0.191219f
C71 minus.n28 a_n1952_n1088# 0.810523f
C72 drain_left.t0 a_n1952_n1088# 0.094266f
C73 drain_left.t1 a_n1952_n1088# 0.015128f
C74 drain_left.t2 a_n1952_n1088# 0.015128f
C75 drain_left.n0 a_n1952_n1088# 0.058784f
C76 drain_left.n1 a_n1952_n1088# 0.403735f
C77 drain_left.t6 a_n1952_n1088# 0.015128f
C78 drain_left.t5 a_n1952_n1088# 0.015128f
C79 drain_left.n2 a_n1952_n1088# 0.05938f
C80 drain_left.n3 a_n1952_n1088# 0.785865f
C81 drain_left.t7 a_n1952_n1088# 0.094266f
C82 drain_left.t3 a_n1952_n1088# 0.015128f
C83 drain_left.t9 a_n1952_n1088# 0.015128f
C84 drain_left.n4 a_n1952_n1088# 0.058784f
C85 drain_left.n5 a_n1952_n1088# 0.445566f
C86 drain_left.t4 a_n1952_n1088# 0.015128f
C87 drain_left.t8 a_n1952_n1088# 0.015128f
C88 drain_left.n6 a_n1952_n1088# 0.058784f
C89 drain_left.n7 a_n1952_n1088# 0.412758f
C90 source.t11 a_n1952_n1088# 0.117035f
C91 source.n0 a_n1952_n1088# 0.555327f
C92 source.t19 a_n1952_n1088# 0.021027f
C93 source.t18 a_n1952_n1088# 0.021027f
C94 source.n1 a_n1952_n1088# 0.068195f
C95 source.n2 a_n1952_n1088# 0.315687f
C96 source.t17 a_n1952_n1088# 0.021027f
C97 source.t14 a_n1952_n1088# 0.021027f
C98 source.n3 a_n1952_n1088# 0.068195f
C99 source.n4 a_n1952_n1088# 0.317904f
C100 source.t2 a_n1952_n1088# 0.117035f
C101 source.n5 a_n1952_n1088# 0.326412f
C102 source.t7 a_n1952_n1088# 0.021027f
C103 source.t0 a_n1952_n1088# 0.021027f
C104 source.n6 a_n1952_n1088# 0.068195f
C105 source.n7 a_n1952_n1088# 0.315687f
C106 source.t6 a_n1952_n1088# 0.021027f
C107 source.t4 a_n1952_n1088# 0.021027f
C108 source.n8 a_n1952_n1088# 0.068195f
C109 source.n9 a_n1952_n1088# 0.842503f
C110 source.t10 a_n1952_n1088# 0.021027f
C111 source.t12 a_n1952_n1088# 0.021027f
C112 source.n10 a_n1952_n1088# 0.068195f
C113 source.n11 a_n1952_n1088# 0.842504f
C114 source.t15 a_n1952_n1088# 0.021027f
C115 source.t16 a_n1952_n1088# 0.021027f
C116 source.n12 a_n1952_n1088# 0.068195f
C117 source.n13 a_n1952_n1088# 0.315687f
C118 source.t13 a_n1952_n1088# 0.117035f
C119 source.n14 a_n1952_n1088# 0.326412f
C120 source.t1 a_n1952_n1088# 0.021027f
C121 source.t9 a_n1952_n1088# 0.021027f
C122 source.n15 a_n1952_n1088# 0.068195f
C123 source.n16 a_n1952_n1088# 0.317905f
C124 source.t3 a_n1952_n1088# 0.021027f
C125 source.t8 a_n1952_n1088# 0.021027f
C126 source.n17 a_n1952_n1088# 0.068195f
C127 source.n18 a_n1952_n1088# 0.315687f
C128 source.t5 a_n1952_n1088# 0.117035f
C129 source.n19 a_n1952_n1088# 0.461918f
C130 source.n20 a_n1952_n1088# 0.55144f
C131 plus.n0 a_n1952_n1088# 0.02832f
C132 plus.t1 a_n1952_n1088# 0.067223f
C133 plus.t5 a_n1952_n1088# 0.067223f
C134 plus.n1 a_n1952_n1088# 0.02832f
C135 plus.t0 a_n1952_n1088# 0.067223f
C136 plus.n2 a_n1952_n1088# 0.066829f
C137 plus.t2 a_n1952_n1088# 0.080622f
C138 plus.n3 a_n1952_n1088# 0.056013f
C139 plus.t6 a_n1952_n1088# 0.067223f
C140 plus.n4 a_n1952_n1088# 0.069683f
C141 plus.n5 a_n1952_n1088# 0.006426f
C142 plus.n6 a_n1952_n1088# 0.118287f
C143 plus.n7 a_n1952_n1088# 0.02832f
C144 plus.n8 a_n1952_n1088# 0.02832f
C145 plus.n9 a_n1952_n1088# 0.006426f
C146 plus.n10 a_n1952_n1088# 0.066829f
C147 plus.n11 a_n1952_n1088# 0.006426f
C148 plus.n12 a_n1952_n1088# 0.065258f
C149 plus.n13 a_n1952_n1088# 0.203861f
C150 plus.n14 a_n1952_n1088# 0.02832f
C151 plus.t9 a_n1952_n1088# 0.067223f
C152 plus.n15 a_n1952_n1088# 0.02832f
C153 plus.t8 a_n1952_n1088# 0.067223f
C154 plus.t7 a_n1952_n1088# 0.067223f
C155 plus.n16 a_n1952_n1088# 0.066829f
C156 plus.t4 a_n1952_n1088# 0.080622f
C157 plus.n17 a_n1952_n1088# 0.056013f
C158 plus.t3 a_n1952_n1088# 0.067223f
C159 plus.n18 a_n1952_n1088# 0.069683f
C160 plus.n19 a_n1952_n1088# 0.006426f
C161 plus.n20 a_n1952_n1088# 0.118287f
C162 plus.n21 a_n1952_n1088# 0.02832f
C163 plus.n22 a_n1952_n1088# 0.02832f
C164 plus.n23 a_n1952_n1088# 0.006426f
C165 plus.n24 a_n1952_n1088# 0.066829f
C166 plus.n25 a_n1952_n1088# 0.006426f
C167 plus.n26 a_n1952_n1088# 0.065258f
C168 plus.n27 a_n1952_n1088# 0.649786f
.ends

