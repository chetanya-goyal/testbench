* NGSPICE file created from diffpair421.ext - technology: sky130A

.subckt diffpair421 minus drain_right drain_left source plus
X0 drain_right minus source a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X1 a_n1064_n3292# a_n1064_n3292# a_n1064_n3292# a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.25
X2 source plus drain_left a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X3 drain_left plus source a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X4 source minus drain_right a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X5 a_n1064_n3292# a_n1064_n3292# a_n1064_n3292# a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X6 drain_left plus source a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X7 source minus drain_right a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X8 a_n1064_n3292# a_n1064_n3292# a_n1064_n3292# a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X9 drain_right minus source a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X10 source plus drain_left a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X11 a_n1064_n3292# a_n1064_n3292# a_n1064_n3292# a_n1064_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
.ends

