* NGSPICE file created from diffpair566.ext - technology: sky130A

.subckt diffpair566 minus drain_right drain_left source plus
X0 drain_right.t13 minus.t0 source.t19 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X1 source.t22 minus.t1 drain_right.t12 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X2 drain_right.t11 minus.t2 source.t25 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X3 source.t3 plus.t0 drain_left.t13 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X4 a_n1756_n4888# a_n1756_n4888# a_n1756_n4888# a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=76 ps=327.6 w=20 l=0.15
X5 a_n1756_n4888# a_n1756_n4888# a_n1756_n4888# a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X6 drain_left.t12 plus.t1 source.t8 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X7 a_n1756_n4888# a_n1756_n4888# a_n1756_n4888# a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X8 drain_left.t11 plus.t2 source.t12 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X9 a_n1756_n4888# a_n1756_n4888# a_n1756_n4888# a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X10 source.t14 minus.t3 drain_right.t10 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X11 source.t2 plus.t3 drain_left.t10 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X12 drain_right.t9 minus.t4 source.t17 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X13 drain_right.t8 minus.t5 source.t20 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X14 drain_right.t7 minus.t6 source.t24 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X15 source.t18 minus.t7 drain_right.t6 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X16 drain_left.t9 plus.t4 source.t11 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X17 drain_left.t8 plus.t5 source.t4 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X18 drain_right.t5 minus.t8 source.t26 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X19 drain_right.t4 minus.t9 source.t16 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X20 source.t23 minus.t10 drain_right.t3 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X21 drain_left.t7 plus.t6 source.t13 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X22 source.t1 plus.t7 drain_left.t6 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X23 source.t27 minus.t11 drain_right.t2 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X24 source.t15 minus.t12 drain_right.t1 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X25 drain_left.t5 plus.t8 source.t7 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X26 drain_left.t4 plus.t9 source.t10 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X27 source.t5 plus.t10 drain_left.t3 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X28 source.t6 plus.t11 drain_left.t2 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X29 source.t9 plus.t12 drain_left.t1 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X30 drain_right.t0 minus.t13 source.t21 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X31 drain_left.t0 plus.t13 source.t0 a_n1756_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
R0 minus.n15 minus.t9 3487.93
R1 minus.n3 minus.t4 3487.93
R2 minus.n32 minus.t0 3487.93
R3 minus.n20 minus.t2 3487.93
R4 minus.n1 minus.t7 3422.2
R5 minus.n14 minus.t11 3422.2
R6 minus.n12 minus.t5 3422.2
R7 minus.n6 minus.t8 3422.2
R8 minus.n4 minus.t3 3422.2
R9 minus.n18 minus.t1 3422.2
R10 minus.n31 minus.t12 3422.2
R11 minus.n29 minus.t6 3422.2
R12 minus.n23 minus.t13 3422.2
R13 minus.n21 minus.t10 3422.2
R14 minus.n3 minus.n2 161.489
R15 minus.n20 minus.n19 161.489
R16 minus.n16 minus.n15 161.3
R17 minus.n13 minus.n0 161.3
R18 minus.n11 minus.n10 161.3
R19 minus.n9 minus.n1 161.3
R20 minus.n8 minus.n7 161.3
R21 minus.n5 minus.n2 161.3
R22 minus.n33 minus.n32 161.3
R23 minus.n30 minus.n17 161.3
R24 minus.n28 minus.n27 161.3
R25 minus.n26 minus.n18 161.3
R26 minus.n25 minus.n24 161.3
R27 minus.n22 minus.n19 161.3
R28 minus.n11 minus.n1 73.0308
R29 minus.n7 minus.n1 73.0308
R30 minus.n24 minus.n18 73.0308
R31 minus.n28 minus.n18 73.0308
R32 minus.n13 minus.n12 51.1217
R33 minus.n6 minus.n5 51.1217
R34 minus.n23 minus.n22 51.1217
R35 minus.n30 minus.n29 51.1217
R36 minus.n14 minus.n13 43.8187
R37 minus.n5 minus.n4 43.8187
R38 minus.n22 minus.n21 43.8187
R39 minus.n31 minus.n30 43.8187
R40 minus.n34 minus.n16 41.9039
R41 minus.n15 minus.n14 29.2126
R42 minus.n4 minus.n3 29.2126
R43 minus.n21 minus.n20 29.2126
R44 minus.n32 minus.n31 29.2126
R45 minus.n12 minus.n11 21.9096
R46 minus.n7 minus.n6 21.9096
R47 minus.n24 minus.n23 21.9096
R48 minus.n29 minus.n28 21.9096
R49 minus.n34 minus.n33 6.57058
R50 minus.n16 minus.n0 0.189894
R51 minus.n10 minus.n0 0.189894
R52 minus.n10 minus.n9 0.189894
R53 minus.n9 minus.n8 0.189894
R54 minus.n8 minus.n2 0.189894
R55 minus.n25 minus.n19 0.189894
R56 minus.n26 minus.n25 0.189894
R57 minus.n27 minus.n26 0.189894
R58 minus.n27 minus.n17 0.189894
R59 minus.n33 minus.n17 0.189894
R60 minus minus.n34 0.188
R61 source.n0 source.t7 44.6397
R62 source.n7 source.t17 44.6396
R63 source.n27 source.t19 44.6395
R64 source.n20 source.t11 44.6395
R65 source.n2 source.n1 43.1397
R66 source.n4 source.n3 43.1397
R67 source.n6 source.n5 43.1397
R68 source.n9 source.n8 43.1397
R69 source.n11 source.n10 43.1397
R70 source.n13 source.n12 43.1397
R71 source.n26 source.n25 43.1396
R72 source.n24 source.n23 43.1396
R73 source.n22 source.n21 43.1396
R74 source.n19 source.n18 43.1396
R75 source.n17 source.n16 43.1396
R76 source.n15 source.n14 43.1396
R77 source.n15 source.n13 28.469
R78 source.n28 source.n0 22.3656
R79 source.n28 source.n27 5.5436
R80 source.n25 source.t24 1.5005
R81 source.n25 source.t15 1.5005
R82 source.n23 source.t21 1.5005
R83 source.n23 source.t22 1.5005
R84 source.n21 source.t25 1.5005
R85 source.n21 source.t23 1.5005
R86 source.n18 source.t8 1.5005
R87 source.n18 source.t5 1.5005
R88 source.n16 source.t13 1.5005
R89 source.n16 source.t2 1.5005
R90 source.n14 source.t12 1.5005
R91 source.n14 source.t3 1.5005
R92 source.n1 source.t0 1.5005
R93 source.n1 source.t6 1.5005
R94 source.n3 source.t10 1.5005
R95 source.n3 source.t1 1.5005
R96 source.n5 source.t4 1.5005
R97 source.n5 source.t9 1.5005
R98 source.n8 source.t26 1.5005
R99 source.n8 source.t14 1.5005
R100 source.n10 source.t20 1.5005
R101 source.n10 source.t18 1.5005
R102 source.n12 source.t16 1.5005
R103 source.n12 source.t27 1.5005
R104 source.n7 source.n6 0.7505
R105 source.n22 source.n20 0.7505
R106 source.n13 source.n11 0.560845
R107 source.n11 source.n9 0.560845
R108 source.n9 source.n7 0.560845
R109 source.n6 source.n4 0.560845
R110 source.n4 source.n2 0.560845
R111 source.n2 source.n0 0.560845
R112 source.n17 source.n15 0.560845
R113 source.n19 source.n17 0.560845
R114 source.n20 source.n19 0.560845
R115 source.n24 source.n22 0.560845
R116 source.n26 source.n24 0.560845
R117 source.n27 source.n26 0.560845
R118 source source.n28 0.188
R119 drain_right.n1 drain_right.t11 61.8786
R120 drain_right.n11 drain_right.t4 61.3184
R121 drain_right.n8 drain_right.n6 60.3788
R122 drain_right.n4 drain_right.n2 60.3788
R123 drain_right.n8 drain_right.n7 59.8185
R124 drain_right.n10 drain_right.n9 59.8185
R125 drain_right.n4 drain_right.n3 59.8184
R126 drain_right.n1 drain_right.n0 59.8184
R127 drain_right drain_right.n5 36.0964
R128 drain_right drain_right.n11 5.93339
R129 drain_right.n2 drain_right.t1 1.5005
R130 drain_right.n2 drain_right.t13 1.5005
R131 drain_right.n3 drain_right.t12 1.5005
R132 drain_right.n3 drain_right.t7 1.5005
R133 drain_right.n0 drain_right.t3 1.5005
R134 drain_right.n0 drain_right.t0 1.5005
R135 drain_right.n6 drain_right.t10 1.5005
R136 drain_right.n6 drain_right.t9 1.5005
R137 drain_right.n7 drain_right.t6 1.5005
R138 drain_right.n7 drain_right.t5 1.5005
R139 drain_right.n9 drain_right.t2 1.5005
R140 drain_right.n9 drain_right.t8 1.5005
R141 drain_right.n11 drain_right.n10 0.560845
R142 drain_right.n10 drain_right.n8 0.560845
R143 drain_right.n5 drain_right.n1 0.365413
R144 drain_right.n5 drain_right.n4 0.0852402
R145 plus.n3 plus.t5 3487.93
R146 plus.n15 plus.t8 3487.93
R147 plus.n20 plus.t4 3487.93
R148 plus.n32 plus.t2 3487.93
R149 plus.n1 plus.t7 3422.2
R150 plus.n4 plus.t12 3422.2
R151 plus.n6 plus.t9 3422.2
R152 plus.n12 plus.t13 3422.2
R153 plus.n14 plus.t11 3422.2
R154 plus.n18 plus.t3 3422.2
R155 plus.n21 plus.t10 3422.2
R156 plus.n23 plus.t1 3422.2
R157 plus.n29 plus.t6 3422.2
R158 plus.n31 plus.t0 3422.2
R159 plus.n3 plus.n2 161.489
R160 plus.n20 plus.n19 161.489
R161 plus.n5 plus.n2 161.3
R162 plus.n8 plus.n7 161.3
R163 plus.n9 plus.n1 161.3
R164 plus.n11 plus.n10 161.3
R165 plus.n13 plus.n0 161.3
R166 plus.n16 plus.n15 161.3
R167 plus.n22 plus.n19 161.3
R168 plus.n25 plus.n24 161.3
R169 plus.n26 plus.n18 161.3
R170 plus.n28 plus.n27 161.3
R171 plus.n30 plus.n17 161.3
R172 plus.n33 plus.n32 161.3
R173 plus.n7 plus.n1 73.0308
R174 plus.n11 plus.n1 73.0308
R175 plus.n28 plus.n18 73.0308
R176 plus.n24 plus.n18 73.0308
R177 plus.n6 plus.n5 51.1217
R178 plus.n13 plus.n12 51.1217
R179 plus.n30 plus.n29 51.1217
R180 plus.n23 plus.n22 51.1217
R181 plus.n5 plus.n4 43.8187
R182 plus.n14 plus.n13 43.8187
R183 plus.n31 plus.n30 43.8187
R184 plus.n22 plus.n21 43.8187
R185 plus plus.n33 32.7547
R186 plus.n4 plus.n3 29.2126
R187 plus.n15 plus.n14 29.2126
R188 plus.n32 plus.n31 29.2126
R189 plus.n21 plus.n20 29.2126
R190 plus.n7 plus.n6 21.9096
R191 plus.n12 plus.n11 21.9096
R192 plus.n29 plus.n28 21.9096
R193 plus.n24 plus.n23 21.9096
R194 plus plus.n16 15.2448
R195 plus.n8 plus.n2 0.189894
R196 plus.n9 plus.n8 0.189894
R197 plus.n10 plus.n9 0.189894
R198 plus.n10 plus.n0 0.189894
R199 plus.n16 plus.n0 0.189894
R200 plus.n33 plus.n17 0.189894
R201 plus.n27 plus.n17 0.189894
R202 plus.n27 plus.n26 0.189894
R203 plus.n26 plus.n25 0.189894
R204 plus.n25 plus.n19 0.189894
R205 drain_left.n7 drain_left.t8 61.8788
R206 drain_left.n1 drain_left.t11 61.8786
R207 drain_left.n4 drain_left.n2 60.3788
R208 drain_left.n11 drain_left.n10 59.8185
R209 drain_left.n9 drain_left.n8 59.8185
R210 drain_left.n7 drain_left.n6 59.8185
R211 drain_left.n4 drain_left.n3 59.8184
R212 drain_left.n1 drain_left.n0 59.8184
R213 drain_left drain_left.n5 36.6497
R214 drain_left drain_left.n11 6.21356
R215 drain_left.n2 drain_left.t3 1.5005
R216 drain_left.n2 drain_left.t9 1.5005
R217 drain_left.n3 drain_left.t10 1.5005
R218 drain_left.n3 drain_left.t12 1.5005
R219 drain_left.n0 drain_left.t13 1.5005
R220 drain_left.n0 drain_left.t7 1.5005
R221 drain_left.n10 drain_left.t2 1.5005
R222 drain_left.n10 drain_left.t5 1.5005
R223 drain_left.n8 drain_left.t6 1.5005
R224 drain_left.n8 drain_left.t0 1.5005
R225 drain_left.n6 drain_left.t1 1.5005
R226 drain_left.n6 drain_left.t4 1.5005
R227 drain_left.n9 drain_left.n7 0.560845
R228 drain_left.n11 drain_left.n9 0.560845
R229 drain_left.n5 drain_left.n1 0.365413
R230 drain_left.n5 drain_left.n4 0.0852402
C0 source minus 4.12923f
C1 drain_left minus 0.171187f
C2 source drain_left 45.833103f
C3 drain_right plus 0.327552f
C4 plus minus 6.80545f
C5 source plus 4.14434f
C6 drain_left plus 5.1773f
C7 drain_right minus 5.01189f
C8 source drain_right 45.8165f
C9 drain_left drain_right 0.904571f
C10 drain_right a_n1756_n4888# 9.20186f
C11 drain_left a_n1756_n4888# 9.47571f
C12 source a_n1756_n4888# 9.031098f
C13 minus a_n1756_n4888# 6.999496f
C14 plus a_n1756_n4888# 9.74832f
C15 drain_left.t11 a_n1756_n4888# 5.20335f
C16 drain_left.t13 a_n1756_n4888# 0.624223f
C17 drain_left.t7 a_n1756_n4888# 0.624223f
C18 drain_left.n0 a_n1756_n4888# 4.19095f
C19 drain_left.n1 a_n1756_n4888# 0.688087f
C20 drain_left.t3 a_n1756_n4888# 0.624223f
C21 drain_left.t9 a_n1756_n4888# 0.624223f
C22 drain_left.n2 a_n1756_n4888# 4.19396f
C23 drain_left.t10 a_n1756_n4888# 0.624223f
C24 drain_left.t12 a_n1756_n4888# 0.624223f
C25 drain_left.n3 a_n1756_n4888# 4.19095f
C26 drain_left.n4 a_n1756_n4888# 0.602881f
C27 drain_left.n5 a_n1756_n4888# 1.76243f
C28 drain_left.t8 a_n1756_n4888# 5.20337f
C29 drain_left.t1 a_n1756_n4888# 0.624223f
C30 drain_left.t4 a_n1756_n4888# 0.624223f
C31 drain_left.n6 a_n1756_n4888# 4.19095f
C32 drain_left.n7 a_n1756_n4888# 0.702833f
C33 drain_left.t6 a_n1756_n4888# 0.624223f
C34 drain_left.t0 a_n1756_n4888# 0.624223f
C35 drain_left.n8 a_n1756_n4888# 4.19095f
C36 drain_left.n9 a_n1756_n4888# 0.314111f
C37 drain_left.t2 a_n1756_n4888# 0.624223f
C38 drain_left.t5 a_n1756_n4888# 0.624223f
C39 drain_left.n10 a_n1756_n4888# 4.19095f
C40 drain_left.n11 a_n1756_n4888# 0.531803f
C41 plus.n0 a_n1756_n4888# 0.056425f
C42 plus.t11 a_n1756_n4888# 0.476763f
C43 plus.t13 a_n1756_n4888# 0.476763f
C44 plus.t7 a_n1756_n4888# 0.476763f
C45 plus.n1 a_n1756_n4888# 0.204521f
C46 plus.n2 a_n1756_n4888# 0.131896f
C47 plus.t9 a_n1756_n4888# 0.476763f
C48 plus.t12 a_n1756_n4888# 0.476763f
C49 plus.t5 a_n1756_n4888# 0.48033f
C50 plus.n3 a_n1756_n4888# 0.20974f
C51 plus.n4 a_n1756_n4888# 0.185803f
C52 plus.n5 a_n1756_n4888# 0.023937f
C53 plus.n6 a_n1756_n4888# 0.185803f
C54 plus.n7 a_n1756_n4888# 0.023937f
C55 plus.n8 a_n1756_n4888# 0.056425f
C56 plus.n9 a_n1756_n4888# 0.056425f
C57 plus.n10 a_n1756_n4888# 0.056425f
C58 plus.n11 a_n1756_n4888# 0.023937f
C59 plus.n12 a_n1756_n4888# 0.185803f
C60 plus.n13 a_n1756_n4888# 0.023937f
C61 plus.n14 a_n1756_n4888# 0.185803f
C62 plus.t8 a_n1756_n4888# 0.48033f
C63 plus.n15 a_n1756_n4888# 0.209652f
C64 plus.n16 a_n1756_n4888# 0.865929f
C65 plus.n17 a_n1756_n4888# 0.056425f
C66 plus.t2 a_n1756_n4888# 0.48033f
C67 plus.t0 a_n1756_n4888# 0.476763f
C68 plus.t6 a_n1756_n4888# 0.476763f
C69 plus.t3 a_n1756_n4888# 0.476763f
C70 plus.n18 a_n1756_n4888# 0.204521f
C71 plus.n19 a_n1756_n4888# 0.131896f
C72 plus.t1 a_n1756_n4888# 0.476763f
C73 plus.t10 a_n1756_n4888# 0.476763f
C74 plus.t4 a_n1756_n4888# 0.48033f
C75 plus.n20 a_n1756_n4888# 0.20974f
C76 plus.n21 a_n1756_n4888# 0.185803f
C77 plus.n22 a_n1756_n4888# 0.023937f
C78 plus.n23 a_n1756_n4888# 0.185803f
C79 plus.n24 a_n1756_n4888# 0.023937f
C80 plus.n25 a_n1756_n4888# 0.056425f
C81 plus.n26 a_n1756_n4888# 0.056425f
C82 plus.n27 a_n1756_n4888# 0.056425f
C83 plus.n28 a_n1756_n4888# 0.023937f
C84 plus.n29 a_n1756_n4888# 0.185803f
C85 plus.n30 a_n1756_n4888# 0.023937f
C86 plus.n31 a_n1756_n4888# 0.185803f
C87 plus.n32 a_n1756_n4888# 0.209652f
C88 plus.n33 a_n1756_n4888# 1.97119f
C89 drain_right.t11 a_n1756_n4888# 5.19333f
C90 drain_right.t3 a_n1756_n4888# 0.623021f
C91 drain_right.t0 a_n1756_n4888# 0.623021f
C92 drain_right.n0 a_n1756_n4888# 4.18288f
C93 drain_right.n1 a_n1756_n4888# 0.686761f
C94 drain_right.t1 a_n1756_n4888# 0.623021f
C95 drain_right.t13 a_n1756_n4888# 0.623021f
C96 drain_right.n2 a_n1756_n4888# 4.18589f
C97 drain_right.t12 a_n1756_n4888# 0.623021f
C98 drain_right.t7 a_n1756_n4888# 0.623021f
C99 drain_right.n3 a_n1756_n4888# 4.18288f
C100 drain_right.n4 a_n1756_n4888# 0.60172f
C101 drain_right.n5 a_n1756_n4888# 1.70482f
C102 drain_right.t10 a_n1756_n4888# 0.623021f
C103 drain_right.t9 a_n1756_n4888# 0.623021f
C104 drain_right.n6 a_n1756_n4888# 4.18588f
C105 drain_right.t6 a_n1756_n4888# 0.623021f
C106 drain_right.t5 a_n1756_n4888# 0.623021f
C107 drain_right.n7 a_n1756_n4888# 4.18287f
C108 drain_right.n8 a_n1756_n4888# 0.634484f
C109 drain_right.t2 a_n1756_n4888# 0.623021f
C110 drain_right.t8 a_n1756_n4888# 0.623021f
C111 drain_right.n9 a_n1756_n4888# 4.18287f
C112 drain_right.n10 a_n1756_n4888# 0.313506f
C113 drain_right.t4 a_n1756_n4888# 5.1898f
C114 drain_right.n11 a_n1756_n4888# 0.609682f
C115 source.t7 a_n1756_n4888# 5.10534f
C116 source.n0 a_n1756_n4888# 2.07279f
C117 source.t0 a_n1756_n4888# 0.627756f
C118 source.t6 a_n1756_n4888# 0.627756f
C119 source.n1 a_n1756_n4888# 4.13106f
C120 source.n2 a_n1756_n4888# 0.363858f
C121 source.t10 a_n1756_n4888# 0.627756f
C122 source.t1 a_n1756_n4888# 0.627756f
C123 source.n3 a_n1756_n4888# 4.13106f
C124 source.n4 a_n1756_n4888# 0.363858f
C125 source.t4 a_n1756_n4888# 0.627756f
C126 source.t9 a_n1756_n4888# 0.627756f
C127 source.n5 a_n1756_n4888# 4.13106f
C128 source.n6 a_n1756_n4888# 0.379879f
C129 source.t17 a_n1756_n4888# 5.10535f
C130 source.n7 a_n1756_n4888# 0.53556f
C131 source.t26 a_n1756_n4888# 0.627756f
C132 source.t14 a_n1756_n4888# 0.627756f
C133 source.n8 a_n1756_n4888# 4.13106f
C134 source.n9 a_n1756_n4888# 0.363858f
C135 source.t20 a_n1756_n4888# 0.627756f
C136 source.t18 a_n1756_n4888# 0.627756f
C137 source.n10 a_n1756_n4888# 4.13106f
C138 source.n11 a_n1756_n4888# 0.363858f
C139 source.t16 a_n1756_n4888# 0.627756f
C140 source.t27 a_n1756_n4888# 0.627756f
C141 source.n12 a_n1756_n4888# 4.13106f
C142 source.n13 a_n1756_n4888# 2.42962f
C143 source.t12 a_n1756_n4888# 0.627756f
C144 source.t3 a_n1756_n4888# 0.627756f
C145 source.n14 a_n1756_n4888# 4.13107f
C146 source.n15 a_n1756_n4888# 2.42961f
C147 source.t13 a_n1756_n4888# 0.627756f
C148 source.t2 a_n1756_n4888# 0.627756f
C149 source.n16 a_n1756_n4888# 4.13107f
C150 source.n17 a_n1756_n4888# 0.363851f
C151 source.t8 a_n1756_n4888# 0.627756f
C152 source.t5 a_n1756_n4888# 0.627756f
C153 source.n18 a_n1756_n4888# 4.13107f
C154 source.n19 a_n1756_n4888# 0.363851f
C155 source.t11 a_n1756_n4888# 5.10532f
C156 source.n20 a_n1756_n4888# 0.535586f
C157 source.t25 a_n1756_n4888# 0.627756f
C158 source.t23 a_n1756_n4888# 0.627756f
C159 source.n21 a_n1756_n4888# 4.13107f
C160 source.n22 a_n1756_n4888# 0.379872f
C161 source.t21 a_n1756_n4888# 0.627756f
C162 source.t22 a_n1756_n4888# 0.627756f
C163 source.n23 a_n1756_n4888# 4.13107f
C164 source.n24 a_n1756_n4888# 0.363851f
C165 source.t24 a_n1756_n4888# 0.627756f
C166 source.t15 a_n1756_n4888# 0.627756f
C167 source.n25 a_n1756_n4888# 4.13107f
C168 source.n26 a_n1756_n4888# 0.363851f
C169 source.t19 a_n1756_n4888# 5.10532f
C170 source.n27 a_n1756_n4888# 0.661067f
C171 source.n28 a_n1756_n4888# 2.36076f
C172 minus.n0 a_n1756_n4888# 0.055332f
C173 minus.t9 a_n1756_n4888# 0.471025f
C174 minus.t11 a_n1756_n4888# 0.467527f
C175 minus.t5 a_n1756_n4888# 0.467527f
C176 minus.t7 a_n1756_n4888# 0.467527f
C177 minus.n1 a_n1756_n4888# 0.200559f
C178 minus.n2 a_n1756_n4888# 0.129341f
C179 minus.t8 a_n1756_n4888# 0.467527f
C180 minus.t3 a_n1756_n4888# 0.467527f
C181 minus.t4 a_n1756_n4888# 0.471025f
C182 minus.n3 a_n1756_n4888# 0.205677f
C183 minus.n4 a_n1756_n4888# 0.182204f
C184 minus.n5 a_n1756_n4888# 0.023473f
C185 minus.n6 a_n1756_n4888# 0.182204f
C186 minus.n7 a_n1756_n4888# 0.023473f
C187 minus.n8 a_n1756_n4888# 0.055332f
C188 minus.n9 a_n1756_n4888# 0.055332f
C189 minus.n10 a_n1756_n4888# 0.055332f
C190 minus.n11 a_n1756_n4888# 0.023473f
C191 minus.n12 a_n1756_n4888# 0.182204f
C192 minus.n13 a_n1756_n4888# 0.023473f
C193 minus.n14 a_n1756_n4888# 0.182204f
C194 minus.n15 a_n1756_n4888# 0.20559f
C195 minus.n16 a_n1756_n4888# 2.44482f
C196 minus.n17 a_n1756_n4888# 0.055332f
C197 minus.t12 a_n1756_n4888# 0.467527f
C198 minus.t6 a_n1756_n4888# 0.467527f
C199 minus.t1 a_n1756_n4888# 0.467527f
C200 minus.n18 a_n1756_n4888# 0.200559f
C201 minus.n19 a_n1756_n4888# 0.129341f
C202 minus.t13 a_n1756_n4888# 0.467527f
C203 minus.t10 a_n1756_n4888# 0.467527f
C204 minus.t2 a_n1756_n4888# 0.471025f
C205 minus.n20 a_n1756_n4888# 0.205677f
C206 minus.n21 a_n1756_n4888# 0.182204f
C207 minus.n22 a_n1756_n4888# 0.023473f
C208 minus.n23 a_n1756_n4888# 0.182204f
C209 minus.n24 a_n1756_n4888# 0.023473f
C210 minus.n25 a_n1756_n4888# 0.055332f
C211 minus.n26 a_n1756_n4888# 0.055332f
C212 minus.n27 a_n1756_n4888# 0.055332f
C213 minus.n28 a_n1756_n4888# 0.023473f
C214 minus.n29 a_n1756_n4888# 0.182204f
C215 minus.n30 a_n1756_n4888# 0.023473f
C216 minus.n31 a_n1756_n4888# 0.182204f
C217 minus.t0 a_n1756_n4888# 0.471025f
C218 minus.n32 a_n1756_n4888# 0.20559f
C219 minus.n33 a_n1756_n4888# 0.370918f
C220 minus.n34 a_n1756_n4888# 2.91815f
.ends

