* NGSPICE file created from diffpair641.ext - technology: sky130A

.subckt diffpair641 minus drain_right drain_left source plus
X0 drain_right minus source a_n1106_n5892# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X1 drain_left plus source a_n1106_n5892# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X2 drain_right minus source a_n1106_n5892# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X3 source plus drain_left a_n1106_n5892# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X4 a_n1106_n5892# a_n1106_n5892# a_n1106_n5892# a_n1106_n5892# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=95 ps=407.6 w=25 l=0.15
X5 source plus drain_left a_n1106_n5892# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X6 drain_left plus source a_n1106_n5892# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X7 source minus drain_right a_n1106_n5892# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X8 a_n1106_n5892# a_n1106_n5892# a_n1106_n5892# a_n1106_n5892# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X9 a_n1106_n5892# a_n1106_n5892# a_n1106_n5892# a_n1106_n5892# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X10 a_n1106_n5892# a_n1106_n5892# a_n1106_n5892# a_n1106_n5892# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X11 source minus drain_right a_n1106_n5892# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
.ends

