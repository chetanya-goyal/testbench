* NGSPICE file created from diffpair350.ext - technology: sky130A

.subckt diffpair350 minus drain_right drain_left source plus
X0 drain_right minus source a_n968_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=3.51 ps=18.78 w=9 l=0.3
X1 drain_left plus source a_n968_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=3.51 ps=18.78 w=9 l=0.3
X2 drain_right minus source a_n968_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=3.51 ps=18.78 w=9 l=0.3
X3 a_n968_n2692# a_n968_n2692# a_n968_n2692# a_n968_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.3
X4 drain_left plus source a_n968_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=3.51 ps=18.78 w=9 l=0.3
X5 a_n968_n2692# a_n968_n2692# a_n968_n2692# a_n968_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X6 a_n968_n2692# a_n968_n2692# a_n968_n2692# a_n968_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X7 a_n968_n2692# a_n968_n2692# a_n968_n2692# a_n968_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
.ends

