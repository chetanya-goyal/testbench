* NGSPICE file created from diffpair374.ext - technology: sky130A

.subckt diffpair374 minus drain_right drain_left source plus
X0 a_n1832_n2688# a_n1832_n2688# a_n1832_n2688# a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.6
X1 drain_right.t9 minus.t0 source.t11 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X2 drain_right.t8 minus.t1 source.t16 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X3 source.t1 plus.t0 drain_left.t9 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X4 a_n1832_n2688# a_n1832_n2688# a_n1832_n2688# a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X5 drain_right.t7 minus.t2 source.t9 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X6 drain_left.t8 plus.t1 source.t19 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X7 drain_left.t7 plus.t2 source.t3 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X8 source.t17 minus.t3 drain_right.t6 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X9 drain_right.t5 minus.t4 source.t12 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X10 source.t4 plus.t3 drain_left.t6 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X11 source.t13 minus.t5 drain_right.t4 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X12 drain_left.t5 plus.t4 source.t6 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X13 drain_right.t3 minus.t6 source.t14 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X14 source.t2 plus.t5 drain_left.t4 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X15 drain_left.t3 plus.t6 source.t18 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X16 source.t15 minus.t7 drain_right.t2 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X17 drain_left.t2 plus.t7 source.t5 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X18 source.t0 plus.t8 drain_left.t1 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X19 a_n1832_n2688# a_n1832_n2688# a_n1832_n2688# a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X20 drain_left.t0 plus.t9 source.t7 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X21 a_n1832_n2688# a_n1832_n2688# a_n1832_n2688# a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X22 drain_right.t1 minus.t8 source.t8 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X23 source.t10 minus.t9 drain_right.t0 a_n1832_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
R0 minus.n3 minus.t6 453.173
R1 minus.n13 minus.t2 453.173
R2 minus.n2 minus.t5 426.973
R3 minus.n1 minus.t4 426.973
R4 minus.n6 minus.t3 426.973
R5 minus.n8 minus.t1 426.973
R6 minus.n12 minus.t9 426.973
R7 minus.n11 minus.t0 426.973
R8 minus.n16 minus.t7 426.973
R9 minus.n18 minus.t8 426.973
R10 minus.n9 minus.n8 161.3
R11 minus.n7 minus.n0 161.3
R12 minus.n6 minus.n5 161.3
R13 minus.n19 minus.n18 161.3
R14 minus.n17 minus.n10 161.3
R15 minus.n16 minus.n15 161.3
R16 minus.n4 minus.n1 80.6037
R17 minus.n14 minus.n11 80.6037
R18 minus.n2 minus.n1 48.2005
R19 minus.n6 minus.n1 48.2005
R20 minus.n12 minus.n11 48.2005
R21 minus.n16 minus.n11 48.2005
R22 minus.n8 minus.n7 45.2793
R23 minus.n18 minus.n17 45.2793
R24 minus.n4 minus.n3 45.1669
R25 minus.n14 minus.n13 45.1669
R26 minus.n20 minus.n9 33.8888
R27 minus.n3 minus.n2 14.3992
R28 minus.n13 minus.n12 14.3992
R29 minus.n20 minus.n19 6.60088
R30 minus.n7 minus.n6 2.92171
R31 minus.n17 minus.n16 2.92171
R32 minus.n5 minus.n4 0.285035
R33 minus.n15 minus.n14 0.285035
R34 minus.n9 minus.n0 0.189894
R35 minus.n5 minus.n0 0.189894
R36 minus.n15 minus.n10 0.189894
R37 minus.n19 minus.n10 0.189894
R38 minus minus.n20 0.188
R39 source.n5 source.t14 51.0588
R40 source.n19 source.t8 51.0586
R41 source.n14 source.t5 51.0586
R42 source.n0 source.t19 51.0586
R43 source.n2 source.n1 48.8588
R44 source.n4 source.n3 48.8588
R45 source.n7 source.n6 48.8588
R46 source.n9 source.n8 48.8588
R47 source.n18 source.n17 48.8586
R48 source.n16 source.n15 48.8586
R49 source.n13 source.n12 48.8586
R50 source.n11 source.n10 48.8586
R51 source.n11 source.n9 20.6184
R52 source.n20 source.n0 14.1529
R53 source.n20 source.n19 5.66429
R54 source.n17 source.t11 2.2005
R55 source.n17 source.t15 2.2005
R56 source.n15 source.t9 2.2005
R57 source.n15 source.t10 2.2005
R58 source.n12 source.t3 2.2005
R59 source.n12 source.t1 2.2005
R60 source.n10 source.t7 2.2005
R61 source.n10 source.t0 2.2005
R62 source.n1 source.t6 2.2005
R63 source.n1 source.t4 2.2005
R64 source.n3 source.t18 2.2005
R65 source.n3 source.t2 2.2005
R66 source.n6 source.t12 2.2005
R67 source.n6 source.t13 2.2005
R68 source.n8 source.t16 2.2005
R69 source.n8 source.t17 2.2005
R70 source.n5 source.n4 0.87119
R71 source.n16 source.n14 0.87119
R72 source.n9 source.n7 0.802224
R73 source.n7 source.n5 0.802224
R74 source.n4 source.n2 0.802224
R75 source.n2 source.n0 0.802224
R76 source.n13 source.n11 0.802224
R77 source.n14 source.n13 0.802224
R78 source.n18 source.n16 0.802224
R79 source.n19 source.n18 0.802224
R80 source source.n20 0.188
R81 drain_right.n1 drain_right.t7 68.5391
R82 drain_right.n7 drain_right.t8 67.7376
R83 drain_right.n6 drain_right.n4 66.3391
R84 drain_right.n3 drain_right.n2 66.0833
R85 drain_right.n6 drain_right.n5 65.5376
R86 drain_right.n1 drain_right.n0 65.5373
R87 drain_right drain_right.n3 27.9484
R88 drain_right drain_right.n7 6.05408
R89 drain_right.n2 drain_right.t2 2.2005
R90 drain_right.n2 drain_right.t1 2.2005
R91 drain_right.n0 drain_right.t0 2.2005
R92 drain_right.n0 drain_right.t9 2.2005
R93 drain_right.n4 drain_right.t4 2.2005
R94 drain_right.n4 drain_right.t3 2.2005
R95 drain_right.n5 drain_right.t6 2.2005
R96 drain_right.n5 drain_right.t5 2.2005
R97 drain_right.n7 drain_right.n6 0.802224
R98 drain_right.n3 drain_right.n1 0.145585
R99 plus.n3 plus.t6 453.173
R100 plus.n13 plus.t7 453.173
R101 plus.n8 plus.t1 426.973
R102 plus.n6 plus.t3 426.973
R103 plus.n5 plus.t4 426.973
R104 plus.n4 plus.t5 426.973
R105 plus.n18 plus.t9 426.973
R106 plus.n16 plus.t8 426.973
R107 plus.n15 plus.t2 426.973
R108 plus.n14 plus.t0 426.973
R109 plus.n6 plus.n1 161.3
R110 plus.n7 plus.n0 161.3
R111 plus.n9 plus.n8 161.3
R112 plus.n16 plus.n11 161.3
R113 plus.n17 plus.n10 161.3
R114 plus.n19 plus.n18 161.3
R115 plus.n5 plus.n2 80.6037
R116 plus.n15 plus.n12 80.6037
R117 plus.n6 plus.n5 48.2005
R118 plus.n5 plus.n4 48.2005
R119 plus.n16 plus.n15 48.2005
R120 plus.n15 plus.n14 48.2005
R121 plus.n8 plus.n7 45.2793
R122 plus.n18 plus.n17 45.2793
R123 plus.n3 plus.n2 45.1669
R124 plus.n13 plus.n12 45.1669
R125 plus plus.n19 28.9062
R126 plus.n4 plus.n3 14.3992
R127 plus.n14 plus.n13 14.3992
R128 plus plus.n9 11.1085
R129 plus.n7 plus.n6 2.92171
R130 plus.n17 plus.n16 2.92171
R131 plus.n2 plus.n1 0.285035
R132 plus.n12 plus.n11 0.285035
R133 plus.n1 plus.n0 0.189894
R134 plus.n9 plus.n0 0.189894
R135 plus.n19 plus.n10 0.189894
R136 plus.n11 plus.n10 0.189894
R137 drain_left.n5 drain_left.t3 68.5393
R138 drain_left.n1 drain_left.t0 68.5391
R139 drain_left.n3 drain_left.n2 66.0833
R140 drain_left.n5 drain_left.n4 65.5376
R141 drain_left.n7 drain_left.n6 65.5374
R142 drain_left.n1 drain_left.n0 65.5373
R143 drain_left drain_left.n3 28.5017
R144 drain_left drain_left.n7 6.45494
R145 drain_left.n2 drain_left.t9 2.2005
R146 drain_left.n2 drain_left.t2 2.2005
R147 drain_left.n0 drain_left.t1 2.2005
R148 drain_left.n0 drain_left.t7 2.2005
R149 drain_left.n6 drain_left.t6 2.2005
R150 drain_left.n6 drain_left.t8 2.2005
R151 drain_left.n4 drain_left.t4 2.2005
R152 drain_left.n4 drain_left.t5 2.2005
R153 drain_left.n7 drain_left.n5 0.802224
R154 drain_left.n3 drain_left.n1 0.145585
C0 drain_right source 12.1373f
C1 drain_left plus 4.89939f
C2 drain_right plus 0.334433f
C3 drain_left drain_right 0.908917f
C4 minus source 4.61984f
C5 plus minus 4.87424f
C6 plus source 4.63427f
C7 drain_left minus 0.172117f
C8 drain_right minus 4.72344f
C9 drain_left source 12.1429f
C10 drain_right a_n1832_n2688# 6.03959f
C11 drain_left a_n1832_n2688# 6.32691f
C12 source a_n1832_n2688# 5.365478f
C13 minus a_n1832_n2688# 6.941984f
C14 plus a_n1832_n2688# 8.52905f
C15 drain_left.t0 a_n1832_n2688# 1.98592f
C16 drain_left.t1 a_n1832_n2688# 0.178016f
C17 drain_left.t7 a_n1832_n2688# 0.178016f
C18 drain_left.n0 a_n1832_n2688# 1.55705f
C19 drain_left.n1 a_n1832_n2688# 0.612723f
C20 drain_left.t9 a_n1832_n2688# 0.178016f
C21 drain_left.t2 a_n1832_n2688# 0.178016f
C22 drain_left.n2 a_n1832_n2688# 1.55969f
C23 drain_left.n3 a_n1832_n2688# 1.38685f
C24 drain_left.t3 a_n1832_n2688# 1.98592f
C25 drain_left.t4 a_n1832_n2688# 0.178016f
C26 drain_left.t5 a_n1832_n2688# 0.178016f
C27 drain_left.n4 a_n1832_n2688# 1.55705f
C28 drain_left.n5 a_n1832_n2688# 0.661677f
C29 drain_left.t6 a_n1832_n2688# 0.178016f
C30 drain_left.t8 a_n1832_n2688# 0.178016f
C31 drain_left.n6 a_n1832_n2688# 1.55704f
C32 drain_left.n7 a_n1832_n2688# 0.548081f
C33 plus.n0 a_n1832_n2688# 0.046089f
C34 plus.t1 a_n1832_n2688# 0.71376f
C35 plus.t3 a_n1832_n2688# 0.71376f
C36 plus.n1 a_n1832_n2688# 0.0615f
C37 plus.t4 a_n1832_n2688# 0.71376f
C38 plus.n2 a_n1832_n2688# 0.222771f
C39 plus.t5 a_n1832_n2688# 0.71376f
C40 plus.t6 a_n1832_n2688# 0.73122f
C41 plus.n3 a_n1832_n2688# 0.286782f
C42 plus.n4 a_n1832_n2688# 0.311796f
C43 plus.n5 a_n1832_n2688# 0.312569f
C44 plus.n6 a_n1832_n2688# 0.302679f
C45 plus.n7 a_n1832_n2688# 0.010459f
C46 plus.n8 a_n1832_n2688# 0.301542f
C47 plus.n9 a_n1832_n2688# 0.463979f
C48 plus.n10 a_n1832_n2688# 0.046089f
C49 plus.t9 a_n1832_n2688# 0.71376f
C50 plus.n11 a_n1832_n2688# 0.0615f
C51 plus.t8 a_n1832_n2688# 0.71376f
C52 plus.n12 a_n1832_n2688# 0.222771f
C53 plus.t2 a_n1832_n2688# 0.71376f
C54 plus.t7 a_n1832_n2688# 0.73122f
C55 plus.n13 a_n1832_n2688# 0.286782f
C56 plus.t0 a_n1832_n2688# 0.71376f
C57 plus.n14 a_n1832_n2688# 0.311796f
C58 plus.n15 a_n1832_n2688# 0.312569f
C59 plus.n16 a_n1832_n2688# 0.302679f
C60 plus.n17 a_n1832_n2688# 0.010459f
C61 plus.n18 a_n1832_n2688# 0.301542f
C62 plus.n19 a_n1832_n2688# 1.28429f
C63 drain_right.t7 a_n1832_n2688# 1.97392f
C64 drain_right.t0 a_n1832_n2688# 0.176941f
C65 drain_right.t9 a_n1832_n2688# 0.176941f
C66 drain_right.n0 a_n1832_n2688# 1.54764f
C67 drain_right.n1 a_n1832_n2688# 0.609022f
C68 drain_right.t2 a_n1832_n2688# 0.176941f
C69 drain_right.t1 a_n1832_n2688# 0.176941f
C70 drain_right.n2 a_n1832_n2688# 1.55027f
C71 drain_right.n3 a_n1832_n2688# 1.32724f
C72 drain_right.t4 a_n1832_n2688# 0.176941f
C73 drain_right.t3 a_n1832_n2688# 0.176941f
C74 drain_right.n4 a_n1832_n2688# 1.55172f
C75 drain_right.t6 a_n1832_n2688# 0.176941f
C76 drain_right.t5 a_n1832_n2688# 0.176941f
C77 drain_right.n5 a_n1832_n2688# 1.54765f
C78 drain_right.n6 a_n1832_n2688# 0.661588f
C79 drain_right.t8 a_n1832_n2688# 1.97002f
C80 drain_right.n7 a_n1832_n2688# 0.557179f
C81 source.t19 a_n1832_n2688# 2.01511f
C82 source.n0 a_n1832_n2688# 1.19578f
C83 source.t6 a_n1832_n2688# 0.188973f
C84 source.t4 a_n1832_n2688# 0.188973f
C85 source.n1 a_n1832_n2688# 1.58196f
C86 source.n2 a_n1832_n2688# 0.384926f
C87 source.t18 a_n1832_n2688# 0.188973f
C88 source.t2 a_n1832_n2688# 0.188973f
C89 source.n3 a_n1832_n2688# 1.58196f
C90 source.n4 a_n1832_n2688# 0.390831f
C91 source.t14 a_n1832_n2688# 2.01511f
C92 source.n5 a_n1832_n2688# 0.473058f
C93 source.t12 a_n1832_n2688# 0.188973f
C94 source.t13 a_n1832_n2688# 0.188973f
C95 source.n6 a_n1832_n2688# 1.58196f
C96 source.n7 a_n1832_n2688# 0.384926f
C97 source.t16 a_n1832_n2688# 0.188973f
C98 source.t17 a_n1832_n2688# 0.188973f
C99 source.n8 a_n1832_n2688# 1.58196f
C100 source.n9 a_n1832_n2688# 1.57551f
C101 source.t7 a_n1832_n2688# 0.188973f
C102 source.t0 a_n1832_n2688# 0.188973f
C103 source.n10 a_n1832_n2688# 1.58195f
C104 source.n11 a_n1832_n2688# 1.57551f
C105 source.t3 a_n1832_n2688# 0.188973f
C106 source.t1 a_n1832_n2688# 0.188973f
C107 source.n12 a_n1832_n2688# 1.58195f
C108 source.n13 a_n1832_n2688# 0.384931f
C109 source.t5 a_n1832_n2688# 2.01511f
C110 source.n14 a_n1832_n2688# 0.473063f
C111 source.t9 a_n1832_n2688# 0.188973f
C112 source.t10 a_n1832_n2688# 0.188973f
C113 source.n15 a_n1832_n2688# 1.58195f
C114 source.n16 a_n1832_n2688# 0.390835f
C115 source.t11 a_n1832_n2688# 0.188973f
C116 source.t15 a_n1832_n2688# 0.188973f
C117 source.n17 a_n1832_n2688# 1.58195f
C118 source.n18 a_n1832_n2688# 0.384931f
C119 source.t8 a_n1832_n2688# 2.01511f
C120 source.n19 a_n1832_n2688# 0.606281f
C121 source.n20 a_n1832_n2688# 1.39504f
C122 minus.n0 a_n1832_n2688# 0.045157f
C123 minus.t4 a_n1832_n2688# 0.69932f
C124 minus.n1 a_n1832_n2688# 0.306246f
C125 minus.t3 a_n1832_n2688# 0.69932f
C126 minus.t6 a_n1832_n2688# 0.716427f
C127 minus.t5 a_n1832_n2688# 0.69932f
C128 minus.n2 a_n1832_n2688# 0.305488f
C129 minus.n3 a_n1832_n2688# 0.28098f
C130 minus.n4 a_n1832_n2688# 0.218264f
C131 minus.n5 a_n1832_n2688# 0.060256f
C132 minus.n6 a_n1832_n2688# 0.296556f
C133 minus.n7 a_n1832_n2688# 0.010247f
C134 minus.t1 a_n1832_n2688# 0.69932f
C135 minus.n8 a_n1832_n2688# 0.295442f
C136 minus.n9 a_n1832_n2688# 1.44145f
C137 minus.n10 a_n1832_n2688# 0.045157f
C138 minus.t0 a_n1832_n2688# 0.69932f
C139 minus.n11 a_n1832_n2688# 0.306246f
C140 minus.t2 a_n1832_n2688# 0.716427f
C141 minus.t9 a_n1832_n2688# 0.69932f
C142 minus.n12 a_n1832_n2688# 0.305488f
C143 minus.n13 a_n1832_n2688# 0.28098f
C144 minus.n14 a_n1832_n2688# 0.218264f
C145 minus.n15 a_n1832_n2688# 0.060256f
C146 minus.t7 a_n1832_n2688# 0.69932f
C147 minus.n16 a_n1832_n2688# 0.296556f
C148 minus.n17 a_n1832_n2688# 0.010247f
C149 minus.t8 a_n1832_n2688# 0.69932f
C150 minus.n18 a_n1832_n2688# 0.295442f
C151 minus.n19 a_n1832_n2688# 0.305906f
C152 minus.n20 a_n1832_n2688# 1.7583f
.ends

