* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t9 plus.t0 source.t14 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X1 source.t6 minus.t0 drain_right.t9 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X2 drain_left.t8 plus.t1 source.t10 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X3 a_n1952_n1288# a_n1952_n1288# a_n1952_n1288# a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.7
X4 drain_left.t7 plus.t2 source.t12 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X5 drain_left.t6 plus.t3 source.t11 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X6 a_n1952_n1288# a_n1952_n1288# a_n1952_n1288# a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X7 drain_left.t5 plus.t4 source.t19 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X8 source.t17 plus.t5 drain_left.t4 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X9 drain_right.t8 minus.t1 source.t8 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X10 a_n1952_n1288# a_n1952_n1288# a_n1952_n1288# a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X11 drain_right.t7 minus.t2 source.t3 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X12 source.t15 plus.t6 drain_left.t3 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X13 source.t5 minus.t3 drain_right.t6 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X14 drain_right.t5 minus.t4 source.t7 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X15 drain_right.t4 minus.t5 source.t9 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X16 source.t16 plus.t7 drain_left.t2 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X17 source.t4 minus.t6 drain_right.t3 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X18 drain_right.t2 minus.t7 source.t1 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X19 drain_right.t1 minus.t8 source.t0 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X20 source.t18 plus.t8 drain_left.t1 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X21 drain_left.t0 plus.t9 source.t13 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X22 source.t2 minus.t9 drain_right.t0 a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X23 a_n1952_n1288# a_n1952_n1288# a_n1952_n1288# a_n1952_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
R0 plus.n6 plus.n5 161.3
R1 plus.n7 plus.n2 161.3
R2 plus.n9 plus.n8 161.3
R3 plus.n10 plus.n1 161.3
R4 plus.n11 plus.n0 161.3
R5 plus.n13 plus.n12 161.3
R6 plus.n20 plus.n19 161.3
R7 plus.n21 plus.n16 161.3
R8 plus.n23 plus.n22 161.3
R9 plus.n24 plus.n15 161.3
R10 plus.n25 plus.n14 161.3
R11 plus.n27 plus.n26 161.3
R12 plus.n3 plus.t3 147.725
R13 plus.n17 plus.t9 147.725
R14 plus.n12 plus.t2 124.977
R15 plus.n10 plus.t6 124.977
R16 plus.n2 plus.t0 124.977
R17 plus.n4 plus.t7 124.977
R18 plus.n26 plus.t4 124.977
R19 plus.n24 plus.t5 124.977
R20 plus.n16 plus.t1 124.977
R21 plus.n18 plus.t8 124.977
R22 plus.n6 plus.n3 44.8741
R23 plus.n20 plus.n17 44.8741
R24 plus.n12 plus.n11 30.6732
R25 plus.n26 plus.n25 30.6732
R26 plus plus.n27 26.7471
R27 plus.n10 plus.n9 26.2914
R28 plus.n5 plus.n4 26.2914
R29 plus.n24 plus.n23 26.2914
R30 plus.n19 plus.n18 26.2914
R31 plus.n9 plus.n2 21.9096
R32 plus.n5 plus.n2 21.9096
R33 plus.n23 plus.n16 21.9096
R34 plus.n19 plus.n16 21.9096
R35 plus.n4 plus.n3 19.0667
R36 plus.n18 plus.n17 19.0667
R37 plus.n11 plus.n10 17.5278
R38 plus.n25 plus.n24 17.5278
R39 plus plus.n13 8.49482
R40 plus.n7 plus.n6 0.189894
R41 plus.n8 plus.n7 0.189894
R42 plus.n8 plus.n1 0.189894
R43 plus.n1 plus.n0 0.189894
R44 plus.n13 plus.n0 0.189894
R45 plus.n27 plus.n14 0.189894
R46 plus.n15 plus.n14 0.189894
R47 plus.n22 plus.n15 0.189894
R48 plus.n22 plus.n21 0.189894
R49 plus.n21 plus.n20 0.189894
R50 source.n42 source.n40 289.615
R51 source.n30 source.n28 289.615
R52 source.n2 source.n0 289.615
R53 source.n14 source.n12 289.615
R54 source.n43 source.n42 185
R55 source.n31 source.n30 185
R56 source.n3 source.n2 185
R57 source.n15 source.n14 185
R58 source.t0 source.n41 167.117
R59 source.t13 source.n29 167.117
R60 source.t12 source.n1 167.117
R61 source.t7 source.n13 167.117
R62 source.n9 source.n8 84.1169
R63 source.n11 source.n10 84.1169
R64 source.n21 source.n20 84.1169
R65 source.n23 source.n22 84.1169
R66 source.n39 source.n38 84.1168
R67 source.n37 source.n36 84.1168
R68 source.n27 source.n26 84.1168
R69 source.n25 source.n24 84.1168
R70 source.n42 source.t0 52.3082
R71 source.n30 source.t13 52.3082
R72 source.n2 source.t12 52.3082
R73 source.n14 source.t7 52.3082
R74 source.n47 source.n46 31.4096
R75 source.n35 source.n34 31.4096
R76 source.n7 source.n6 31.4096
R77 source.n19 source.n18 31.4096
R78 source.n25 source.n23 15.4878
R79 source.n38 source.t1 9.9005
R80 source.n38 source.t4 9.9005
R81 source.n36 source.t9 9.9005
R82 source.n36 source.t5 9.9005
R83 source.n26 source.t10 9.9005
R84 source.n26 source.t18 9.9005
R85 source.n24 source.t19 9.9005
R86 source.n24 source.t17 9.9005
R87 source.n8 source.t14 9.9005
R88 source.n8 source.t15 9.9005
R89 source.n10 source.t11 9.9005
R90 source.n10 source.t16 9.9005
R91 source.n20 source.t3 9.9005
R92 source.n20 source.t6 9.9005
R93 source.n22 source.t8 9.9005
R94 source.n22 source.t2 9.9005
R95 source.n43 source.n41 9.71174
R96 source.n31 source.n29 9.71174
R97 source.n3 source.n1 9.71174
R98 source.n15 source.n13 9.71174
R99 source.n46 source.n45 9.45567
R100 source.n34 source.n33 9.45567
R101 source.n6 source.n5 9.45567
R102 source.n18 source.n17 9.45567
R103 source.n45 source.n44 9.3005
R104 source.n33 source.n32 9.3005
R105 source.n5 source.n4 9.3005
R106 source.n17 source.n16 9.3005
R107 source.n48 source.n7 8.893
R108 source.n46 source.n40 8.14595
R109 source.n34 source.n28 8.14595
R110 source.n6 source.n0 8.14595
R111 source.n18 source.n12 8.14595
R112 source.n44 source.n43 7.3702
R113 source.n32 source.n31 7.3702
R114 source.n4 source.n3 7.3702
R115 source.n16 source.n15 7.3702
R116 source.n44 source.n40 5.81868
R117 source.n32 source.n28 5.81868
R118 source.n4 source.n0 5.81868
R119 source.n16 source.n12 5.81868
R120 source.n48 source.n47 5.7074
R121 source.n45 source.n41 3.44771
R122 source.n33 source.n29 3.44771
R123 source.n5 source.n1 3.44771
R124 source.n17 source.n13 3.44771
R125 source.n19 source.n11 0.914293
R126 source.n37 source.n35 0.914293
R127 source.n23 source.n21 0.888431
R128 source.n21 source.n19 0.888431
R129 source.n11 source.n9 0.888431
R130 source.n9 source.n7 0.888431
R131 source.n27 source.n25 0.888431
R132 source.n35 source.n27 0.888431
R133 source.n39 source.n37 0.888431
R134 source.n47 source.n39 0.888431
R135 source source.n48 0.188
R136 drain_left.n2 drain_left.n0 289.615
R137 drain_left.n13 drain_left.n11 289.615
R138 drain_left.n3 drain_left.n2 185
R139 drain_left.n14 drain_left.n13 185
R140 drain_left.t5 drain_left.n1 167.117
R141 drain_left.t6 drain_left.n12 167.117
R142 drain_left.n10 drain_left.n9 101.406
R143 drain_left.n21 drain_left.n20 100.796
R144 drain_left.n19 drain_left.n18 100.796
R145 drain_left.n8 drain_left.n7 100.796
R146 drain_left.n2 drain_left.t5 52.3082
R147 drain_left.n13 drain_left.t6 52.3082
R148 drain_left.n8 drain_left.n6 48.9763
R149 drain_left.n19 drain_left.n17 48.9763
R150 drain_left drain_left.n10 23.565
R151 drain_left.n9 drain_left.t1 9.9005
R152 drain_left.n9 drain_left.t0 9.9005
R153 drain_left.n7 drain_left.t4 9.9005
R154 drain_left.n7 drain_left.t8 9.9005
R155 drain_left.n20 drain_left.t3 9.9005
R156 drain_left.n20 drain_left.t7 9.9005
R157 drain_left.n18 drain_left.t2 9.9005
R158 drain_left.n18 drain_left.t9 9.9005
R159 drain_left.n3 drain_left.n1 9.71174
R160 drain_left.n14 drain_left.n12 9.71174
R161 drain_left.n6 drain_left.n5 9.45567
R162 drain_left.n17 drain_left.n16 9.45567
R163 drain_left.n5 drain_left.n4 9.3005
R164 drain_left.n16 drain_left.n15 9.3005
R165 drain_left.n6 drain_left.n0 8.14595
R166 drain_left.n17 drain_left.n11 8.14595
R167 drain_left.n4 drain_left.n3 7.3702
R168 drain_left.n15 drain_left.n14 7.3702
R169 drain_left drain_left.n21 6.54115
R170 drain_left.n4 drain_left.n0 5.81868
R171 drain_left.n15 drain_left.n11 5.81868
R172 drain_left.n5 drain_left.n1 3.44771
R173 drain_left.n16 drain_left.n12 3.44771
R174 drain_left.n21 drain_left.n19 0.888431
R175 drain_left.n10 drain_left.n8 0.167137
R176 minus.n13 minus.n12 161.3
R177 minus.n11 minus.n0 161.3
R178 minus.n10 minus.n9 161.3
R179 minus.n8 minus.n1 161.3
R180 minus.n7 minus.n6 161.3
R181 minus.n5 minus.n2 161.3
R182 minus.n27 minus.n26 161.3
R183 minus.n25 minus.n14 161.3
R184 minus.n24 minus.n23 161.3
R185 minus.n22 minus.n15 161.3
R186 minus.n21 minus.n20 161.3
R187 minus.n19 minus.n16 161.3
R188 minus.n3 minus.t4 147.725
R189 minus.n17 minus.t5 147.725
R190 minus.n4 minus.t0 124.977
R191 minus.n6 minus.t2 124.977
R192 minus.n10 minus.t9 124.977
R193 minus.n12 minus.t1 124.977
R194 minus.n18 minus.t3 124.977
R195 minus.n20 minus.t7 124.977
R196 minus.n24 minus.t6 124.977
R197 minus.n26 minus.t8 124.977
R198 minus.n3 minus.n2 44.8741
R199 minus.n17 minus.n16 44.8741
R200 minus.n12 minus.n11 30.6732
R201 minus.n26 minus.n25 30.6732
R202 minus.n28 minus.n13 29.0782
R203 minus.n5 minus.n4 26.2914
R204 minus.n10 minus.n1 26.2914
R205 minus.n19 minus.n18 26.2914
R206 minus.n24 minus.n15 26.2914
R207 minus.n6 minus.n5 21.9096
R208 minus.n6 minus.n1 21.9096
R209 minus.n20 minus.n19 21.9096
R210 minus.n20 minus.n15 21.9096
R211 minus.n4 minus.n3 19.0667
R212 minus.n18 minus.n17 19.0667
R213 minus.n11 minus.n10 17.5278
R214 minus.n25 minus.n24 17.5278
R215 minus.n28 minus.n27 6.63876
R216 minus.n13 minus.n0 0.189894
R217 minus.n9 minus.n0 0.189894
R218 minus.n9 minus.n8 0.189894
R219 minus.n8 minus.n7 0.189894
R220 minus.n7 minus.n2 0.189894
R221 minus.n21 minus.n16 0.189894
R222 minus.n22 minus.n21 0.189894
R223 minus.n23 minus.n22 0.189894
R224 minus.n23 minus.n14 0.189894
R225 minus.n27 minus.n14 0.189894
R226 minus minus.n28 0.188
R227 drain_right.n2 drain_right.n0 289.615
R228 drain_right.n16 drain_right.n14 289.615
R229 drain_right.n3 drain_right.n2 185
R230 drain_right.n17 drain_right.n16 185
R231 drain_right.t4 drain_right.n1 167.117
R232 drain_right.t8 drain_right.n15 167.117
R233 drain_right.n13 drain_right.n11 101.683
R234 drain_right.n10 drain_right.n9 101.406
R235 drain_right.n13 drain_right.n12 100.796
R236 drain_right.n8 drain_right.n7 100.796
R237 drain_right.n2 drain_right.t4 52.3082
R238 drain_right.n16 drain_right.t8 52.3082
R239 drain_right.n8 drain_right.n6 48.9763
R240 drain_right.n21 drain_right.n20 48.0884
R241 drain_right drain_right.n10 23.0118
R242 drain_right.n9 drain_right.t3 9.9005
R243 drain_right.n9 drain_right.t1 9.9005
R244 drain_right.n7 drain_right.t6 9.9005
R245 drain_right.n7 drain_right.t2 9.9005
R246 drain_right.n11 drain_right.t9 9.9005
R247 drain_right.n11 drain_right.t5 9.9005
R248 drain_right.n12 drain_right.t0 9.9005
R249 drain_right.n12 drain_right.t7 9.9005
R250 drain_right.n3 drain_right.n1 9.71174
R251 drain_right.n17 drain_right.n15 9.71174
R252 drain_right.n6 drain_right.n5 9.45567
R253 drain_right.n20 drain_right.n19 9.45567
R254 drain_right.n5 drain_right.n4 9.3005
R255 drain_right.n19 drain_right.n18 9.3005
R256 drain_right.n6 drain_right.n0 8.14595
R257 drain_right.n20 drain_right.n14 8.14595
R258 drain_right.n4 drain_right.n3 7.3702
R259 drain_right.n18 drain_right.n17 7.3702
R260 drain_right drain_right.n21 6.09718
R261 drain_right.n4 drain_right.n0 5.81868
R262 drain_right.n18 drain_right.n14 5.81868
R263 drain_right.n5 drain_right.n1 3.44771
R264 drain_right.n19 drain_right.n15 3.44771
R265 drain_right.n21 drain_right.n13 0.888431
R266 drain_right.n10 drain_right.n8 0.167137
C0 plus minus 3.73292f
C1 drain_left source 4.53542f
C2 drain_right source 4.53523f
C3 drain_left drain_right 0.965971f
C4 plus source 1.86166f
C5 drain_left plus 1.6793f
C6 drain_right plus 0.352787f
C7 minus source 1.84762f
C8 drain_left minus 0.178286f
C9 drain_right minus 1.48947f
C10 drain_right a_n1952_n1288# 3.772876f
C11 drain_left a_n1952_n1288# 4.03083f
C12 source a_n1952_n1288# 2.611252f
C13 minus a_n1952_n1288# 6.811874f
C14 plus a_n1952_n1288# 7.337094f
C15 drain_right.n0 a_n1952_n1288# 0.026677f
C16 drain_right.n1 a_n1952_n1288# 0.059027f
C17 drain_right.t4 a_n1952_n1288# 0.044297f
C18 drain_right.n2 a_n1952_n1288# 0.046197f
C19 drain_right.n3 a_n1952_n1288# 0.014892f
C20 drain_right.n4 a_n1952_n1288# 0.009822f
C21 drain_right.n5 a_n1952_n1288# 0.13011f
C22 drain_right.n6 a_n1952_n1288# 0.043449f
C23 drain_right.t6 a_n1952_n1288# 0.028887f
C24 drain_right.t2 a_n1952_n1288# 0.028887f
C25 drain_right.n7 a_n1952_n1288# 0.181477f
C26 drain_right.n8 a_n1952_n1288# 0.289888f
C27 drain_right.t3 a_n1952_n1288# 0.028887f
C28 drain_right.t1 a_n1952_n1288# 0.028887f
C29 drain_right.n9 a_n1952_n1288# 0.1829f
C30 drain_right.n10 a_n1952_n1288# 0.755753f
C31 drain_right.t9 a_n1952_n1288# 0.028887f
C32 drain_right.t5 a_n1952_n1288# 0.028887f
C33 drain_right.n11 a_n1952_n1288# 0.183677f
C34 drain_right.t0 a_n1952_n1288# 0.028887f
C35 drain_right.t7 a_n1952_n1288# 0.028887f
C36 drain_right.n12 a_n1952_n1288# 0.181478f
C37 drain_right.n13 a_n1952_n1288# 0.494129f
C38 drain_right.n14 a_n1952_n1288# 0.026677f
C39 drain_right.n15 a_n1952_n1288# 0.059027f
C40 drain_right.t8 a_n1952_n1288# 0.044297f
C41 drain_right.n16 a_n1952_n1288# 0.046197f
C42 drain_right.n17 a_n1952_n1288# 0.014892f
C43 drain_right.n18 a_n1952_n1288# 0.009822f
C44 drain_right.n19 a_n1952_n1288# 0.13011f
C45 drain_right.n20 a_n1952_n1288# 0.041873f
C46 drain_right.n21 a_n1952_n1288# 0.254899f
C47 minus.n0 a_n1952_n1288# 0.02399f
C48 minus.n1 a_n1952_n1288# 0.005444f
C49 minus.t9 a_n1952_n1288# 0.104006f
C50 minus.n2 a_n1952_n1288# 0.100201f
C51 minus.t4 a_n1952_n1288# 0.115126f
C52 minus.n3 a_n1952_n1288# 0.063365f
C53 minus.t0 a_n1952_n1288# 0.104006f
C54 minus.n4 a_n1952_n1288# 0.074715f
C55 minus.n5 a_n1952_n1288# 0.005444f
C56 minus.t2 a_n1952_n1288# 0.104006f
C57 minus.n6 a_n1952_n1288# 0.072298f
C58 minus.n7 a_n1952_n1288# 0.02399f
C59 minus.n8 a_n1952_n1288# 0.02399f
C60 minus.n9 a_n1952_n1288# 0.02399f
C61 minus.n10 a_n1952_n1288# 0.072298f
C62 minus.n11 a_n1952_n1288# 0.005444f
C63 minus.t1 a_n1952_n1288# 0.104006f
C64 minus.n12 a_n1952_n1288# 0.070967f
C65 minus.n13 a_n1952_n1288# 0.594631f
C66 minus.n14 a_n1952_n1288# 0.02399f
C67 minus.n15 a_n1952_n1288# 0.005444f
C68 minus.n16 a_n1952_n1288# 0.100201f
C69 minus.t5 a_n1952_n1288# 0.115126f
C70 minus.n17 a_n1952_n1288# 0.063365f
C71 minus.t3 a_n1952_n1288# 0.104006f
C72 minus.n18 a_n1952_n1288# 0.074715f
C73 minus.n19 a_n1952_n1288# 0.005444f
C74 minus.t7 a_n1952_n1288# 0.104006f
C75 minus.n20 a_n1952_n1288# 0.072298f
C76 minus.n21 a_n1952_n1288# 0.02399f
C77 minus.n22 a_n1952_n1288# 0.02399f
C78 minus.n23 a_n1952_n1288# 0.02399f
C79 minus.t6 a_n1952_n1288# 0.104006f
C80 minus.n24 a_n1952_n1288# 0.072298f
C81 minus.n25 a_n1952_n1288# 0.005444f
C82 minus.t8 a_n1952_n1288# 0.104006f
C83 minus.n26 a_n1952_n1288# 0.070967f
C84 minus.n27 a_n1952_n1288# 0.164631f
C85 minus.n28 a_n1952_n1288# 0.730412f
C86 drain_left.n0 a_n1952_n1288# 0.02626f
C87 drain_left.n1 a_n1952_n1288# 0.058104f
C88 drain_left.t5 a_n1952_n1288# 0.043604f
C89 drain_left.n2 a_n1952_n1288# 0.045474f
C90 drain_left.n3 a_n1952_n1288# 0.014659f
C91 drain_left.n4 a_n1952_n1288# 0.009668f
C92 drain_left.n5 a_n1952_n1288# 0.128075f
C93 drain_left.n6 a_n1952_n1288# 0.042769f
C94 drain_left.t4 a_n1952_n1288# 0.028435f
C95 drain_left.t8 a_n1952_n1288# 0.028435f
C96 drain_left.n7 a_n1952_n1288# 0.178639f
C97 drain_left.n8 a_n1952_n1288# 0.285355f
C98 drain_left.t1 a_n1952_n1288# 0.028435f
C99 drain_left.t0 a_n1952_n1288# 0.028435f
C100 drain_left.n9 a_n1952_n1288# 0.180039f
C101 drain_left.n10 a_n1952_n1288# 0.77915f
C102 drain_left.n11 a_n1952_n1288# 0.02626f
C103 drain_left.n12 a_n1952_n1288# 0.058104f
C104 drain_left.t6 a_n1952_n1288# 0.043604f
C105 drain_left.n13 a_n1952_n1288# 0.045474f
C106 drain_left.n14 a_n1952_n1288# 0.014659f
C107 drain_left.n15 a_n1952_n1288# 0.009668f
C108 drain_left.n16 a_n1952_n1288# 0.128075f
C109 drain_left.n17 a_n1952_n1288# 0.042769f
C110 drain_left.t2 a_n1952_n1288# 0.028435f
C111 drain_left.t9 a_n1952_n1288# 0.028435f
C112 drain_left.n18 a_n1952_n1288# 0.17864f
C113 drain_left.n19 a_n1952_n1288# 0.324667f
C114 drain_left.t3 a_n1952_n1288# 0.028435f
C115 drain_left.t7 a_n1952_n1288# 0.028435f
C116 drain_left.n20 a_n1952_n1288# 0.17864f
C117 drain_left.n21 a_n1952_n1288# 0.399798f
C118 source.n0 a_n1952_n1288# 0.033279f
C119 source.n1 a_n1952_n1288# 0.073634f
C120 source.t12 a_n1952_n1288# 0.055259f
C121 source.n2 a_n1952_n1288# 0.057629f
C122 source.n3 a_n1952_n1288# 0.018577f
C123 source.n4 a_n1952_n1288# 0.012252f
C124 source.n5 a_n1952_n1288# 0.162308f
C125 source.n6 a_n1952_n1288# 0.036482f
C126 source.n7 a_n1952_n1288# 0.389142f
C127 source.t14 a_n1952_n1288# 0.036036f
C128 source.t15 a_n1952_n1288# 0.036036f
C129 source.n8 a_n1952_n1288# 0.192647f
C130 source.n9 a_n1952_n1288# 0.307738f
C131 source.t11 a_n1952_n1288# 0.036036f
C132 source.t16 a_n1952_n1288# 0.036036f
C133 source.n10 a_n1952_n1288# 0.192647f
C134 source.n11 a_n1952_n1288# 0.309638f
C135 source.n12 a_n1952_n1288# 0.033279f
C136 source.n13 a_n1952_n1288# 0.073634f
C137 source.t7 a_n1952_n1288# 0.055259f
C138 source.n14 a_n1952_n1288# 0.057629f
C139 source.n15 a_n1952_n1288# 0.018577f
C140 source.n16 a_n1952_n1288# 0.012252f
C141 source.n17 a_n1952_n1288# 0.162308f
C142 source.n18 a_n1952_n1288# 0.036482f
C143 source.n19 a_n1952_n1288# 0.151142f
C144 source.t3 a_n1952_n1288# 0.036036f
C145 source.t6 a_n1952_n1288# 0.036036f
C146 source.n20 a_n1952_n1288# 0.192647f
C147 source.n21 a_n1952_n1288# 0.307738f
C148 source.t8 a_n1952_n1288# 0.036036f
C149 source.t2 a_n1952_n1288# 0.036036f
C150 source.n22 a_n1952_n1288# 0.192647f
C151 source.n23 a_n1952_n1288# 0.831229f
C152 source.t19 a_n1952_n1288# 0.036036f
C153 source.t17 a_n1952_n1288# 0.036036f
C154 source.n24 a_n1952_n1288# 0.192646f
C155 source.n25 a_n1952_n1288# 0.83123f
C156 source.t10 a_n1952_n1288# 0.036036f
C157 source.t18 a_n1952_n1288# 0.036036f
C158 source.n26 a_n1952_n1288# 0.192646f
C159 source.n27 a_n1952_n1288# 0.307739f
C160 source.n28 a_n1952_n1288# 0.033279f
C161 source.n29 a_n1952_n1288# 0.073634f
C162 source.t13 a_n1952_n1288# 0.055259f
C163 source.n30 a_n1952_n1288# 0.057629f
C164 source.n31 a_n1952_n1288# 0.018577f
C165 source.n32 a_n1952_n1288# 0.012252f
C166 source.n33 a_n1952_n1288# 0.162308f
C167 source.n34 a_n1952_n1288# 0.036482f
C168 source.n35 a_n1952_n1288# 0.151142f
C169 source.t9 a_n1952_n1288# 0.036036f
C170 source.t5 a_n1952_n1288# 0.036036f
C171 source.n36 a_n1952_n1288# 0.192646f
C172 source.n37 a_n1952_n1288# 0.309639f
C173 source.t1 a_n1952_n1288# 0.036036f
C174 source.t4 a_n1952_n1288# 0.036036f
C175 source.n38 a_n1952_n1288# 0.192646f
C176 source.n39 a_n1952_n1288# 0.307739f
C177 source.n40 a_n1952_n1288# 0.033279f
C178 source.n41 a_n1952_n1288# 0.073634f
C179 source.t0 a_n1952_n1288# 0.055259f
C180 source.n42 a_n1952_n1288# 0.057629f
C181 source.n43 a_n1952_n1288# 0.018577f
C182 source.n44 a_n1952_n1288# 0.012252f
C183 source.n45 a_n1952_n1288# 0.162308f
C184 source.n46 a_n1952_n1288# 0.036482f
C185 source.n47 a_n1952_n1288# 0.267255f
C186 source.n48 a_n1952_n1288# 0.574816f
C187 plus.n0 a_n1952_n1288# 0.024309f
C188 plus.t2 a_n1952_n1288# 0.105388f
C189 plus.t6 a_n1952_n1288# 0.105388f
C190 plus.n1 a_n1952_n1288# 0.024309f
C191 plus.t0 a_n1952_n1288# 0.105388f
C192 plus.n2 a_n1952_n1288# 0.073259f
C193 plus.t3 a_n1952_n1288# 0.116656f
C194 plus.n3 a_n1952_n1288# 0.064207f
C195 plus.t7 a_n1952_n1288# 0.105388f
C196 plus.n4 a_n1952_n1288# 0.075708f
C197 plus.n5 a_n1952_n1288# 0.005516f
C198 plus.n6 a_n1952_n1288# 0.101532f
C199 plus.n7 a_n1952_n1288# 0.024309f
C200 plus.n8 a_n1952_n1288# 0.024309f
C201 plus.n9 a_n1952_n1288# 0.005516f
C202 plus.n10 a_n1952_n1288# 0.073259f
C203 plus.n11 a_n1952_n1288# 0.005516f
C204 plus.n12 a_n1952_n1288# 0.07191f
C205 plus.n13 a_n1952_n1288# 0.182106f
C206 plus.n14 a_n1952_n1288# 0.024309f
C207 plus.t4 a_n1952_n1288# 0.105388f
C208 plus.n15 a_n1952_n1288# 0.024309f
C209 plus.t5 a_n1952_n1288# 0.105388f
C210 plus.t1 a_n1952_n1288# 0.105388f
C211 plus.n16 a_n1952_n1288# 0.073259f
C212 plus.t9 a_n1952_n1288# 0.116656f
C213 plus.n17 a_n1952_n1288# 0.064207f
C214 plus.t8 a_n1952_n1288# 0.105388f
C215 plus.n18 a_n1952_n1288# 0.075708f
C216 plus.n19 a_n1952_n1288# 0.005516f
C217 plus.n20 a_n1952_n1288# 0.101532f
C218 plus.n21 a_n1952_n1288# 0.024309f
C219 plus.n22 a_n1952_n1288# 0.024309f
C220 plus.n23 a_n1952_n1288# 0.005516f
C221 plus.n24 a_n1952_n1288# 0.073259f
C222 plus.n25 a_n1952_n1288# 0.005516f
C223 plus.n26 a_n1952_n1288# 0.07191f
C224 plus.n27 a_n1952_n1288# 0.575041f
.ends

