* NGSPICE file created from diffpair35.ext - technology: sky130A

.subckt diffpair35 minus drain_right drain_left source plus
X0 drain_left.t11 plus.t0 source.t12 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X1 source.t7 minus.t0 drain_right.t11 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X2 drain_right.t10 minus.t1 source.t10 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X3 source.t0 minus.t2 drain_right.t9 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X4 source.t13 plus.t1 drain_left.t10 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X5 source.t19 plus.t2 drain_left.t9 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X6 a_n1598_n1088# a_n1598_n1088# a_n1598_n1088# a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.3
X7 source.t16 plus.t3 drain_left.t8 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X8 drain_right.t8 minus.t3 source.t11 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X9 drain_right.t7 minus.t4 source.t1 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X10 drain_left.t7 plus.t4 source.t23 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X11 a_n1598_n1088# a_n1598_n1088# a_n1598_n1088# a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X12 a_n1598_n1088# a_n1598_n1088# a_n1598_n1088# a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X13 source.t6 minus.t5 drain_right.t6 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X14 source.t17 plus.t5 drain_left.t6 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X15 drain_left.t5 plus.t6 source.t20 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X16 drain_left.t4 plus.t7 source.t22 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X17 source.t9 minus.t6 drain_right.t5 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X18 drain_right.t4 minus.t7 source.t3 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X19 source.t5 minus.t8 drain_right.t3 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X20 drain_left.t3 plus.t8 source.t18 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X21 source.t21 plus.t9 drain_left.t2 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X22 source.t15 plus.t10 drain_left.t1 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X23 drain_right.t2 minus.t9 source.t8 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X24 drain_right.t1 minus.t10 source.t2 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X25 source.t4 minus.t11 drain_right.t0 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X26 a_n1598_n1088# a_n1598_n1088# a_n1598_n1088# a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X27 drain_left.t0 plus.t11 source.t14 a_n1598_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
R0 plus.n2 plus.t3 232.237
R1 plus.n13 plus.t8 232.237
R2 plus.n17 plus.t7 232.237
R3 plus.n28 plus.t2 232.237
R4 plus.n3 plus.t6 184.768
R5 plus.n4 plus.t10 184.768
R6 plus.n10 plus.t11 184.768
R7 plus.n12 plus.t5 184.768
R8 plus.n19 plus.t1 184.768
R9 plus.n18 plus.t0 184.768
R10 plus.n25 plus.t9 184.768
R11 plus.n27 plus.t4 184.768
R12 plus.n6 plus.n2 161.489
R13 plus.n21 plus.n17 161.489
R14 plus.n6 plus.n5 161.3
R15 plus.n7 plus.n1 161.3
R16 plus.n9 plus.n8 161.3
R17 plus.n11 plus.n0 161.3
R18 plus.n14 plus.n13 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n22 plus.n16 161.3
R21 plus.n24 plus.n23 161.3
R22 plus.n26 plus.n15 161.3
R23 plus.n29 plus.n28 161.3
R24 plus.n9 plus.n1 73.0308
R25 plus.n24 plus.n16 73.0308
R26 plus.n5 plus.n4 63.5369
R27 plus.n11 plus.n10 63.5369
R28 plus.n26 plus.n25 63.5369
R29 plus.n20 plus.n18 63.5369
R30 plus.n3 plus.n2 44.549
R31 plus.n13 plus.n12 44.549
R32 plus.n28 plus.n27 44.549
R33 plus.n19 plus.n17 44.549
R34 plus.n5 plus.n3 28.4823
R35 plus.n12 plus.n11 28.4823
R36 plus.n27 plus.n26 28.4823
R37 plus.n20 plus.n19 28.4823
R38 plus plus.n29 24.9005
R39 plus.n4 plus.n1 9.49444
R40 plus.n10 plus.n9 9.49444
R41 plus.n25 plus.n24 9.49444
R42 plus.n18 plus.n16 9.49444
R43 plus plus.n14 7.98914
R44 plus.n7 plus.n6 0.189894
R45 plus.n8 plus.n7 0.189894
R46 plus.n8 plus.n0 0.189894
R47 plus.n14 plus.n0 0.189894
R48 plus.n29 plus.n15 0.189894
R49 plus.n23 plus.n15 0.189894
R50 plus.n23 plus.n22 0.189894
R51 plus.n22 plus.n21 0.189894
R52 source.n0 source.t18 243.255
R53 source.n5 source.t16 243.255
R54 source.n6 source.t3 243.255
R55 source.n11 source.t7 243.255
R56 source.n23 source.t1 243.254
R57 source.n18 source.t5 243.254
R58 source.n17 source.t22 243.254
R59 source.n12 source.t19 243.254
R60 source.n2 source.n1 223.454
R61 source.n4 source.n3 223.454
R62 source.n8 source.n7 223.454
R63 source.n10 source.n9 223.454
R64 source.n22 source.n21 223.453
R65 source.n20 source.n19 223.453
R66 source.n16 source.n15 223.453
R67 source.n14 source.n13 223.453
R68 source.n21 source.t8 19.8005
R69 source.n21 source.t6 19.8005
R70 source.n19 source.t11 19.8005
R71 source.n19 source.t0 19.8005
R72 source.n15 source.t12 19.8005
R73 source.n15 source.t13 19.8005
R74 source.n13 source.t23 19.8005
R75 source.n13 source.t21 19.8005
R76 source.n1 source.t14 19.8005
R77 source.n1 source.t17 19.8005
R78 source.n3 source.t20 19.8005
R79 source.n3 source.t15 19.8005
R80 source.n7 source.t10 19.8005
R81 source.n7 source.t4 19.8005
R82 source.n9 source.t2 19.8005
R83 source.n9 source.t9 19.8005
R84 source.n12 source.n11 13.4975
R85 source.n24 source.n0 7.96301
R86 source.n24 source.n23 5.53498
R87 source.n11 source.n10 0.543603
R88 source.n10 source.n8 0.543603
R89 source.n8 source.n6 0.543603
R90 source.n5 source.n4 0.543603
R91 source.n4 source.n2 0.543603
R92 source.n2 source.n0 0.543603
R93 source.n14 source.n12 0.543603
R94 source.n16 source.n14 0.543603
R95 source.n17 source.n16 0.543603
R96 source.n20 source.n18 0.543603
R97 source.n22 source.n20 0.543603
R98 source.n23 source.n22 0.543603
R99 source.n6 source.n5 0.470328
R100 source.n18 source.n17 0.470328
R101 source source.n24 0.188
R102 drain_left.n6 drain_left.n4 240.675
R103 drain_left.n3 drain_left.n2 240.619
R104 drain_left.n3 drain_left.n0 240.619
R105 drain_left.n8 drain_left.n7 240.132
R106 drain_left.n6 drain_left.n5 240.132
R107 drain_left.n3 drain_left.n1 240.131
R108 drain_left drain_left.n3 21.7493
R109 drain_left.n1 drain_left.t2 19.8005
R110 drain_left.n1 drain_left.t11 19.8005
R111 drain_left.n2 drain_left.t10 19.8005
R112 drain_left.n2 drain_left.t4 19.8005
R113 drain_left.n0 drain_left.t9 19.8005
R114 drain_left.n0 drain_left.t7 19.8005
R115 drain_left.n7 drain_left.t6 19.8005
R116 drain_left.n7 drain_left.t3 19.8005
R117 drain_left.n5 drain_left.t1 19.8005
R118 drain_left.n5 drain_left.t0 19.8005
R119 drain_left.n4 drain_left.t8 19.8005
R120 drain_left.n4 drain_left.t5 19.8005
R121 drain_left drain_left.n8 6.19632
R122 drain_left.n8 drain_left.n6 0.543603
R123 minus.n13 minus.t0 232.237
R124 minus.n2 minus.t7 232.237
R125 minus.n28 minus.t4 232.237
R126 minus.n17 minus.t8 232.237
R127 minus.n12 minus.t10 184.768
R128 minus.n10 minus.t6 184.768
R129 minus.n3 minus.t1 184.768
R130 minus.n4 minus.t11 184.768
R131 minus.n27 minus.t5 184.768
R132 minus.n25 minus.t9 184.768
R133 minus.n19 minus.t2 184.768
R134 minus.n18 minus.t3 184.768
R135 minus.n6 minus.n2 161.489
R136 minus.n21 minus.n17 161.489
R137 minus.n14 minus.n13 161.3
R138 minus.n11 minus.n0 161.3
R139 minus.n9 minus.n8 161.3
R140 minus.n7 minus.n1 161.3
R141 minus.n6 minus.n5 161.3
R142 minus.n29 minus.n28 161.3
R143 minus.n26 minus.n15 161.3
R144 minus.n24 minus.n23 161.3
R145 minus.n22 minus.n16 161.3
R146 minus.n21 minus.n20 161.3
R147 minus.n9 minus.n1 73.0308
R148 minus.n24 minus.n16 73.0308
R149 minus.n11 minus.n10 63.5369
R150 minus.n5 minus.n3 63.5369
R151 minus.n20 minus.n19 63.5369
R152 minus.n26 minus.n25 63.5369
R153 minus.n13 minus.n12 44.549
R154 minus.n4 minus.n2 44.549
R155 minus.n18 minus.n17 44.549
R156 minus.n28 minus.n27 44.549
R157 minus.n12 minus.n11 28.4823
R158 minus.n5 minus.n4 28.4823
R159 minus.n20 minus.n18 28.4823
R160 minus.n27 minus.n26 28.4823
R161 minus.n30 minus.n14 26.8528
R162 minus.n10 minus.n9 9.49444
R163 minus.n3 minus.n1 9.49444
R164 minus.n19 minus.n16 9.49444
R165 minus.n25 minus.n24 9.49444
R166 minus.n30 minus.n29 6.51186
R167 minus.n14 minus.n0 0.189894
R168 minus.n8 minus.n0 0.189894
R169 minus.n8 minus.n7 0.189894
R170 minus.n7 minus.n6 0.189894
R171 minus.n22 minus.n21 0.189894
R172 minus.n23 minus.n22 0.189894
R173 minus.n23 minus.n15 0.189894
R174 minus.n29 minus.n15 0.189894
R175 minus minus.n30 0.188
R176 drain_right.n6 drain_right.n4 240.675
R177 drain_right.n3 drain_right.n2 240.619
R178 drain_right.n3 drain_right.n0 240.619
R179 drain_right.n6 drain_right.n5 240.132
R180 drain_right.n8 drain_right.n7 240.132
R181 drain_right.n3 drain_right.n1 240.131
R182 drain_right drain_right.n3 21.196
R183 drain_right.n1 drain_right.t9 19.8005
R184 drain_right.n1 drain_right.t2 19.8005
R185 drain_right.n2 drain_right.t6 19.8005
R186 drain_right.n2 drain_right.t7 19.8005
R187 drain_right.n0 drain_right.t3 19.8005
R188 drain_right.n0 drain_right.t8 19.8005
R189 drain_right.n4 drain_right.t0 19.8005
R190 drain_right.n4 drain_right.t4 19.8005
R191 drain_right.n5 drain_right.t5 19.8005
R192 drain_right.n5 drain_right.t10 19.8005
R193 drain_right.n7 drain_right.t11 19.8005
R194 drain_right.n7 drain_right.t1 19.8005
R195 drain_right drain_right.n8 6.19632
R196 drain_right.n8 drain_right.n6 0.543603
C0 minus drain_left 0.178004f
C1 plus drain_left 0.945804f
C2 minus drain_right 0.792406f
C3 plus drain_right 0.315444f
C4 source drain_left 4.08036f
C5 minus plus 3.11588f
C6 source drain_right 4.08011f
C7 source minus 1.01439f
C8 source plus 1.02826f
C9 drain_right drain_left 0.786281f
C10 drain_right a_n1598_n1088# 3.26591f
C11 drain_left a_n1598_n1088# 3.47665f
C12 source a_n1598_n1088# 2.405054f
C13 minus a_n1598_n1088# 5.299895f
C14 plus a_n1598_n1088# 5.975736f
C15 drain_right.t3 a_n1598_n1088# 0.01935f
C16 drain_right.t8 a_n1598_n1088# 0.01935f
C17 drain_right.n0 a_n1598_n1088# 0.075721f
C18 drain_right.t9 a_n1598_n1088# 0.01935f
C19 drain_right.t2 a_n1598_n1088# 0.01935f
C20 drain_right.n1 a_n1598_n1088# 0.075187f
C21 drain_right.t6 a_n1598_n1088# 0.01935f
C22 drain_right.t7 a_n1598_n1088# 0.01935f
C23 drain_right.n2 a_n1598_n1088# 0.075721f
C24 drain_right.n3 a_n1598_n1088# 1.29569f
C25 drain_right.t0 a_n1598_n1088# 0.01935f
C26 drain_right.t4 a_n1598_n1088# 0.01935f
C27 drain_right.n4 a_n1598_n1088# 0.075789f
C28 drain_right.t5 a_n1598_n1088# 0.01935f
C29 drain_right.t10 a_n1598_n1088# 0.01935f
C30 drain_right.n5 a_n1598_n1088# 0.075187f
C31 drain_right.n6 a_n1598_n1088# 0.523129f
C32 drain_right.t11 a_n1598_n1088# 0.01935f
C33 drain_right.t1 a_n1598_n1088# 0.01935f
C34 drain_right.n7 a_n1598_n1088# 0.075187f
C35 drain_right.n8 a_n1598_n1088# 0.460746f
C36 minus.n0 a_n1598_n1088# 0.033236f
C37 minus.t0 a_n1598_n1088# 0.037734f
C38 minus.t10 a_n1598_n1088# 0.030737f
C39 minus.t6 a_n1598_n1088# 0.030737f
C40 minus.n1 a_n1598_n1088# 0.012357f
C41 minus.t7 a_n1598_n1088# 0.037734f
C42 minus.n2 a_n1598_n1088# 0.040972f
C43 minus.t1 a_n1598_n1088# 0.030737f
C44 minus.n3 a_n1598_n1088# 0.031668f
C45 minus.t11 a_n1598_n1088# 0.030737f
C46 minus.n4 a_n1598_n1088# 0.031668f
C47 minus.n5 a_n1598_n1088# 0.013689f
C48 minus.n6 a_n1598_n1088# 0.075643f
C49 minus.n7 a_n1598_n1088# 0.033236f
C50 minus.n8 a_n1598_n1088# 0.033236f
C51 minus.n9 a_n1598_n1088# 0.012357f
C52 minus.n10 a_n1598_n1088# 0.031668f
C53 minus.n11 a_n1598_n1088# 0.013689f
C54 minus.n12 a_n1598_n1088# 0.031668f
C55 minus.n13 a_n1598_n1088# 0.040923f
C56 minus.n14 a_n1598_n1088# 0.711937f
C57 minus.n15 a_n1598_n1088# 0.033236f
C58 minus.t5 a_n1598_n1088# 0.030737f
C59 minus.t9 a_n1598_n1088# 0.030737f
C60 minus.n16 a_n1598_n1088# 0.012357f
C61 minus.t8 a_n1598_n1088# 0.037734f
C62 minus.n17 a_n1598_n1088# 0.040972f
C63 minus.t3 a_n1598_n1088# 0.030737f
C64 minus.n18 a_n1598_n1088# 0.031668f
C65 minus.t2 a_n1598_n1088# 0.030737f
C66 minus.n19 a_n1598_n1088# 0.031668f
C67 minus.n20 a_n1598_n1088# 0.013689f
C68 minus.n21 a_n1598_n1088# 0.075643f
C69 minus.n22 a_n1598_n1088# 0.033236f
C70 minus.n23 a_n1598_n1088# 0.033236f
C71 minus.n24 a_n1598_n1088# 0.012357f
C72 minus.n25 a_n1598_n1088# 0.031668f
C73 minus.n26 a_n1598_n1088# 0.013689f
C74 minus.n27 a_n1598_n1088# 0.031668f
C75 minus.t4 a_n1598_n1088# 0.037734f
C76 minus.n28 a_n1598_n1088# 0.040923f
C77 minus.n29 a_n1598_n1088# 0.218217f
C78 minus.n30 a_n1598_n1088# 0.879162f
C79 drain_left.t9 a_n1598_n1088# 0.018908f
C80 drain_left.t7 a_n1598_n1088# 0.018908f
C81 drain_left.n0 a_n1598_n1088# 0.073992f
C82 drain_left.t2 a_n1598_n1088# 0.018908f
C83 drain_left.t11 a_n1598_n1088# 0.018908f
C84 drain_left.n1 a_n1598_n1088# 0.07347f
C85 drain_left.t10 a_n1598_n1088# 0.018908f
C86 drain_left.t4 a_n1598_n1088# 0.018908f
C87 drain_left.n2 a_n1598_n1088# 0.073992f
C88 drain_left.n3 a_n1598_n1088# 1.31243f
C89 drain_left.t8 a_n1598_n1088# 0.018908f
C90 drain_left.t5 a_n1598_n1088# 0.018908f
C91 drain_left.n4 a_n1598_n1088# 0.074059f
C92 drain_left.t1 a_n1598_n1088# 0.018908f
C93 drain_left.t0 a_n1598_n1088# 0.018908f
C94 drain_left.n5 a_n1598_n1088# 0.07347f
C95 drain_left.n6 a_n1598_n1088# 0.511186f
C96 drain_left.t6 a_n1598_n1088# 0.018908f
C97 drain_left.t3 a_n1598_n1088# 0.018908f
C98 drain_left.n7 a_n1598_n1088# 0.07347f
C99 drain_left.n8 a_n1598_n1088# 0.450228f
C100 source.t18 a_n1598_n1088# 0.122525f
C101 source.n0 a_n1598_n1088# 0.526104f
C102 source.t14 a_n1598_n1088# 0.022014f
C103 source.t17 a_n1598_n1088# 0.022014f
C104 source.n1 a_n1598_n1088# 0.071394f
C105 source.n2 a_n1598_n1088# 0.268592f
C106 source.t20 a_n1598_n1088# 0.022014f
C107 source.t15 a_n1598_n1088# 0.022014f
C108 source.n3 a_n1598_n1088# 0.071394f
C109 source.n4 a_n1598_n1088# 0.268592f
C110 source.t16 a_n1598_n1088# 0.122525f
C111 source.n5 a_n1598_n1088# 0.27092f
C112 source.t3 a_n1598_n1088# 0.122525f
C113 source.n6 a_n1598_n1088# 0.27092f
C114 source.t10 a_n1598_n1088# 0.022014f
C115 source.t4 a_n1598_n1088# 0.022014f
C116 source.n7 a_n1598_n1088# 0.071394f
C117 source.n8 a_n1598_n1088# 0.268592f
C118 source.t2 a_n1598_n1088# 0.022014f
C119 source.t9 a_n1598_n1088# 0.022014f
C120 source.n9 a_n1598_n1088# 0.071394f
C121 source.n10 a_n1598_n1088# 0.268592f
C122 source.t7 a_n1598_n1088# 0.122525f
C123 source.n11 a_n1598_n1088# 0.749326f
C124 source.t19 a_n1598_n1088# 0.122525f
C125 source.n12 a_n1598_n1088# 0.749326f
C126 source.t23 a_n1598_n1088# 0.022014f
C127 source.t21 a_n1598_n1088# 0.022014f
C128 source.n13 a_n1598_n1088# 0.071394f
C129 source.n14 a_n1598_n1088# 0.268592f
C130 source.t12 a_n1598_n1088# 0.022014f
C131 source.t13 a_n1598_n1088# 0.022014f
C132 source.n15 a_n1598_n1088# 0.071394f
C133 source.n16 a_n1598_n1088# 0.268592f
C134 source.t22 a_n1598_n1088# 0.122525f
C135 source.n17 a_n1598_n1088# 0.27092f
C136 source.t5 a_n1598_n1088# 0.122525f
C137 source.n18 a_n1598_n1088# 0.27092f
C138 source.t11 a_n1598_n1088# 0.022014f
C139 source.t0 a_n1598_n1088# 0.022014f
C140 source.n19 a_n1598_n1088# 0.071394f
C141 source.n20 a_n1598_n1088# 0.268592f
C142 source.t8 a_n1598_n1088# 0.022014f
C143 source.t6 a_n1598_n1088# 0.022014f
C144 source.n21 a_n1598_n1088# 0.071394f
C145 source.n22 a_n1598_n1088# 0.268592f
C146 source.t1 a_n1598_n1088# 0.122525f
C147 source.n23 a_n1598_n1088# 0.428175f
C148 source.n24 a_n1598_n1088# 0.564187f
C149 plus.n0 a_n1598_n1088# 0.033972f
C150 plus.t5 a_n1598_n1088# 0.031418f
C151 plus.t11 a_n1598_n1088# 0.031418f
C152 plus.n1 a_n1598_n1088# 0.012631f
C153 plus.t3 a_n1598_n1088# 0.03857f
C154 plus.n2 a_n1598_n1088# 0.04188f
C155 plus.t6 a_n1598_n1088# 0.031418f
C156 plus.n3 a_n1598_n1088# 0.03237f
C157 plus.t10 a_n1598_n1088# 0.031418f
C158 plus.n4 a_n1598_n1088# 0.03237f
C159 plus.n5 a_n1598_n1088# 0.013993f
C160 plus.n6 a_n1598_n1088# 0.07732f
C161 plus.n7 a_n1598_n1088# 0.033972f
C162 plus.n8 a_n1598_n1088# 0.033972f
C163 plus.n9 a_n1598_n1088# 0.012631f
C164 plus.n10 a_n1598_n1088# 0.03237f
C165 plus.n11 a_n1598_n1088# 0.013993f
C166 plus.n12 a_n1598_n1088# 0.03237f
C167 plus.t8 a_n1598_n1088# 0.03857f
C168 plus.n13 a_n1598_n1088# 0.041829f
C169 plus.n14 a_n1598_n1088# 0.233915f
C170 plus.n15 a_n1598_n1088# 0.033972f
C171 plus.t2 a_n1598_n1088# 0.03857f
C172 plus.t4 a_n1598_n1088# 0.031418f
C173 plus.t9 a_n1598_n1088# 0.031418f
C174 plus.n16 a_n1598_n1088# 0.012631f
C175 plus.t7 a_n1598_n1088# 0.03857f
C176 plus.n17 a_n1598_n1088# 0.04188f
C177 plus.t0 a_n1598_n1088# 0.031418f
C178 plus.n18 a_n1598_n1088# 0.03237f
C179 plus.t1 a_n1598_n1088# 0.031418f
C180 plus.n19 a_n1598_n1088# 0.03237f
C181 plus.n20 a_n1598_n1088# 0.013993f
C182 plus.n21 a_n1598_n1088# 0.07732f
C183 plus.n22 a_n1598_n1088# 0.033972f
C184 plus.n23 a_n1598_n1088# 0.033972f
C185 plus.n24 a_n1598_n1088# 0.012631f
C186 plus.n25 a_n1598_n1088# 0.03237f
C187 plus.n26 a_n1598_n1088# 0.013993f
C188 plus.n27 a_n1598_n1088# 0.03237f
C189 plus.n28 a_n1598_n1088# 0.041829f
C190 plus.n29 a_n1598_n1088# 0.708f
.ends

