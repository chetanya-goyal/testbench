* NGSPICE file created from diffpair469.ext - technology: sky130A

.subckt diffpair469 minus drain_right drain_left source plus
X0 source.t47 minus.t0 drain_right.t15 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X1 a_n3394_n3288# a_n3394_n3288# a_n3394_n3288# a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.7
X2 drain_right.t14 minus.t1 source.t46 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X3 source.t10 plus.t0 drain_left.t23 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X4 drain_left.t22 plus.t1 source.t23 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X5 drain_left.t21 plus.t2 source.t22 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X6 source.t12 plus.t3 drain_left.t20 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X7 source.t45 minus.t2 drain_right.t19 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X8 source.t11 plus.t4 drain_left.t19 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X9 source.t44 minus.t3 drain_right.t18 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X10 drain_right.t3 minus.t4 source.t43 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X11 drain_left.t18 plus.t5 source.t13 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X12 source.t17 plus.t6 drain_left.t17 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X13 source.t0 plus.t7 drain_left.t16 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X14 drain_right.t2 minus.t5 source.t42 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X15 drain_right.t23 minus.t6 source.t41 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X16 drain_right.t22 minus.t7 source.t40 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X17 a_n3394_n3288# a_n3394_n3288# a_n3394_n3288# a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X18 drain_right.t9 minus.t8 source.t39 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X19 source.t20 plus.t8 drain_left.t15 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X20 drain_right.t8 minus.t9 source.t38 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X21 drain_left.t14 plus.t9 source.t1 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X22 drain_left.t13 plus.t10 source.t14 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X23 drain_right.t1 minus.t10 source.t37 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X24 drain_left.t12 plus.t11 source.t16 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X25 source.t36 minus.t11 drain_right.t0 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X26 drain_right.t7 minus.t12 source.t35 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X27 source.t9 plus.t12 drain_left.t11 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X28 drain_left.t10 plus.t13 source.t15 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X29 drain_left.t9 plus.t14 source.t2 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X30 drain_right.t6 minus.t13 source.t34 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X31 a_n3394_n3288# a_n3394_n3288# a_n3394_n3288# a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X32 source.t8 plus.t15 drain_left.t8 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X33 drain_left.t7 plus.t16 source.t19 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X34 source.t7 plus.t17 drain_left.t6 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X35 drain_left.t5 plus.t18 source.t5 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X36 source.t33 minus.t14 drain_right.t5 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.7
X37 drain_left.t4 plus.t19 source.t4 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X38 a_n3394_n3288# a_n3394_n3288# a_n3394_n3288# a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X39 source.t32 minus.t15 drain_right.t4 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X40 drain_right.t11 minus.t16 source.t31 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X41 source.t30 minus.t17 drain_right.t10 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X42 source.t21 plus.t20 drain_left.t3 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X43 source.t29 minus.t18 drain_right.t13 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X44 drain_left.t2 plus.t21 source.t18 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.7
X45 source.t28 minus.t19 drain_right.t12 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X46 source.t3 plus.t22 drain_left.t1 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X47 drain_right.t17 minus.t20 source.t27 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X48 source.t26 minus.t21 drain_right.t16 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X49 source.t25 minus.t22 drain_right.t21 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X50 source.t6 plus.t23 drain_left.t0 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
X51 source.t24 minus.t23 drain_right.t20 a_n3394_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.7
R0 minus.n11 minus.t13 495.62
R1 minus.n53 minus.t2 495.62
R2 minus.n10 minus.t3 469.262
R3 minus.n14 minus.t10 469.262
R4 minus.n16 minus.t21 469.262
R5 minus.n20 minus.t9 469.262
R6 minus.n22 minus.t22 469.262
R7 minus.n26 minus.t8 469.262
R8 minus.n28 minus.t18 469.262
R9 minus.n32 minus.t7 469.262
R10 minus.n34 minus.t15 469.262
R11 minus.n38 minus.t5 469.262
R12 minus.n40 minus.t14 469.262
R13 minus.n52 minus.t4 469.262
R14 minus.n56 minus.t19 469.262
R15 minus.n58 minus.t20 469.262
R16 minus.n62 minus.t23 469.262
R17 minus.n64 minus.t16 469.262
R18 minus.n68 minus.t17 469.262
R19 minus.n70 minus.t12 469.262
R20 minus.n74 minus.t11 469.262
R21 minus.n76 minus.t6 469.262
R22 minus.n80 minus.t0 469.262
R23 minus.n82 minus.t1 469.262
R24 minus.n41 minus.n40 161.3
R25 minus.n39 minus.n0 161.3
R26 minus.n38 minus.n37 161.3
R27 minus.n36 minus.n1 161.3
R28 minus.n35 minus.n34 161.3
R29 minus.n33 minus.n2 161.3
R30 minus.n32 minus.n31 161.3
R31 minus.n30 minus.n3 161.3
R32 minus.n29 minus.n28 161.3
R33 minus.n27 minus.n4 161.3
R34 minus.n26 minus.n25 161.3
R35 minus.n24 minus.n5 161.3
R36 minus.n23 minus.n22 161.3
R37 minus.n21 minus.n6 161.3
R38 minus.n20 minus.n19 161.3
R39 minus.n18 minus.n7 161.3
R40 minus.n17 minus.n16 161.3
R41 minus.n15 minus.n8 161.3
R42 minus.n14 minus.n13 161.3
R43 minus.n12 minus.n9 161.3
R44 minus.n83 minus.n82 161.3
R45 minus.n81 minus.n42 161.3
R46 minus.n80 minus.n79 161.3
R47 minus.n78 minus.n43 161.3
R48 minus.n77 minus.n76 161.3
R49 minus.n75 minus.n44 161.3
R50 minus.n74 minus.n73 161.3
R51 minus.n72 minus.n45 161.3
R52 minus.n71 minus.n70 161.3
R53 minus.n69 minus.n46 161.3
R54 minus.n68 minus.n67 161.3
R55 minus.n66 minus.n47 161.3
R56 minus.n65 minus.n64 161.3
R57 minus.n63 minus.n48 161.3
R58 minus.n62 minus.n61 161.3
R59 minus.n60 minus.n49 161.3
R60 minus.n59 minus.n58 161.3
R61 minus.n57 minus.n50 161.3
R62 minus.n56 minus.n55 161.3
R63 minus.n54 minus.n51 161.3
R64 minus.n40 minus.n39 46.0096
R65 minus.n82 minus.n81 46.0096
R66 minus.n12 minus.n11 45.0871
R67 minus.n54 minus.n53 45.0871
R68 minus.n84 minus.n41 42.1558
R69 minus.n10 minus.n9 41.6278
R70 minus.n38 minus.n1 41.6278
R71 minus.n52 minus.n51 41.6278
R72 minus.n80 minus.n43 41.6278
R73 minus.n15 minus.n14 37.246
R74 minus.n34 minus.n33 37.246
R75 minus.n57 minus.n56 37.246
R76 minus.n76 minus.n75 37.246
R77 minus.n16 minus.n7 32.8641
R78 minus.n32 minus.n3 32.8641
R79 minus.n58 minus.n49 32.8641
R80 minus.n74 minus.n45 32.8641
R81 minus.n21 minus.n20 28.4823
R82 minus.n28 minus.n27 28.4823
R83 minus.n63 minus.n62 28.4823
R84 minus.n70 minus.n69 28.4823
R85 minus.n26 minus.n5 24.1005
R86 minus.n22 minus.n5 24.1005
R87 minus.n64 minus.n47 24.1005
R88 minus.n68 minus.n47 24.1005
R89 minus.n22 minus.n21 19.7187
R90 minus.n27 minus.n26 19.7187
R91 minus.n64 minus.n63 19.7187
R92 minus.n69 minus.n68 19.7187
R93 minus.n20 minus.n7 15.3369
R94 minus.n28 minus.n3 15.3369
R95 minus.n62 minus.n49 15.3369
R96 minus.n70 minus.n45 15.3369
R97 minus.n11 minus.n10 14.1472
R98 minus.n53 minus.n52 14.1472
R99 minus.n16 minus.n15 10.955
R100 minus.n33 minus.n32 10.955
R101 minus.n58 minus.n57 10.955
R102 minus.n75 minus.n74 10.955
R103 minus.n84 minus.n83 6.67853
R104 minus.n14 minus.n9 6.57323
R105 minus.n34 minus.n1 6.57323
R106 minus.n56 minus.n51 6.57323
R107 minus.n76 minus.n43 6.57323
R108 minus.n39 minus.n38 2.19141
R109 minus.n81 minus.n80 2.19141
R110 minus.n41 minus.n0 0.189894
R111 minus.n37 minus.n0 0.189894
R112 minus.n37 minus.n36 0.189894
R113 minus.n36 minus.n35 0.189894
R114 minus.n35 minus.n2 0.189894
R115 minus.n31 minus.n2 0.189894
R116 minus.n31 minus.n30 0.189894
R117 minus.n30 minus.n29 0.189894
R118 minus.n29 minus.n4 0.189894
R119 minus.n25 minus.n4 0.189894
R120 minus.n25 minus.n24 0.189894
R121 minus.n24 minus.n23 0.189894
R122 minus.n23 minus.n6 0.189894
R123 minus.n19 minus.n6 0.189894
R124 minus.n19 minus.n18 0.189894
R125 minus.n18 minus.n17 0.189894
R126 minus.n17 minus.n8 0.189894
R127 minus.n13 minus.n8 0.189894
R128 minus.n13 minus.n12 0.189894
R129 minus.n55 minus.n54 0.189894
R130 minus.n55 minus.n50 0.189894
R131 minus.n59 minus.n50 0.189894
R132 minus.n60 minus.n59 0.189894
R133 minus.n61 minus.n60 0.189894
R134 minus.n61 minus.n48 0.189894
R135 minus.n65 minus.n48 0.189894
R136 minus.n66 minus.n65 0.189894
R137 minus.n67 minus.n66 0.189894
R138 minus.n67 minus.n46 0.189894
R139 minus.n71 minus.n46 0.189894
R140 minus.n72 minus.n71 0.189894
R141 minus.n73 minus.n72 0.189894
R142 minus.n73 minus.n44 0.189894
R143 minus.n77 minus.n44 0.189894
R144 minus.n78 minus.n77 0.189894
R145 minus.n79 minus.n78 0.189894
R146 minus.n79 minus.n42 0.189894
R147 minus.n83 minus.n42 0.189894
R148 minus minus.n84 0.188
R149 drain_right.n7 drain_right.n5 60.4404
R150 drain_right.n2 drain_right.n0 60.4404
R151 drain_right.n13 drain_right.n11 60.4404
R152 drain_right.n13 drain_right.n12 59.5527
R153 drain_right.n15 drain_right.n14 59.5527
R154 drain_right.n17 drain_right.n16 59.5527
R155 drain_right.n19 drain_right.n18 59.5527
R156 drain_right.n21 drain_right.n20 59.5527
R157 drain_right.n7 drain_right.n6 59.5525
R158 drain_right.n9 drain_right.n8 59.5525
R159 drain_right.n4 drain_right.n3 59.5525
R160 drain_right.n2 drain_right.n1 59.5525
R161 drain_right drain_right.n10 35.2492
R162 drain_right drain_right.n21 6.54115
R163 drain_right.n5 drain_right.t15 1.6505
R164 drain_right.n5 drain_right.t14 1.6505
R165 drain_right.n6 drain_right.t0 1.6505
R166 drain_right.n6 drain_right.t23 1.6505
R167 drain_right.n8 drain_right.t10 1.6505
R168 drain_right.n8 drain_right.t7 1.6505
R169 drain_right.n3 drain_right.t20 1.6505
R170 drain_right.n3 drain_right.t11 1.6505
R171 drain_right.n1 drain_right.t12 1.6505
R172 drain_right.n1 drain_right.t17 1.6505
R173 drain_right.n0 drain_right.t19 1.6505
R174 drain_right.n0 drain_right.t3 1.6505
R175 drain_right.n11 drain_right.t18 1.6505
R176 drain_right.n11 drain_right.t6 1.6505
R177 drain_right.n12 drain_right.t16 1.6505
R178 drain_right.n12 drain_right.t1 1.6505
R179 drain_right.n14 drain_right.t21 1.6505
R180 drain_right.n14 drain_right.t8 1.6505
R181 drain_right.n16 drain_right.t13 1.6505
R182 drain_right.n16 drain_right.t9 1.6505
R183 drain_right.n18 drain_right.t4 1.6505
R184 drain_right.n18 drain_right.t22 1.6505
R185 drain_right.n20 drain_right.t5 1.6505
R186 drain_right.n20 drain_right.t2 1.6505
R187 drain_right.n9 drain_right.n7 0.888431
R188 drain_right.n4 drain_right.n2 0.888431
R189 drain_right.n21 drain_right.n19 0.888431
R190 drain_right.n19 drain_right.n17 0.888431
R191 drain_right.n17 drain_right.n15 0.888431
R192 drain_right.n15 drain_right.n13 0.888431
R193 drain_right.n10 drain_right.n9 0.389119
R194 drain_right.n10 drain_right.n4 0.389119
R195 source.n562 source.n502 289.615
R196 source.n486 source.n426 289.615
R197 source.n420 source.n360 289.615
R198 source.n344 source.n284 289.615
R199 source.n60 source.n0 289.615
R200 source.n136 source.n76 289.615
R201 source.n202 source.n142 289.615
R202 source.n278 source.n218 289.615
R203 source.n522 source.n521 185
R204 source.n527 source.n526 185
R205 source.n529 source.n528 185
R206 source.n518 source.n517 185
R207 source.n535 source.n534 185
R208 source.n537 source.n536 185
R209 source.n514 source.n513 185
R210 source.n544 source.n543 185
R211 source.n545 source.n512 185
R212 source.n547 source.n546 185
R213 source.n510 source.n509 185
R214 source.n553 source.n552 185
R215 source.n555 source.n554 185
R216 source.n506 source.n505 185
R217 source.n561 source.n560 185
R218 source.n563 source.n562 185
R219 source.n446 source.n445 185
R220 source.n451 source.n450 185
R221 source.n453 source.n452 185
R222 source.n442 source.n441 185
R223 source.n459 source.n458 185
R224 source.n461 source.n460 185
R225 source.n438 source.n437 185
R226 source.n468 source.n467 185
R227 source.n469 source.n436 185
R228 source.n471 source.n470 185
R229 source.n434 source.n433 185
R230 source.n477 source.n476 185
R231 source.n479 source.n478 185
R232 source.n430 source.n429 185
R233 source.n485 source.n484 185
R234 source.n487 source.n486 185
R235 source.n380 source.n379 185
R236 source.n385 source.n384 185
R237 source.n387 source.n386 185
R238 source.n376 source.n375 185
R239 source.n393 source.n392 185
R240 source.n395 source.n394 185
R241 source.n372 source.n371 185
R242 source.n402 source.n401 185
R243 source.n403 source.n370 185
R244 source.n405 source.n404 185
R245 source.n368 source.n367 185
R246 source.n411 source.n410 185
R247 source.n413 source.n412 185
R248 source.n364 source.n363 185
R249 source.n419 source.n418 185
R250 source.n421 source.n420 185
R251 source.n304 source.n303 185
R252 source.n309 source.n308 185
R253 source.n311 source.n310 185
R254 source.n300 source.n299 185
R255 source.n317 source.n316 185
R256 source.n319 source.n318 185
R257 source.n296 source.n295 185
R258 source.n326 source.n325 185
R259 source.n327 source.n294 185
R260 source.n329 source.n328 185
R261 source.n292 source.n291 185
R262 source.n335 source.n334 185
R263 source.n337 source.n336 185
R264 source.n288 source.n287 185
R265 source.n343 source.n342 185
R266 source.n345 source.n344 185
R267 source.n61 source.n60 185
R268 source.n59 source.n58 185
R269 source.n4 source.n3 185
R270 source.n53 source.n52 185
R271 source.n51 source.n50 185
R272 source.n8 source.n7 185
R273 source.n45 source.n44 185
R274 source.n43 source.n10 185
R275 source.n42 source.n41 185
R276 source.n13 source.n11 185
R277 source.n36 source.n35 185
R278 source.n34 source.n33 185
R279 source.n17 source.n16 185
R280 source.n28 source.n27 185
R281 source.n26 source.n25 185
R282 source.n21 source.n20 185
R283 source.n137 source.n136 185
R284 source.n135 source.n134 185
R285 source.n80 source.n79 185
R286 source.n129 source.n128 185
R287 source.n127 source.n126 185
R288 source.n84 source.n83 185
R289 source.n121 source.n120 185
R290 source.n119 source.n86 185
R291 source.n118 source.n117 185
R292 source.n89 source.n87 185
R293 source.n112 source.n111 185
R294 source.n110 source.n109 185
R295 source.n93 source.n92 185
R296 source.n104 source.n103 185
R297 source.n102 source.n101 185
R298 source.n97 source.n96 185
R299 source.n203 source.n202 185
R300 source.n201 source.n200 185
R301 source.n146 source.n145 185
R302 source.n195 source.n194 185
R303 source.n193 source.n192 185
R304 source.n150 source.n149 185
R305 source.n187 source.n186 185
R306 source.n185 source.n152 185
R307 source.n184 source.n183 185
R308 source.n155 source.n153 185
R309 source.n178 source.n177 185
R310 source.n176 source.n175 185
R311 source.n159 source.n158 185
R312 source.n170 source.n169 185
R313 source.n168 source.n167 185
R314 source.n163 source.n162 185
R315 source.n279 source.n278 185
R316 source.n277 source.n276 185
R317 source.n222 source.n221 185
R318 source.n271 source.n270 185
R319 source.n269 source.n268 185
R320 source.n226 source.n225 185
R321 source.n263 source.n262 185
R322 source.n261 source.n228 185
R323 source.n260 source.n259 185
R324 source.n231 source.n229 185
R325 source.n254 source.n253 185
R326 source.n252 source.n251 185
R327 source.n235 source.n234 185
R328 source.n246 source.n245 185
R329 source.n244 source.n243 185
R330 source.n239 source.n238 185
R331 source.n523 source.t46 149.524
R332 source.n447 source.t45 149.524
R333 source.n381 source.t18 149.524
R334 source.n305 source.t7 149.524
R335 source.n22 source.t22 149.524
R336 source.n98 source.t0 149.524
R337 source.n164 source.t34 149.524
R338 source.n240 source.t33 149.524
R339 source.n527 source.n521 104.615
R340 source.n528 source.n527 104.615
R341 source.n528 source.n517 104.615
R342 source.n535 source.n517 104.615
R343 source.n536 source.n535 104.615
R344 source.n536 source.n513 104.615
R345 source.n544 source.n513 104.615
R346 source.n545 source.n544 104.615
R347 source.n546 source.n545 104.615
R348 source.n546 source.n509 104.615
R349 source.n553 source.n509 104.615
R350 source.n554 source.n553 104.615
R351 source.n554 source.n505 104.615
R352 source.n561 source.n505 104.615
R353 source.n562 source.n561 104.615
R354 source.n451 source.n445 104.615
R355 source.n452 source.n451 104.615
R356 source.n452 source.n441 104.615
R357 source.n459 source.n441 104.615
R358 source.n460 source.n459 104.615
R359 source.n460 source.n437 104.615
R360 source.n468 source.n437 104.615
R361 source.n469 source.n468 104.615
R362 source.n470 source.n469 104.615
R363 source.n470 source.n433 104.615
R364 source.n477 source.n433 104.615
R365 source.n478 source.n477 104.615
R366 source.n478 source.n429 104.615
R367 source.n485 source.n429 104.615
R368 source.n486 source.n485 104.615
R369 source.n385 source.n379 104.615
R370 source.n386 source.n385 104.615
R371 source.n386 source.n375 104.615
R372 source.n393 source.n375 104.615
R373 source.n394 source.n393 104.615
R374 source.n394 source.n371 104.615
R375 source.n402 source.n371 104.615
R376 source.n403 source.n402 104.615
R377 source.n404 source.n403 104.615
R378 source.n404 source.n367 104.615
R379 source.n411 source.n367 104.615
R380 source.n412 source.n411 104.615
R381 source.n412 source.n363 104.615
R382 source.n419 source.n363 104.615
R383 source.n420 source.n419 104.615
R384 source.n309 source.n303 104.615
R385 source.n310 source.n309 104.615
R386 source.n310 source.n299 104.615
R387 source.n317 source.n299 104.615
R388 source.n318 source.n317 104.615
R389 source.n318 source.n295 104.615
R390 source.n326 source.n295 104.615
R391 source.n327 source.n326 104.615
R392 source.n328 source.n327 104.615
R393 source.n328 source.n291 104.615
R394 source.n335 source.n291 104.615
R395 source.n336 source.n335 104.615
R396 source.n336 source.n287 104.615
R397 source.n343 source.n287 104.615
R398 source.n344 source.n343 104.615
R399 source.n60 source.n59 104.615
R400 source.n59 source.n3 104.615
R401 source.n52 source.n3 104.615
R402 source.n52 source.n51 104.615
R403 source.n51 source.n7 104.615
R404 source.n44 source.n7 104.615
R405 source.n44 source.n43 104.615
R406 source.n43 source.n42 104.615
R407 source.n42 source.n11 104.615
R408 source.n35 source.n11 104.615
R409 source.n35 source.n34 104.615
R410 source.n34 source.n16 104.615
R411 source.n27 source.n16 104.615
R412 source.n27 source.n26 104.615
R413 source.n26 source.n20 104.615
R414 source.n136 source.n135 104.615
R415 source.n135 source.n79 104.615
R416 source.n128 source.n79 104.615
R417 source.n128 source.n127 104.615
R418 source.n127 source.n83 104.615
R419 source.n120 source.n83 104.615
R420 source.n120 source.n119 104.615
R421 source.n119 source.n118 104.615
R422 source.n118 source.n87 104.615
R423 source.n111 source.n87 104.615
R424 source.n111 source.n110 104.615
R425 source.n110 source.n92 104.615
R426 source.n103 source.n92 104.615
R427 source.n103 source.n102 104.615
R428 source.n102 source.n96 104.615
R429 source.n202 source.n201 104.615
R430 source.n201 source.n145 104.615
R431 source.n194 source.n145 104.615
R432 source.n194 source.n193 104.615
R433 source.n193 source.n149 104.615
R434 source.n186 source.n149 104.615
R435 source.n186 source.n185 104.615
R436 source.n185 source.n184 104.615
R437 source.n184 source.n153 104.615
R438 source.n177 source.n153 104.615
R439 source.n177 source.n176 104.615
R440 source.n176 source.n158 104.615
R441 source.n169 source.n158 104.615
R442 source.n169 source.n168 104.615
R443 source.n168 source.n162 104.615
R444 source.n278 source.n277 104.615
R445 source.n277 source.n221 104.615
R446 source.n270 source.n221 104.615
R447 source.n270 source.n269 104.615
R448 source.n269 source.n225 104.615
R449 source.n262 source.n225 104.615
R450 source.n262 source.n261 104.615
R451 source.n261 source.n260 104.615
R452 source.n260 source.n229 104.615
R453 source.n253 source.n229 104.615
R454 source.n253 source.n252 104.615
R455 source.n252 source.n234 104.615
R456 source.n245 source.n234 104.615
R457 source.n245 source.n244 104.615
R458 source.n244 source.n238 104.615
R459 source.t46 source.n521 52.3082
R460 source.t45 source.n445 52.3082
R461 source.t18 source.n379 52.3082
R462 source.t7 source.n303 52.3082
R463 source.t22 source.n20 52.3082
R464 source.t0 source.n96 52.3082
R465 source.t34 source.n162 52.3082
R466 source.t33 source.n238 52.3082
R467 source.n67 source.n66 42.8739
R468 source.n69 source.n68 42.8739
R469 source.n71 source.n70 42.8739
R470 source.n73 source.n72 42.8739
R471 source.n75 source.n74 42.8739
R472 source.n209 source.n208 42.8739
R473 source.n211 source.n210 42.8739
R474 source.n213 source.n212 42.8739
R475 source.n215 source.n214 42.8739
R476 source.n217 source.n216 42.8739
R477 source.n501 source.n500 42.8737
R478 source.n499 source.n498 42.8737
R479 source.n497 source.n496 42.8737
R480 source.n495 source.n494 42.8737
R481 source.n493 source.n492 42.8737
R482 source.n359 source.n358 42.8737
R483 source.n357 source.n356 42.8737
R484 source.n355 source.n354 42.8737
R485 source.n353 source.n352 42.8737
R486 source.n351 source.n350 42.8737
R487 source.n567 source.n566 29.8581
R488 source.n491 source.n490 29.8581
R489 source.n425 source.n424 29.8581
R490 source.n349 source.n348 29.8581
R491 source.n65 source.n64 29.8581
R492 source.n141 source.n140 29.8581
R493 source.n207 source.n206 29.8581
R494 source.n283 source.n282 29.8581
R495 source.n349 source.n283 22.1757
R496 source.n568 source.n65 16.4688
R497 source.n547 source.n512 13.1884
R498 source.n471 source.n436 13.1884
R499 source.n405 source.n370 13.1884
R500 source.n329 source.n294 13.1884
R501 source.n45 source.n10 13.1884
R502 source.n121 source.n86 13.1884
R503 source.n187 source.n152 13.1884
R504 source.n263 source.n228 13.1884
R505 source.n543 source.n542 12.8005
R506 source.n548 source.n510 12.8005
R507 source.n467 source.n466 12.8005
R508 source.n472 source.n434 12.8005
R509 source.n401 source.n400 12.8005
R510 source.n406 source.n368 12.8005
R511 source.n325 source.n324 12.8005
R512 source.n330 source.n292 12.8005
R513 source.n46 source.n8 12.8005
R514 source.n41 source.n12 12.8005
R515 source.n122 source.n84 12.8005
R516 source.n117 source.n88 12.8005
R517 source.n188 source.n150 12.8005
R518 source.n183 source.n154 12.8005
R519 source.n264 source.n226 12.8005
R520 source.n259 source.n230 12.8005
R521 source.n541 source.n514 12.0247
R522 source.n552 source.n551 12.0247
R523 source.n465 source.n438 12.0247
R524 source.n476 source.n475 12.0247
R525 source.n399 source.n372 12.0247
R526 source.n410 source.n409 12.0247
R527 source.n323 source.n296 12.0247
R528 source.n334 source.n333 12.0247
R529 source.n50 source.n49 12.0247
R530 source.n40 source.n13 12.0247
R531 source.n126 source.n125 12.0247
R532 source.n116 source.n89 12.0247
R533 source.n192 source.n191 12.0247
R534 source.n182 source.n155 12.0247
R535 source.n268 source.n267 12.0247
R536 source.n258 source.n231 12.0247
R537 source.n538 source.n537 11.249
R538 source.n555 source.n508 11.249
R539 source.n462 source.n461 11.249
R540 source.n479 source.n432 11.249
R541 source.n396 source.n395 11.249
R542 source.n413 source.n366 11.249
R543 source.n320 source.n319 11.249
R544 source.n337 source.n290 11.249
R545 source.n53 source.n6 11.249
R546 source.n37 source.n36 11.249
R547 source.n129 source.n82 11.249
R548 source.n113 source.n112 11.249
R549 source.n195 source.n148 11.249
R550 source.n179 source.n178 11.249
R551 source.n271 source.n224 11.249
R552 source.n255 source.n254 11.249
R553 source.n534 source.n516 10.4732
R554 source.n556 source.n506 10.4732
R555 source.n458 source.n440 10.4732
R556 source.n480 source.n430 10.4732
R557 source.n392 source.n374 10.4732
R558 source.n414 source.n364 10.4732
R559 source.n316 source.n298 10.4732
R560 source.n338 source.n288 10.4732
R561 source.n54 source.n4 10.4732
R562 source.n33 source.n15 10.4732
R563 source.n130 source.n80 10.4732
R564 source.n109 source.n91 10.4732
R565 source.n196 source.n146 10.4732
R566 source.n175 source.n157 10.4732
R567 source.n272 source.n222 10.4732
R568 source.n251 source.n233 10.4732
R569 source.n523 source.n522 10.2747
R570 source.n447 source.n446 10.2747
R571 source.n381 source.n380 10.2747
R572 source.n305 source.n304 10.2747
R573 source.n22 source.n21 10.2747
R574 source.n98 source.n97 10.2747
R575 source.n164 source.n163 10.2747
R576 source.n240 source.n239 10.2747
R577 source.n533 source.n518 9.69747
R578 source.n560 source.n559 9.69747
R579 source.n457 source.n442 9.69747
R580 source.n484 source.n483 9.69747
R581 source.n391 source.n376 9.69747
R582 source.n418 source.n417 9.69747
R583 source.n315 source.n300 9.69747
R584 source.n342 source.n341 9.69747
R585 source.n58 source.n57 9.69747
R586 source.n32 source.n17 9.69747
R587 source.n134 source.n133 9.69747
R588 source.n108 source.n93 9.69747
R589 source.n200 source.n199 9.69747
R590 source.n174 source.n159 9.69747
R591 source.n276 source.n275 9.69747
R592 source.n250 source.n235 9.69747
R593 source.n566 source.n565 9.45567
R594 source.n490 source.n489 9.45567
R595 source.n424 source.n423 9.45567
R596 source.n348 source.n347 9.45567
R597 source.n64 source.n63 9.45567
R598 source.n140 source.n139 9.45567
R599 source.n206 source.n205 9.45567
R600 source.n282 source.n281 9.45567
R601 source.n565 source.n564 9.3005
R602 source.n504 source.n503 9.3005
R603 source.n559 source.n558 9.3005
R604 source.n557 source.n556 9.3005
R605 source.n508 source.n507 9.3005
R606 source.n551 source.n550 9.3005
R607 source.n549 source.n548 9.3005
R608 source.n525 source.n524 9.3005
R609 source.n520 source.n519 9.3005
R610 source.n531 source.n530 9.3005
R611 source.n533 source.n532 9.3005
R612 source.n516 source.n515 9.3005
R613 source.n539 source.n538 9.3005
R614 source.n541 source.n540 9.3005
R615 source.n542 source.n511 9.3005
R616 source.n489 source.n488 9.3005
R617 source.n428 source.n427 9.3005
R618 source.n483 source.n482 9.3005
R619 source.n481 source.n480 9.3005
R620 source.n432 source.n431 9.3005
R621 source.n475 source.n474 9.3005
R622 source.n473 source.n472 9.3005
R623 source.n449 source.n448 9.3005
R624 source.n444 source.n443 9.3005
R625 source.n455 source.n454 9.3005
R626 source.n457 source.n456 9.3005
R627 source.n440 source.n439 9.3005
R628 source.n463 source.n462 9.3005
R629 source.n465 source.n464 9.3005
R630 source.n466 source.n435 9.3005
R631 source.n423 source.n422 9.3005
R632 source.n362 source.n361 9.3005
R633 source.n417 source.n416 9.3005
R634 source.n415 source.n414 9.3005
R635 source.n366 source.n365 9.3005
R636 source.n409 source.n408 9.3005
R637 source.n407 source.n406 9.3005
R638 source.n383 source.n382 9.3005
R639 source.n378 source.n377 9.3005
R640 source.n389 source.n388 9.3005
R641 source.n391 source.n390 9.3005
R642 source.n374 source.n373 9.3005
R643 source.n397 source.n396 9.3005
R644 source.n399 source.n398 9.3005
R645 source.n400 source.n369 9.3005
R646 source.n347 source.n346 9.3005
R647 source.n286 source.n285 9.3005
R648 source.n341 source.n340 9.3005
R649 source.n339 source.n338 9.3005
R650 source.n290 source.n289 9.3005
R651 source.n333 source.n332 9.3005
R652 source.n331 source.n330 9.3005
R653 source.n307 source.n306 9.3005
R654 source.n302 source.n301 9.3005
R655 source.n313 source.n312 9.3005
R656 source.n315 source.n314 9.3005
R657 source.n298 source.n297 9.3005
R658 source.n321 source.n320 9.3005
R659 source.n323 source.n322 9.3005
R660 source.n324 source.n293 9.3005
R661 source.n24 source.n23 9.3005
R662 source.n19 source.n18 9.3005
R663 source.n30 source.n29 9.3005
R664 source.n32 source.n31 9.3005
R665 source.n15 source.n14 9.3005
R666 source.n38 source.n37 9.3005
R667 source.n40 source.n39 9.3005
R668 source.n12 source.n9 9.3005
R669 source.n63 source.n62 9.3005
R670 source.n2 source.n1 9.3005
R671 source.n57 source.n56 9.3005
R672 source.n55 source.n54 9.3005
R673 source.n6 source.n5 9.3005
R674 source.n49 source.n48 9.3005
R675 source.n47 source.n46 9.3005
R676 source.n100 source.n99 9.3005
R677 source.n95 source.n94 9.3005
R678 source.n106 source.n105 9.3005
R679 source.n108 source.n107 9.3005
R680 source.n91 source.n90 9.3005
R681 source.n114 source.n113 9.3005
R682 source.n116 source.n115 9.3005
R683 source.n88 source.n85 9.3005
R684 source.n139 source.n138 9.3005
R685 source.n78 source.n77 9.3005
R686 source.n133 source.n132 9.3005
R687 source.n131 source.n130 9.3005
R688 source.n82 source.n81 9.3005
R689 source.n125 source.n124 9.3005
R690 source.n123 source.n122 9.3005
R691 source.n166 source.n165 9.3005
R692 source.n161 source.n160 9.3005
R693 source.n172 source.n171 9.3005
R694 source.n174 source.n173 9.3005
R695 source.n157 source.n156 9.3005
R696 source.n180 source.n179 9.3005
R697 source.n182 source.n181 9.3005
R698 source.n154 source.n151 9.3005
R699 source.n205 source.n204 9.3005
R700 source.n144 source.n143 9.3005
R701 source.n199 source.n198 9.3005
R702 source.n197 source.n196 9.3005
R703 source.n148 source.n147 9.3005
R704 source.n191 source.n190 9.3005
R705 source.n189 source.n188 9.3005
R706 source.n242 source.n241 9.3005
R707 source.n237 source.n236 9.3005
R708 source.n248 source.n247 9.3005
R709 source.n250 source.n249 9.3005
R710 source.n233 source.n232 9.3005
R711 source.n256 source.n255 9.3005
R712 source.n258 source.n257 9.3005
R713 source.n230 source.n227 9.3005
R714 source.n281 source.n280 9.3005
R715 source.n220 source.n219 9.3005
R716 source.n275 source.n274 9.3005
R717 source.n273 source.n272 9.3005
R718 source.n224 source.n223 9.3005
R719 source.n267 source.n266 9.3005
R720 source.n265 source.n264 9.3005
R721 source.n530 source.n529 8.92171
R722 source.n563 source.n504 8.92171
R723 source.n454 source.n453 8.92171
R724 source.n487 source.n428 8.92171
R725 source.n388 source.n387 8.92171
R726 source.n421 source.n362 8.92171
R727 source.n312 source.n311 8.92171
R728 source.n345 source.n286 8.92171
R729 source.n61 source.n2 8.92171
R730 source.n29 source.n28 8.92171
R731 source.n137 source.n78 8.92171
R732 source.n105 source.n104 8.92171
R733 source.n203 source.n144 8.92171
R734 source.n171 source.n170 8.92171
R735 source.n279 source.n220 8.92171
R736 source.n247 source.n246 8.92171
R737 source.n526 source.n520 8.14595
R738 source.n564 source.n502 8.14595
R739 source.n450 source.n444 8.14595
R740 source.n488 source.n426 8.14595
R741 source.n384 source.n378 8.14595
R742 source.n422 source.n360 8.14595
R743 source.n308 source.n302 8.14595
R744 source.n346 source.n284 8.14595
R745 source.n62 source.n0 8.14595
R746 source.n25 source.n19 8.14595
R747 source.n138 source.n76 8.14595
R748 source.n101 source.n95 8.14595
R749 source.n204 source.n142 8.14595
R750 source.n167 source.n161 8.14595
R751 source.n280 source.n218 8.14595
R752 source.n243 source.n237 8.14595
R753 source.n525 source.n522 7.3702
R754 source.n449 source.n446 7.3702
R755 source.n383 source.n380 7.3702
R756 source.n307 source.n304 7.3702
R757 source.n24 source.n21 7.3702
R758 source.n100 source.n97 7.3702
R759 source.n166 source.n163 7.3702
R760 source.n242 source.n239 7.3702
R761 source.n526 source.n525 5.81868
R762 source.n566 source.n502 5.81868
R763 source.n450 source.n449 5.81868
R764 source.n490 source.n426 5.81868
R765 source.n384 source.n383 5.81868
R766 source.n424 source.n360 5.81868
R767 source.n308 source.n307 5.81868
R768 source.n348 source.n284 5.81868
R769 source.n64 source.n0 5.81868
R770 source.n25 source.n24 5.81868
R771 source.n140 source.n76 5.81868
R772 source.n101 source.n100 5.81868
R773 source.n206 source.n142 5.81868
R774 source.n167 source.n166 5.81868
R775 source.n282 source.n218 5.81868
R776 source.n243 source.n242 5.81868
R777 source.n568 source.n567 5.7074
R778 source.n529 source.n520 5.04292
R779 source.n564 source.n563 5.04292
R780 source.n453 source.n444 5.04292
R781 source.n488 source.n487 5.04292
R782 source.n387 source.n378 5.04292
R783 source.n422 source.n421 5.04292
R784 source.n311 source.n302 5.04292
R785 source.n346 source.n345 5.04292
R786 source.n62 source.n61 5.04292
R787 source.n28 source.n19 5.04292
R788 source.n138 source.n137 5.04292
R789 source.n104 source.n95 5.04292
R790 source.n204 source.n203 5.04292
R791 source.n170 source.n161 5.04292
R792 source.n280 source.n279 5.04292
R793 source.n246 source.n237 5.04292
R794 source.n530 source.n518 4.26717
R795 source.n560 source.n504 4.26717
R796 source.n454 source.n442 4.26717
R797 source.n484 source.n428 4.26717
R798 source.n388 source.n376 4.26717
R799 source.n418 source.n362 4.26717
R800 source.n312 source.n300 4.26717
R801 source.n342 source.n286 4.26717
R802 source.n58 source.n2 4.26717
R803 source.n29 source.n17 4.26717
R804 source.n134 source.n78 4.26717
R805 source.n105 source.n93 4.26717
R806 source.n200 source.n144 4.26717
R807 source.n171 source.n159 4.26717
R808 source.n276 source.n220 4.26717
R809 source.n247 source.n235 4.26717
R810 source.n534 source.n533 3.49141
R811 source.n559 source.n506 3.49141
R812 source.n458 source.n457 3.49141
R813 source.n483 source.n430 3.49141
R814 source.n392 source.n391 3.49141
R815 source.n417 source.n364 3.49141
R816 source.n316 source.n315 3.49141
R817 source.n341 source.n288 3.49141
R818 source.n57 source.n4 3.49141
R819 source.n33 source.n32 3.49141
R820 source.n133 source.n80 3.49141
R821 source.n109 source.n108 3.49141
R822 source.n199 source.n146 3.49141
R823 source.n175 source.n174 3.49141
R824 source.n275 source.n222 3.49141
R825 source.n251 source.n250 3.49141
R826 source.n524 source.n523 2.84303
R827 source.n448 source.n447 2.84303
R828 source.n382 source.n381 2.84303
R829 source.n306 source.n305 2.84303
R830 source.n23 source.n22 2.84303
R831 source.n99 source.n98 2.84303
R832 source.n165 source.n164 2.84303
R833 source.n241 source.n240 2.84303
R834 source.n537 source.n516 2.71565
R835 source.n556 source.n555 2.71565
R836 source.n461 source.n440 2.71565
R837 source.n480 source.n479 2.71565
R838 source.n395 source.n374 2.71565
R839 source.n414 source.n413 2.71565
R840 source.n319 source.n298 2.71565
R841 source.n338 source.n337 2.71565
R842 source.n54 source.n53 2.71565
R843 source.n36 source.n15 2.71565
R844 source.n130 source.n129 2.71565
R845 source.n112 source.n91 2.71565
R846 source.n196 source.n195 2.71565
R847 source.n178 source.n157 2.71565
R848 source.n272 source.n271 2.71565
R849 source.n254 source.n233 2.71565
R850 source.n538 source.n514 1.93989
R851 source.n552 source.n508 1.93989
R852 source.n462 source.n438 1.93989
R853 source.n476 source.n432 1.93989
R854 source.n396 source.n372 1.93989
R855 source.n410 source.n366 1.93989
R856 source.n320 source.n296 1.93989
R857 source.n334 source.n290 1.93989
R858 source.n50 source.n6 1.93989
R859 source.n37 source.n13 1.93989
R860 source.n126 source.n82 1.93989
R861 source.n113 source.n89 1.93989
R862 source.n192 source.n148 1.93989
R863 source.n179 source.n155 1.93989
R864 source.n268 source.n224 1.93989
R865 source.n255 source.n231 1.93989
R866 source.n500 source.t41 1.6505
R867 source.n500 source.t47 1.6505
R868 source.n498 source.t35 1.6505
R869 source.n498 source.t36 1.6505
R870 source.n496 source.t31 1.6505
R871 source.n496 source.t30 1.6505
R872 source.n494 source.t27 1.6505
R873 source.n494 source.t24 1.6505
R874 source.n492 source.t43 1.6505
R875 source.n492 source.t28 1.6505
R876 source.n358 source.t4 1.6505
R877 source.n358 source.t3 1.6505
R878 source.n356 source.t1 1.6505
R879 source.n356 source.t20 1.6505
R880 source.n354 source.t23 1.6505
R881 source.n354 source.t10 1.6505
R882 source.n352 source.t2 1.6505
R883 source.n352 source.t21 1.6505
R884 source.n350 source.t19 1.6505
R885 source.n350 source.t8 1.6505
R886 source.n66 source.t13 1.6505
R887 source.n66 source.t9 1.6505
R888 source.n68 source.t14 1.6505
R889 source.n68 source.t6 1.6505
R890 source.n70 source.t15 1.6505
R891 source.n70 source.t12 1.6505
R892 source.n72 source.t16 1.6505
R893 source.n72 source.t17 1.6505
R894 source.n74 source.t5 1.6505
R895 source.n74 source.t11 1.6505
R896 source.n208 source.t37 1.6505
R897 source.n208 source.t44 1.6505
R898 source.n210 source.t38 1.6505
R899 source.n210 source.t26 1.6505
R900 source.n212 source.t39 1.6505
R901 source.n212 source.t25 1.6505
R902 source.n214 source.t40 1.6505
R903 source.n214 source.t29 1.6505
R904 source.n216 source.t42 1.6505
R905 source.n216 source.t32 1.6505
R906 source.n543 source.n541 1.16414
R907 source.n551 source.n510 1.16414
R908 source.n467 source.n465 1.16414
R909 source.n475 source.n434 1.16414
R910 source.n401 source.n399 1.16414
R911 source.n409 source.n368 1.16414
R912 source.n325 source.n323 1.16414
R913 source.n333 source.n292 1.16414
R914 source.n49 source.n8 1.16414
R915 source.n41 source.n40 1.16414
R916 source.n125 source.n84 1.16414
R917 source.n117 source.n116 1.16414
R918 source.n191 source.n150 1.16414
R919 source.n183 source.n182 1.16414
R920 source.n267 source.n226 1.16414
R921 source.n259 source.n258 1.16414
R922 source.n283 source.n217 0.888431
R923 source.n217 source.n215 0.888431
R924 source.n215 source.n213 0.888431
R925 source.n213 source.n211 0.888431
R926 source.n211 source.n209 0.888431
R927 source.n209 source.n207 0.888431
R928 source.n141 source.n75 0.888431
R929 source.n75 source.n73 0.888431
R930 source.n73 source.n71 0.888431
R931 source.n71 source.n69 0.888431
R932 source.n69 source.n67 0.888431
R933 source.n67 source.n65 0.888431
R934 source.n351 source.n349 0.888431
R935 source.n353 source.n351 0.888431
R936 source.n355 source.n353 0.888431
R937 source.n357 source.n355 0.888431
R938 source.n359 source.n357 0.888431
R939 source.n425 source.n359 0.888431
R940 source.n493 source.n491 0.888431
R941 source.n495 source.n493 0.888431
R942 source.n497 source.n495 0.888431
R943 source.n499 source.n497 0.888431
R944 source.n501 source.n499 0.888431
R945 source.n567 source.n501 0.888431
R946 source.n207 source.n141 0.470328
R947 source.n491 source.n425 0.470328
R948 source.n542 source.n512 0.388379
R949 source.n548 source.n547 0.388379
R950 source.n466 source.n436 0.388379
R951 source.n472 source.n471 0.388379
R952 source.n400 source.n370 0.388379
R953 source.n406 source.n405 0.388379
R954 source.n324 source.n294 0.388379
R955 source.n330 source.n329 0.388379
R956 source.n46 source.n45 0.388379
R957 source.n12 source.n10 0.388379
R958 source.n122 source.n121 0.388379
R959 source.n88 source.n86 0.388379
R960 source.n188 source.n187 0.388379
R961 source.n154 source.n152 0.388379
R962 source.n264 source.n263 0.388379
R963 source.n230 source.n228 0.388379
R964 source source.n568 0.188
R965 source.n524 source.n519 0.155672
R966 source.n531 source.n519 0.155672
R967 source.n532 source.n531 0.155672
R968 source.n532 source.n515 0.155672
R969 source.n539 source.n515 0.155672
R970 source.n540 source.n539 0.155672
R971 source.n540 source.n511 0.155672
R972 source.n549 source.n511 0.155672
R973 source.n550 source.n549 0.155672
R974 source.n550 source.n507 0.155672
R975 source.n557 source.n507 0.155672
R976 source.n558 source.n557 0.155672
R977 source.n558 source.n503 0.155672
R978 source.n565 source.n503 0.155672
R979 source.n448 source.n443 0.155672
R980 source.n455 source.n443 0.155672
R981 source.n456 source.n455 0.155672
R982 source.n456 source.n439 0.155672
R983 source.n463 source.n439 0.155672
R984 source.n464 source.n463 0.155672
R985 source.n464 source.n435 0.155672
R986 source.n473 source.n435 0.155672
R987 source.n474 source.n473 0.155672
R988 source.n474 source.n431 0.155672
R989 source.n481 source.n431 0.155672
R990 source.n482 source.n481 0.155672
R991 source.n482 source.n427 0.155672
R992 source.n489 source.n427 0.155672
R993 source.n382 source.n377 0.155672
R994 source.n389 source.n377 0.155672
R995 source.n390 source.n389 0.155672
R996 source.n390 source.n373 0.155672
R997 source.n397 source.n373 0.155672
R998 source.n398 source.n397 0.155672
R999 source.n398 source.n369 0.155672
R1000 source.n407 source.n369 0.155672
R1001 source.n408 source.n407 0.155672
R1002 source.n408 source.n365 0.155672
R1003 source.n415 source.n365 0.155672
R1004 source.n416 source.n415 0.155672
R1005 source.n416 source.n361 0.155672
R1006 source.n423 source.n361 0.155672
R1007 source.n306 source.n301 0.155672
R1008 source.n313 source.n301 0.155672
R1009 source.n314 source.n313 0.155672
R1010 source.n314 source.n297 0.155672
R1011 source.n321 source.n297 0.155672
R1012 source.n322 source.n321 0.155672
R1013 source.n322 source.n293 0.155672
R1014 source.n331 source.n293 0.155672
R1015 source.n332 source.n331 0.155672
R1016 source.n332 source.n289 0.155672
R1017 source.n339 source.n289 0.155672
R1018 source.n340 source.n339 0.155672
R1019 source.n340 source.n285 0.155672
R1020 source.n347 source.n285 0.155672
R1021 source.n63 source.n1 0.155672
R1022 source.n56 source.n1 0.155672
R1023 source.n56 source.n55 0.155672
R1024 source.n55 source.n5 0.155672
R1025 source.n48 source.n5 0.155672
R1026 source.n48 source.n47 0.155672
R1027 source.n47 source.n9 0.155672
R1028 source.n39 source.n9 0.155672
R1029 source.n39 source.n38 0.155672
R1030 source.n38 source.n14 0.155672
R1031 source.n31 source.n14 0.155672
R1032 source.n31 source.n30 0.155672
R1033 source.n30 source.n18 0.155672
R1034 source.n23 source.n18 0.155672
R1035 source.n139 source.n77 0.155672
R1036 source.n132 source.n77 0.155672
R1037 source.n132 source.n131 0.155672
R1038 source.n131 source.n81 0.155672
R1039 source.n124 source.n81 0.155672
R1040 source.n124 source.n123 0.155672
R1041 source.n123 source.n85 0.155672
R1042 source.n115 source.n85 0.155672
R1043 source.n115 source.n114 0.155672
R1044 source.n114 source.n90 0.155672
R1045 source.n107 source.n90 0.155672
R1046 source.n107 source.n106 0.155672
R1047 source.n106 source.n94 0.155672
R1048 source.n99 source.n94 0.155672
R1049 source.n205 source.n143 0.155672
R1050 source.n198 source.n143 0.155672
R1051 source.n198 source.n197 0.155672
R1052 source.n197 source.n147 0.155672
R1053 source.n190 source.n147 0.155672
R1054 source.n190 source.n189 0.155672
R1055 source.n189 source.n151 0.155672
R1056 source.n181 source.n151 0.155672
R1057 source.n181 source.n180 0.155672
R1058 source.n180 source.n156 0.155672
R1059 source.n173 source.n156 0.155672
R1060 source.n173 source.n172 0.155672
R1061 source.n172 source.n160 0.155672
R1062 source.n165 source.n160 0.155672
R1063 source.n281 source.n219 0.155672
R1064 source.n274 source.n219 0.155672
R1065 source.n274 source.n273 0.155672
R1066 source.n273 source.n223 0.155672
R1067 source.n266 source.n223 0.155672
R1068 source.n266 source.n265 0.155672
R1069 source.n265 source.n227 0.155672
R1070 source.n257 source.n227 0.155672
R1071 source.n257 source.n256 0.155672
R1072 source.n256 source.n232 0.155672
R1073 source.n249 source.n232 0.155672
R1074 source.n249 source.n248 0.155672
R1075 source.n248 source.n236 0.155672
R1076 source.n241 source.n236 0.155672
R1077 plus.n11 plus.t7 495.62
R1078 plus.n53 plus.t21 495.62
R1079 plus.n40 plus.t2 469.262
R1080 plus.n38 plus.t12 469.262
R1081 plus.n2 plus.t5 469.262
R1082 plus.n32 plus.t23 469.262
R1083 plus.n4 plus.t10 469.262
R1084 plus.n26 plus.t3 469.262
R1085 plus.n6 plus.t13 469.262
R1086 plus.n20 plus.t6 469.262
R1087 plus.n8 plus.t11 469.262
R1088 plus.n14 plus.t4 469.262
R1089 plus.n10 plus.t18 469.262
R1090 plus.n82 plus.t17 469.262
R1091 plus.n80 plus.t16 469.262
R1092 plus.n44 plus.t15 469.262
R1093 plus.n74 plus.t14 469.262
R1094 plus.n46 plus.t20 469.262
R1095 plus.n68 plus.t1 469.262
R1096 plus.n48 plus.t0 469.262
R1097 plus.n62 plus.t9 469.262
R1098 plus.n50 plus.t8 469.262
R1099 plus.n56 plus.t19 469.262
R1100 plus.n52 plus.t22 469.262
R1101 plus.n13 plus.n12 161.3
R1102 plus.n14 plus.n9 161.3
R1103 plus.n16 plus.n15 161.3
R1104 plus.n17 plus.n8 161.3
R1105 plus.n19 plus.n18 161.3
R1106 plus.n20 plus.n7 161.3
R1107 plus.n22 plus.n21 161.3
R1108 plus.n23 plus.n6 161.3
R1109 plus.n25 plus.n24 161.3
R1110 plus.n26 plus.n5 161.3
R1111 plus.n28 plus.n27 161.3
R1112 plus.n29 plus.n4 161.3
R1113 plus.n31 plus.n30 161.3
R1114 plus.n32 plus.n3 161.3
R1115 plus.n34 plus.n33 161.3
R1116 plus.n35 plus.n2 161.3
R1117 plus.n37 plus.n36 161.3
R1118 plus.n38 plus.n1 161.3
R1119 plus.n39 plus.n0 161.3
R1120 plus.n41 plus.n40 161.3
R1121 plus.n55 plus.n54 161.3
R1122 plus.n56 plus.n51 161.3
R1123 plus.n58 plus.n57 161.3
R1124 plus.n59 plus.n50 161.3
R1125 plus.n61 plus.n60 161.3
R1126 plus.n62 plus.n49 161.3
R1127 plus.n64 plus.n63 161.3
R1128 plus.n65 plus.n48 161.3
R1129 plus.n67 plus.n66 161.3
R1130 plus.n68 plus.n47 161.3
R1131 plus.n70 plus.n69 161.3
R1132 plus.n71 plus.n46 161.3
R1133 plus.n73 plus.n72 161.3
R1134 plus.n74 plus.n45 161.3
R1135 plus.n76 plus.n75 161.3
R1136 plus.n77 plus.n44 161.3
R1137 plus.n79 plus.n78 161.3
R1138 plus.n80 plus.n43 161.3
R1139 plus.n81 plus.n42 161.3
R1140 plus.n83 plus.n82 161.3
R1141 plus.n40 plus.n39 46.0096
R1142 plus.n82 plus.n81 46.0096
R1143 plus.n12 plus.n11 45.0871
R1144 plus.n54 plus.n53 45.0871
R1145 plus.n38 plus.n37 41.6278
R1146 plus.n13 plus.n10 41.6278
R1147 plus.n80 plus.n79 41.6278
R1148 plus.n55 plus.n52 41.6278
R1149 plus.n33 plus.n2 37.246
R1150 plus.n15 plus.n14 37.246
R1151 plus.n75 plus.n44 37.246
R1152 plus.n57 plus.n56 37.246
R1153 plus plus.n83 36.0369
R1154 plus.n32 plus.n31 32.8641
R1155 plus.n19 plus.n8 32.8641
R1156 plus.n74 plus.n73 32.8641
R1157 plus.n61 plus.n50 32.8641
R1158 plus.n27 plus.n4 28.4823
R1159 plus.n21 plus.n20 28.4823
R1160 plus.n69 plus.n46 28.4823
R1161 plus.n63 plus.n62 28.4823
R1162 plus.n25 plus.n6 24.1005
R1163 plus.n26 plus.n25 24.1005
R1164 plus.n68 plus.n67 24.1005
R1165 plus.n67 plus.n48 24.1005
R1166 plus.n27 plus.n26 19.7187
R1167 plus.n21 plus.n6 19.7187
R1168 plus.n69 plus.n68 19.7187
R1169 plus.n63 plus.n48 19.7187
R1170 plus.n31 plus.n4 15.3369
R1171 plus.n20 plus.n19 15.3369
R1172 plus.n73 plus.n46 15.3369
R1173 plus.n62 plus.n61 15.3369
R1174 plus.n11 plus.n10 14.1472
R1175 plus.n53 plus.n52 14.1472
R1176 plus plus.n41 12.3225
R1177 plus.n33 plus.n32 10.955
R1178 plus.n15 plus.n8 10.955
R1179 plus.n75 plus.n74 10.955
R1180 plus.n57 plus.n50 10.955
R1181 plus.n37 plus.n2 6.57323
R1182 plus.n14 plus.n13 6.57323
R1183 plus.n79 plus.n44 6.57323
R1184 plus.n56 plus.n55 6.57323
R1185 plus.n39 plus.n38 2.19141
R1186 plus.n81 plus.n80 2.19141
R1187 plus.n12 plus.n9 0.189894
R1188 plus.n16 plus.n9 0.189894
R1189 plus.n17 plus.n16 0.189894
R1190 plus.n18 plus.n17 0.189894
R1191 plus.n18 plus.n7 0.189894
R1192 plus.n22 plus.n7 0.189894
R1193 plus.n23 plus.n22 0.189894
R1194 plus.n24 plus.n23 0.189894
R1195 plus.n24 plus.n5 0.189894
R1196 plus.n28 plus.n5 0.189894
R1197 plus.n29 plus.n28 0.189894
R1198 plus.n30 plus.n29 0.189894
R1199 plus.n30 plus.n3 0.189894
R1200 plus.n34 plus.n3 0.189894
R1201 plus.n35 plus.n34 0.189894
R1202 plus.n36 plus.n35 0.189894
R1203 plus.n36 plus.n1 0.189894
R1204 plus.n1 plus.n0 0.189894
R1205 plus.n41 plus.n0 0.189894
R1206 plus.n83 plus.n42 0.189894
R1207 plus.n43 plus.n42 0.189894
R1208 plus.n78 plus.n43 0.189894
R1209 plus.n78 plus.n77 0.189894
R1210 plus.n77 plus.n76 0.189894
R1211 plus.n76 plus.n45 0.189894
R1212 plus.n72 plus.n45 0.189894
R1213 plus.n72 plus.n71 0.189894
R1214 plus.n71 plus.n70 0.189894
R1215 plus.n70 plus.n47 0.189894
R1216 plus.n66 plus.n47 0.189894
R1217 plus.n66 plus.n65 0.189894
R1218 plus.n65 plus.n64 0.189894
R1219 plus.n64 plus.n49 0.189894
R1220 plus.n60 plus.n49 0.189894
R1221 plus.n60 plus.n59 0.189894
R1222 plus.n59 plus.n58 0.189894
R1223 plus.n58 plus.n51 0.189894
R1224 plus.n54 plus.n51 0.189894
R1225 drain_left.n13 drain_left.n11 60.4406
R1226 drain_left.n7 drain_left.n5 60.4404
R1227 drain_left.n2 drain_left.n0 60.4404
R1228 drain_left.n19 drain_left.n18 59.5527
R1229 drain_left.n17 drain_left.n16 59.5527
R1230 drain_left.n15 drain_left.n14 59.5527
R1231 drain_left.n13 drain_left.n12 59.5527
R1232 drain_left.n7 drain_left.n6 59.5525
R1233 drain_left.n9 drain_left.n8 59.5525
R1234 drain_left.n4 drain_left.n3 59.5525
R1235 drain_left.n2 drain_left.n1 59.5525
R1236 drain_left.n21 drain_left.n20 59.5525
R1237 drain_left drain_left.n10 35.8024
R1238 drain_left drain_left.n21 6.54115
R1239 drain_left.n5 drain_left.t1 1.6505
R1240 drain_left.n5 drain_left.t2 1.6505
R1241 drain_left.n6 drain_left.t15 1.6505
R1242 drain_left.n6 drain_left.t4 1.6505
R1243 drain_left.n8 drain_left.t23 1.6505
R1244 drain_left.n8 drain_left.t14 1.6505
R1245 drain_left.n3 drain_left.t3 1.6505
R1246 drain_left.n3 drain_left.t22 1.6505
R1247 drain_left.n1 drain_left.t8 1.6505
R1248 drain_left.n1 drain_left.t9 1.6505
R1249 drain_left.n0 drain_left.t6 1.6505
R1250 drain_left.n0 drain_left.t7 1.6505
R1251 drain_left.n20 drain_left.t11 1.6505
R1252 drain_left.n20 drain_left.t21 1.6505
R1253 drain_left.n18 drain_left.t0 1.6505
R1254 drain_left.n18 drain_left.t18 1.6505
R1255 drain_left.n16 drain_left.t20 1.6505
R1256 drain_left.n16 drain_left.t13 1.6505
R1257 drain_left.n14 drain_left.t17 1.6505
R1258 drain_left.n14 drain_left.t10 1.6505
R1259 drain_left.n12 drain_left.t19 1.6505
R1260 drain_left.n12 drain_left.t12 1.6505
R1261 drain_left.n11 drain_left.t16 1.6505
R1262 drain_left.n11 drain_left.t5 1.6505
R1263 drain_left.n9 drain_left.n7 0.888431
R1264 drain_left.n4 drain_left.n2 0.888431
R1265 drain_left.n15 drain_left.n13 0.888431
R1266 drain_left.n17 drain_left.n15 0.888431
R1267 drain_left.n19 drain_left.n17 0.888431
R1268 drain_left.n21 drain_left.n19 0.888431
R1269 drain_left.n10 drain_left.n9 0.389119
R1270 drain_left.n10 drain_left.n4 0.389119
C0 minus plus 7.38089f
C1 minus drain_right 14.939599f
C2 plus drain_left 15.2801f
C3 minus source 15.2298f
C4 drain_right drain_left 1.87044f
C5 drain_right plus 0.498726f
C6 source drain_left 28.3559f
C7 source plus 15.243799f
C8 drain_right source 28.3584f
C9 minus drain_left 0.174517f
C10 drain_right a_n3394_n3288# 7.89082f
C11 drain_left a_n3394_n3288# 8.36606f
C12 source a_n3394_n3288# 9.585801f
C13 minus a_n3394_n3288# 13.745971f
C14 plus a_n3394_n3288# 15.63595f
C15 drain_left.t6 a_n3394_n3288# 0.259395f
C16 drain_left.t7 a_n3394_n3288# 0.259395f
C17 drain_left.n0 a_n3394_n3288# 2.31405f
C18 drain_left.t8 a_n3394_n3288# 0.259395f
C19 drain_left.t9 a_n3394_n3288# 0.259395f
C20 drain_left.n1 a_n3394_n3288# 2.30822f
C21 drain_left.n2 a_n3394_n3288# 0.777387f
C22 drain_left.t3 a_n3394_n3288# 0.259395f
C23 drain_left.t22 a_n3394_n3288# 0.259395f
C24 drain_left.n3 a_n3394_n3288# 2.30822f
C25 drain_left.n4 a_n3394_n3288# 0.343723f
C26 drain_left.t1 a_n3394_n3288# 0.259395f
C27 drain_left.t2 a_n3394_n3288# 0.259395f
C28 drain_left.n5 a_n3394_n3288# 2.31405f
C29 drain_left.t15 a_n3394_n3288# 0.259395f
C30 drain_left.t4 a_n3394_n3288# 0.259395f
C31 drain_left.n6 a_n3394_n3288# 2.30822f
C32 drain_left.n7 a_n3394_n3288# 0.777387f
C33 drain_left.t23 a_n3394_n3288# 0.259395f
C34 drain_left.t14 a_n3394_n3288# 0.259395f
C35 drain_left.n8 a_n3394_n3288# 2.30822f
C36 drain_left.n9 a_n3394_n3288# 0.343723f
C37 drain_left.n10 a_n3394_n3288# 1.80516f
C38 drain_left.t16 a_n3394_n3288# 0.259395f
C39 drain_left.t5 a_n3394_n3288# 0.259395f
C40 drain_left.n11 a_n3394_n3288# 2.31406f
C41 drain_left.t19 a_n3394_n3288# 0.259395f
C42 drain_left.t12 a_n3394_n3288# 0.259395f
C43 drain_left.n12 a_n3394_n3288# 2.30823f
C44 drain_left.n13 a_n3394_n3288# 0.777368f
C45 drain_left.t17 a_n3394_n3288# 0.259395f
C46 drain_left.t10 a_n3394_n3288# 0.259395f
C47 drain_left.n14 a_n3394_n3288# 2.30823f
C48 drain_left.n15 a_n3394_n3288# 0.386092f
C49 drain_left.t20 a_n3394_n3288# 0.259395f
C50 drain_left.t13 a_n3394_n3288# 0.259395f
C51 drain_left.n16 a_n3394_n3288# 2.30823f
C52 drain_left.n17 a_n3394_n3288# 0.386092f
C53 drain_left.t0 a_n3394_n3288# 0.259395f
C54 drain_left.t18 a_n3394_n3288# 0.259395f
C55 drain_left.n18 a_n3394_n3288# 2.30823f
C56 drain_left.n19 a_n3394_n3288# 0.386092f
C57 drain_left.t11 a_n3394_n3288# 0.259395f
C58 drain_left.t21 a_n3394_n3288# 0.259395f
C59 drain_left.n20 a_n3394_n3288# 2.30822f
C60 drain_left.n21 a_n3394_n3288# 0.628053f
C61 plus.n0 a_n3394_n3288# 0.039593f
C62 plus.t2 a_n3394_n3288# 0.948353f
C63 plus.t12 a_n3394_n3288# 0.948353f
C64 plus.n1 a_n3394_n3288# 0.039593f
C65 plus.t5 a_n3394_n3288# 0.948353f
C66 plus.n2 a_n3394_n3288# 0.378221f
C67 plus.n3 a_n3394_n3288# 0.039593f
C68 plus.t23 a_n3394_n3288# 0.948353f
C69 plus.t10 a_n3394_n3288# 0.948353f
C70 plus.n4 a_n3394_n3288# 0.378221f
C71 plus.n5 a_n3394_n3288# 0.039593f
C72 plus.t3 a_n3394_n3288# 0.948353f
C73 plus.t13 a_n3394_n3288# 0.948353f
C74 plus.n6 a_n3394_n3288# 0.378221f
C75 plus.n7 a_n3394_n3288# 0.039593f
C76 plus.t6 a_n3394_n3288# 0.948353f
C77 plus.t11 a_n3394_n3288# 0.948353f
C78 plus.n8 a_n3394_n3288# 0.378221f
C79 plus.n9 a_n3394_n3288# 0.039593f
C80 plus.t4 a_n3394_n3288# 0.948353f
C81 plus.t18 a_n3394_n3288# 0.948353f
C82 plus.n10 a_n3394_n3288# 0.386323f
C83 plus.t7 a_n3394_n3288# 0.968504f
C84 plus.n11 a_n3394_n3288# 0.360177f
C85 plus.n12 a_n3394_n3288# 0.170449f
C86 plus.n13 a_n3394_n3288# 0.008984f
C87 plus.n14 a_n3394_n3288# 0.378221f
C88 plus.n15 a_n3394_n3288# 0.008984f
C89 plus.n16 a_n3394_n3288# 0.039593f
C90 plus.n17 a_n3394_n3288# 0.039593f
C91 plus.n18 a_n3394_n3288# 0.039593f
C92 plus.n19 a_n3394_n3288# 0.008984f
C93 plus.n20 a_n3394_n3288# 0.378221f
C94 plus.n21 a_n3394_n3288# 0.008984f
C95 plus.n22 a_n3394_n3288# 0.039593f
C96 plus.n23 a_n3394_n3288# 0.039593f
C97 plus.n24 a_n3394_n3288# 0.039593f
C98 plus.n25 a_n3394_n3288# 0.008984f
C99 plus.n26 a_n3394_n3288# 0.378221f
C100 plus.n27 a_n3394_n3288# 0.008984f
C101 plus.n28 a_n3394_n3288# 0.039593f
C102 plus.n29 a_n3394_n3288# 0.039593f
C103 plus.n30 a_n3394_n3288# 0.039593f
C104 plus.n31 a_n3394_n3288# 0.008984f
C105 plus.n32 a_n3394_n3288# 0.378221f
C106 plus.n33 a_n3394_n3288# 0.008984f
C107 plus.n34 a_n3394_n3288# 0.039593f
C108 plus.n35 a_n3394_n3288# 0.039593f
C109 plus.n36 a_n3394_n3288# 0.039593f
C110 plus.n37 a_n3394_n3288# 0.008984f
C111 plus.n38 a_n3394_n3288# 0.378221f
C112 plus.n39 a_n3394_n3288# 0.008984f
C113 plus.n40 a_n3394_n3288# 0.378587f
C114 plus.n41 a_n3394_n3288# 0.459805f
C115 plus.n42 a_n3394_n3288# 0.039593f
C116 plus.t17 a_n3394_n3288# 0.948353f
C117 plus.n43 a_n3394_n3288# 0.039593f
C118 plus.t16 a_n3394_n3288# 0.948353f
C119 plus.t15 a_n3394_n3288# 0.948353f
C120 plus.n44 a_n3394_n3288# 0.378221f
C121 plus.n45 a_n3394_n3288# 0.039593f
C122 plus.t14 a_n3394_n3288# 0.948353f
C123 plus.t20 a_n3394_n3288# 0.948353f
C124 plus.n46 a_n3394_n3288# 0.378221f
C125 plus.n47 a_n3394_n3288# 0.039593f
C126 plus.t1 a_n3394_n3288# 0.948353f
C127 plus.t0 a_n3394_n3288# 0.948353f
C128 plus.n48 a_n3394_n3288# 0.378221f
C129 plus.n49 a_n3394_n3288# 0.039593f
C130 plus.t9 a_n3394_n3288# 0.948353f
C131 plus.t8 a_n3394_n3288# 0.948353f
C132 plus.n50 a_n3394_n3288# 0.378221f
C133 plus.n51 a_n3394_n3288# 0.039593f
C134 plus.t19 a_n3394_n3288# 0.948353f
C135 plus.t22 a_n3394_n3288# 0.948353f
C136 plus.n52 a_n3394_n3288# 0.386323f
C137 plus.t21 a_n3394_n3288# 0.968504f
C138 plus.n53 a_n3394_n3288# 0.360177f
C139 plus.n54 a_n3394_n3288# 0.170449f
C140 plus.n55 a_n3394_n3288# 0.008984f
C141 plus.n56 a_n3394_n3288# 0.378221f
C142 plus.n57 a_n3394_n3288# 0.008984f
C143 plus.n58 a_n3394_n3288# 0.039593f
C144 plus.n59 a_n3394_n3288# 0.039593f
C145 plus.n60 a_n3394_n3288# 0.039593f
C146 plus.n61 a_n3394_n3288# 0.008984f
C147 plus.n62 a_n3394_n3288# 0.378221f
C148 plus.n63 a_n3394_n3288# 0.008984f
C149 plus.n64 a_n3394_n3288# 0.039593f
C150 plus.n65 a_n3394_n3288# 0.039593f
C151 plus.n66 a_n3394_n3288# 0.039593f
C152 plus.n67 a_n3394_n3288# 0.008984f
C153 plus.n68 a_n3394_n3288# 0.378221f
C154 plus.n69 a_n3394_n3288# 0.008984f
C155 plus.n70 a_n3394_n3288# 0.039593f
C156 plus.n71 a_n3394_n3288# 0.039593f
C157 plus.n72 a_n3394_n3288# 0.039593f
C158 plus.n73 a_n3394_n3288# 0.008984f
C159 plus.n74 a_n3394_n3288# 0.378221f
C160 plus.n75 a_n3394_n3288# 0.008984f
C161 plus.n76 a_n3394_n3288# 0.039593f
C162 plus.n77 a_n3394_n3288# 0.039593f
C163 plus.n78 a_n3394_n3288# 0.039593f
C164 plus.n79 a_n3394_n3288# 0.008984f
C165 plus.n80 a_n3394_n3288# 0.378221f
C166 plus.n81 a_n3394_n3288# 0.008984f
C167 plus.n82 a_n3394_n3288# 0.378587f
C168 plus.n83 a_n3394_n3288# 1.51961f
C169 source.n0 a_n3394_n3288# 0.032909f
C170 source.n1 a_n3394_n3288# 0.024844f
C171 source.n2 a_n3394_n3288# 0.01335f
C172 source.n3 a_n3394_n3288# 0.031555f
C173 source.n4 a_n3394_n3288# 0.014135f
C174 source.n5 a_n3394_n3288# 0.024844f
C175 source.n6 a_n3394_n3288# 0.01335f
C176 source.n7 a_n3394_n3288# 0.031555f
C177 source.n8 a_n3394_n3288# 0.014135f
C178 source.n9 a_n3394_n3288# 0.024844f
C179 source.n10 a_n3394_n3288# 0.013743f
C180 source.n11 a_n3394_n3288# 0.031555f
C181 source.n12 a_n3394_n3288# 0.01335f
C182 source.n13 a_n3394_n3288# 0.014135f
C183 source.n14 a_n3394_n3288# 0.024844f
C184 source.n15 a_n3394_n3288# 0.01335f
C185 source.n16 a_n3394_n3288# 0.031555f
C186 source.n17 a_n3394_n3288# 0.014135f
C187 source.n18 a_n3394_n3288# 0.024844f
C188 source.n19 a_n3394_n3288# 0.01335f
C189 source.n20 a_n3394_n3288# 0.023666f
C190 source.n21 a_n3394_n3288# 0.022307f
C191 source.t22 a_n3394_n3288# 0.053294f
C192 source.n22 a_n3394_n3288# 0.179123f
C193 source.n23 a_n3394_n3288# 1.25334f
C194 source.n24 a_n3394_n3288# 0.01335f
C195 source.n25 a_n3394_n3288# 0.014135f
C196 source.n26 a_n3394_n3288# 0.031555f
C197 source.n27 a_n3394_n3288# 0.031555f
C198 source.n28 a_n3394_n3288# 0.014135f
C199 source.n29 a_n3394_n3288# 0.01335f
C200 source.n30 a_n3394_n3288# 0.024844f
C201 source.n31 a_n3394_n3288# 0.024844f
C202 source.n32 a_n3394_n3288# 0.01335f
C203 source.n33 a_n3394_n3288# 0.014135f
C204 source.n34 a_n3394_n3288# 0.031555f
C205 source.n35 a_n3394_n3288# 0.031555f
C206 source.n36 a_n3394_n3288# 0.014135f
C207 source.n37 a_n3394_n3288# 0.01335f
C208 source.n38 a_n3394_n3288# 0.024844f
C209 source.n39 a_n3394_n3288# 0.024844f
C210 source.n40 a_n3394_n3288# 0.01335f
C211 source.n41 a_n3394_n3288# 0.014135f
C212 source.n42 a_n3394_n3288# 0.031555f
C213 source.n43 a_n3394_n3288# 0.031555f
C214 source.n44 a_n3394_n3288# 0.031555f
C215 source.n45 a_n3394_n3288# 0.013743f
C216 source.n46 a_n3394_n3288# 0.01335f
C217 source.n47 a_n3394_n3288# 0.024844f
C218 source.n48 a_n3394_n3288# 0.024844f
C219 source.n49 a_n3394_n3288# 0.01335f
C220 source.n50 a_n3394_n3288# 0.014135f
C221 source.n51 a_n3394_n3288# 0.031555f
C222 source.n52 a_n3394_n3288# 0.031555f
C223 source.n53 a_n3394_n3288# 0.014135f
C224 source.n54 a_n3394_n3288# 0.01335f
C225 source.n55 a_n3394_n3288# 0.024844f
C226 source.n56 a_n3394_n3288# 0.024844f
C227 source.n57 a_n3394_n3288# 0.01335f
C228 source.n58 a_n3394_n3288# 0.014135f
C229 source.n59 a_n3394_n3288# 0.031555f
C230 source.n60 a_n3394_n3288# 0.064754f
C231 source.n61 a_n3394_n3288# 0.014135f
C232 source.n62 a_n3394_n3288# 0.01335f
C233 source.n63 a_n3394_n3288# 0.053353f
C234 source.n64 a_n3394_n3288# 0.035737f
C235 source.n65 a_n3394_n3288# 1.0451f
C236 source.t13 a_n3394_n3288# 0.23559f
C237 source.t9 a_n3394_n3288# 0.23559f
C238 source.n66 a_n3394_n3288# 2.01713f
C239 source.n67 a_n3394_n3288# 0.396162f
C240 source.t14 a_n3394_n3288# 0.23559f
C241 source.t6 a_n3394_n3288# 0.23559f
C242 source.n68 a_n3394_n3288# 2.01713f
C243 source.n69 a_n3394_n3288# 0.396162f
C244 source.t15 a_n3394_n3288# 0.23559f
C245 source.t12 a_n3394_n3288# 0.23559f
C246 source.n70 a_n3394_n3288# 2.01713f
C247 source.n71 a_n3394_n3288# 0.396162f
C248 source.t16 a_n3394_n3288# 0.23559f
C249 source.t17 a_n3394_n3288# 0.23559f
C250 source.n72 a_n3394_n3288# 2.01713f
C251 source.n73 a_n3394_n3288# 0.396162f
C252 source.t5 a_n3394_n3288# 0.23559f
C253 source.t11 a_n3394_n3288# 0.23559f
C254 source.n74 a_n3394_n3288# 2.01713f
C255 source.n75 a_n3394_n3288# 0.396162f
C256 source.n76 a_n3394_n3288# 0.032909f
C257 source.n77 a_n3394_n3288# 0.024844f
C258 source.n78 a_n3394_n3288# 0.01335f
C259 source.n79 a_n3394_n3288# 0.031555f
C260 source.n80 a_n3394_n3288# 0.014135f
C261 source.n81 a_n3394_n3288# 0.024844f
C262 source.n82 a_n3394_n3288# 0.01335f
C263 source.n83 a_n3394_n3288# 0.031555f
C264 source.n84 a_n3394_n3288# 0.014135f
C265 source.n85 a_n3394_n3288# 0.024844f
C266 source.n86 a_n3394_n3288# 0.013743f
C267 source.n87 a_n3394_n3288# 0.031555f
C268 source.n88 a_n3394_n3288# 0.01335f
C269 source.n89 a_n3394_n3288# 0.014135f
C270 source.n90 a_n3394_n3288# 0.024844f
C271 source.n91 a_n3394_n3288# 0.01335f
C272 source.n92 a_n3394_n3288# 0.031555f
C273 source.n93 a_n3394_n3288# 0.014135f
C274 source.n94 a_n3394_n3288# 0.024844f
C275 source.n95 a_n3394_n3288# 0.01335f
C276 source.n96 a_n3394_n3288# 0.023666f
C277 source.n97 a_n3394_n3288# 0.022307f
C278 source.t0 a_n3394_n3288# 0.053294f
C279 source.n98 a_n3394_n3288# 0.179123f
C280 source.n99 a_n3394_n3288# 1.25334f
C281 source.n100 a_n3394_n3288# 0.01335f
C282 source.n101 a_n3394_n3288# 0.014135f
C283 source.n102 a_n3394_n3288# 0.031555f
C284 source.n103 a_n3394_n3288# 0.031555f
C285 source.n104 a_n3394_n3288# 0.014135f
C286 source.n105 a_n3394_n3288# 0.01335f
C287 source.n106 a_n3394_n3288# 0.024844f
C288 source.n107 a_n3394_n3288# 0.024844f
C289 source.n108 a_n3394_n3288# 0.01335f
C290 source.n109 a_n3394_n3288# 0.014135f
C291 source.n110 a_n3394_n3288# 0.031555f
C292 source.n111 a_n3394_n3288# 0.031555f
C293 source.n112 a_n3394_n3288# 0.014135f
C294 source.n113 a_n3394_n3288# 0.01335f
C295 source.n114 a_n3394_n3288# 0.024844f
C296 source.n115 a_n3394_n3288# 0.024844f
C297 source.n116 a_n3394_n3288# 0.01335f
C298 source.n117 a_n3394_n3288# 0.014135f
C299 source.n118 a_n3394_n3288# 0.031555f
C300 source.n119 a_n3394_n3288# 0.031555f
C301 source.n120 a_n3394_n3288# 0.031555f
C302 source.n121 a_n3394_n3288# 0.013743f
C303 source.n122 a_n3394_n3288# 0.01335f
C304 source.n123 a_n3394_n3288# 0.024844f
C305 source.n124 a_n3394_n3288# 0.024844f
C306 source.n125 a_n3394_n3288# 0.01335f
C307 source.n126 a_n3394_n3288# 0.014135f
C308 source.n127 a_n3394_n3288# 0.031555f
C309 source.n128 a_n3394_n3288# 0.031555f
C310 source.n129 a_n3394_n3288# 0.014135f
C311 source.n130 a_n3394_n3288# 0.01335f
C312 source.n131 a_n3394_n3288# 0.024844f
C313 source.n132 a_n3394_n3288# 0.024844f
C314 source.n133 a_n3394_n3288# 0.01335f
C315 source.n134 a_n3394_n3288# 0.014135f
C316 source.n135 a_n3394_n3288# 0.031555f
C317 source.n136 a_n3394_n3288# 0.064754f
C318 source.n137 a_n3394_n3288# 0.014135f
C319 source.n138 a_n3394_n3288# 0.01335f
C320 source.n139 a_n3394_n3288# 0.053353f
C321 source.n140 a_n3394_n3288# 0.035737f
C322 source.n141 a_n3394_n3288# 0.127617f
C323 source.n142 a_n3394_n3288# 0.032909f
C324 source.n143 a_n3394_n3288# 0.024844f
C325 source.n144 a_n3394_n3288# 0.01335f
C326 source.n145 a_n3394_n3288# 0.031555f
C327 source.n146 a_n3394_n3288# 0.014135f
C328 source.n147 a_n3394_n3288# 0.024844f
C329 source.n148 a_n3394_n3288# 0.01335f
C330 source.n149 a_n3394_n3288# 0.031555f
C331 source.n150 a_n3394_n3288# 0.014135f
C332 source.n151 a_n3394_n3288# 0.024844f
C333 source.n152 a_n3394_n3288# 0.013743f
C334 source.n153 a_n3394_n3288# 0.031555f
C335 source.n154 a_n3394_n3288# 0.01335f
C336 source.n155 a_n3394_n3288# 0.014135f
C337 source.n156 a_n3394_n3288# 0.024844f
C338 source.n157 a_n3394_n3288# 0.01335f
C339 source.n158 a_n3394_n3288# 0.031555f
C340 source.n159 a_n3394_n3288# 0.014135f
C341 source.n160 a_n3394_n3288# 0.024844f
C342 source.n161 a_n3394_n3288# 0.01335f
C343 source.n162 a_n3394_n3288# 0.023666f
C344 source.n163 a_n3394_n3288# 0.022307f
C345 source.t34 a_n3394_n3288# 0.053294f
C346 source.n164 a_n3394_n3288# 0.179123f
C347 source.n165 a_n3394_n3288# 1.25334f
C348 source.n166 a_n3394_n3288# 0.01335f
C349 source.n167 a_n3394_n3288# 0.014135f
C350 source.n168 a_n3394_n3288# 0.031555f
C351 source.n169 a_n3394_n3288# 0.031555f
C352 source.n170 a_n3394_n3288# 0.014135f
C353 source.n171 a_n3394_n3288# 0.01335f
C354 source.n172 a_n3394_n3288# 0.024844f
C355 source.n173 a_n3394_n3288# 0.024844f
C356 source.n174 a_n3394_n3288# 0.01335f
C357 source.n175 a_n3394_n3288# 0.014135f
C358 source.n176 a_n3394_n3288# 0.031555f
C359 source.n177 a_n3394_n3288# 0.031555f
C360 source.n178 a_n3394_n3288# 0.014135f
C361 source.n179 a_n3394_n3288# 0.01335f
C362 source.n180 a_n3394_n3288# 0.024844f
C363 source.n181 a_n3394_n3288# 0.024844f
C364 source.n182 a_n3394_n3288# 0.01335f
C365 source.n183 a_n3394_n3288# 0.014135f
C366 source.n184 a_n3394_n3288# 0.031555f
C367 source.n185 a_n3394_n3288# 0.031555f
C368 source.n186 a_n3394_n3288# 0.031555f
C369 source.n187 a_n3394_n3288# 0.013743f
C370 source.n188 a_n3394_n3288# 0.01335f
C371 source.n189 a_n3394_n3288# 0.024844f
C372 source.n190 a_n3394_n3288# 0.024844f
C373 source.n191 a_n3394_n3288# 0.01335f
C374 source.n192 a_n3394_n3288# 0.014135f
C375 source.n193 a_n3394_n3288# 0.031555f
C376 source.n194 a_n3394_n3288# 0.031555f
C377 source.n195 a_n3394_n3288# 0.014135f
C378 source.n196 a_n3394_n3288# 0.01335f
C379 source.n197 a_n3394_n3288# 0.024844f
C380 source.n198 a_n3394_n3288# 0.024844f
C381 source.n199 a_n3394_n3288# 0.01335f
C382 source.n200 a_n3394_n3288# 0.014135f
C383 source.n201 a_n3394_n3288# 0.031555f
C384 source.n202 a_n3394_n3288# 0.064754f
C385 source.n203 a_n3394_n3288# 0.014135f
C386 source.n204 a_n3394_n3288# 0.01335f
C387 source.n205 a_n3394_n3288# 0.053353f
C388 source.n206 a_n3394_n3288# 0.035737f
C389 source.n207 a_n3394_n3288# 0.127617f
C390 source.t37 a_n3394_n3288# 0.23559f
C391 source.t44 a_n3394_n3288# 0.23559f
C392 source.n208 a_n3394_n3288# 2.01713f
C393 source.n209 a_n3394_n3288# 0.396162f
C394 source.t38 a_n3394_n3288# 0.23559f
C395 source.t26 a_n3394_n3288# 0.23559f
C396 source.n210 a_n3394_n3288# 2.01713f
C397 source.n211 a_n3394_n3288# 0.396162f
C398 source.t39 a_n3394_n3288# 0.23559f
C399 source.t25 a_n3394_n3288# 0.23559f
C400 source.n212 a_n3394_n3288# 2.01713f
C401 source.n213 a_n3394_n3288# 0.396162f
C402 source.t40 a_n3394_n3288# 0.23559f
C403 source.t29 a_n3394_n3288# 0.23559f
C404 source.n214 a_n3394_n3288# 2.01713f
C405 source.n215 a_n3394_n3288# 0.396162f
C406 source.t42 a_n3394_n3288# 0.23559f
C407 source.t32 a_n3394_n3288# 0.23559f
C408 source.n216 a_n3394_n3288# 2.01713f
C409 source.n217 a_n3394_n3288# 0.396162f
C410 source.n218 a_n3394_n3288# 0.032909f
C411 source.n219 a_n3394_n3288# 0.024844f
C412 source.n220 a_n3394_n3288# 0.01335f
C413 source.n221 a_n3394_n3288# 0.031555f
C414 source.n222 a_n3394_n3288# 0.014135f
C415 source.n223 a_n3394_n3288# 0.024844f
C416 source.n224 a_n3394_n3288# 0.01335f
C417 source.n225 a_n3394_n3288# 0.031555f
C418 source.n226 a_n3394_n3288# 0.014135f
C419 source.n227 a_n3394_n3288# 0.024844f
C420 source.n228 a_n3394_n3288# 0.013743f
C421 source.n229 a_n3394_n3288# 0.031555f
C422 source.n230 a_n3394_n3288# 0.01335f
C423 source.n231 a_n3394_n3288# 0.014135f
C424 source.n232 a_n3394_n3288# 0.024844f
C425 source.n233 a_n3394_n3288# 0.01335f
C426 source.n234 a_n3394_n3288# 0.031555f
C427 source.n235 a_n3394_n3288# 0.014135f
C428 source.n236 a_n3394_n3288# 0.024844f
C429 source.n237 a_n3394_n3288# 0.01335f
C430 source.n238 a_n3394_n3288# 0.023666f
C431 source.n239 a_n3394_n3288# 0.022307f
C432 source.t33 a_n3394_n3288# 0.053294f
C433 source.n240 a_n3394_n3288# 0.179123f
C434 source.n241 a_n3394_n3288# 1.25334f
C435 source.n242 a_n3394_n3288# 0.01335f
C436 source.n243 a_n3394_n3288# 0.014135f
C437 source.n244 a_n3394_n3288# 0.031555f
C438 source.n245 a_n3394_n3288# 0.031555f
C439 source.n246 a_n3394_n3288# 0.014135f
C440 source.n247 a_n3394_n3288# 0.01335f
C441 source.n248 a_n3394_n3288# 0.024844f
C442 source.n249 a_n3394_n3288# 0.024844f
C443 source.n250 a_n3394_n3288# 0.01335f
C444 source.n251 a_n3394_n3288# 0.014135f
C445 source.n252 a_n3394_n3288# 0.031555f
C446 source.n253 a_n3394_n3288# 0.031555f
C447 source.n254 a_n3394_n3288# 0.014135f
C448 source.n255 a_n3394_n3288# 0.01335f
C449 source.n256 a_n3394_n3288# 0.024844f
C450 source.n257 a_n3394_n3288# 0.024844f
C451 source.n258 a_n3394_n3288# 0.01335f
C452 source.n259 a_n3394_n3288# 0.014135f
C453 source.n260 a_n3394_n3288# 0.031555f
C454 source.n261 a_n3394_n3288# 0.031555f
C455 source.n262 a_n3394_n3288# 0.031555f
C456 source.n263 a_n3394_n3288# 0.013743f
C457 source.n264 a_n3394_n3288# 0.01335f
C458 source.n265 a_n3394_n3288# 0.024844f
C459 source.n266 a_n3394_n3288# 0.024844f
C460 source.n267 a_n3394_n3288# 0.01335f
C461 source.n268 a_n3394_n3288# 0.014135f
C462 source.n269 a_n3394_n3288# 0.031555f
C463 source.n270 a_n3394_n3288# 0.031555f
C464 source.n271 a_n3394_n3288# 0.014135f
C465 source.n272 a_n3394_n3288# 0.01335f
C466 source.n273 a_n3394_n3288# 0.024844f
C467 source.n274 a_n3394_n3288# 0.024844f
C468 source.n275 a_n3394_n3288# 0.01335f
C469 source.n276 a_n3394_n3288# 0.014135f
C470 source.n277 a_n3394_n3288# 0.031555f
C471 source.n278 a_n3394_n3288# 0.064754f
C472 source.n279 a_n3394_n3288# 0.014135f
C473 source.n280 a_n3394_n3288# 0.01335f
C474 source.n281 a_n3394_n3288# 0.053353f
C475 source.n282 a_n3394_n3288# 0.035737f
C476 source.n283 a_n3394_n3288# 1.44571f
C477 source.n284 a_n3394_n3288# 0.032909f
C478 source.n285 a_n3394_n3288# 0.024844f
C479 source.n286 a_n3394_n3288# 0.01335f
C480 source.n287 a_n3394_n3288# 0.031555f
C481 source.n288 a_n3394_n3288# 0.014135f
C482 source.n289 a_n3394_n3288# 0.024844f
C483 source.n290 a_n3394_n3288# 0.01335f
C484 source.n291 a_n3394_n3288# 0.031555f
C485 source.n292 a_n3394_n3288# 0.014135f
C486 source.n293 a_n3394_n3288# 0.024844f
C487 source.n294 a_n3394_n3288# 0.013743f
C488 source.n295 a_n3394_n3288# 0.031555f
C489 source.n296 a_n3394_n3288# 0.014135f
C490 source.n297 a_n3394_n3288# 0.024844f
C491 source.n298 a_n3394_n3288# 0.01335f
C492 source.n299 a_n3394_n3288# 0.031555f
C493 source.n300 a_n3394_n3288# 0.014135f
C494 source.n301 a_n3394_n3288# 0.024844f
C495 source.n302 a_n3394_n3288# 0.01335f
C496 source.n303 a_n3394_n3288# 0.023666f
C497 source.n304 a_n3394_n3288# 0.022307f
C498 source.t7 a_n3394_n3288# 0.053294f
C499 source.n305 a_n3394_n3288# 0.179123f
C500 source.n306 a_n3394_n3288# 1.25334f
C501 source.n307 a_n3394_n3288# 0.01335f
C502 source.n308 a_n3394_n3288# 0.014135f
C503 source.n309 a_n3394_n3288# 0.031555f
C504 source.n310 a_n3394_n3288# 0.031555f
C505 source.n311 a_n3394_n3288# 0.014135f
C506 source.n312 a_n3394_n3288# 0.01335f
C507 source.n313 a_n3394_n3288# 0.024844f
C508 source.n314 a_n3394_n3288# 0.024844f
C509 source.n315 a_n3394_n3288# 0.01335f
C510 source.n316 a_n3394_n3288# 0.014135f
C511 source.n317 a_n3394_n3288# 0.031555f
C512 source.n318 a_n3394_n3288# 0.031555f
C513 source.n319 a_n3394_n3288# 0.014135f
C514 source.n320 a_n3394_n3288# 0.01335f
C515 source.n321 a_n3394_n3288# 0.024844f
C516 source.n322 a_n3394_n3288# 0.024844f
C517 source.n323 a_n3394_n3288# 0.01335f
C518 source.n324 a_n3394_n3288# 0.01335f
C519 source.n325 a_n3394_n3288# 0.014135f
C520 source.n326 a_n3394_n3288# 0.031555f
C521 source.n327 a_n3394_n3288# 0.031555f
C522 source.n328 a_n3394_n3288# 0.031555f
C523 source.n329 a_n3394_n3288# 0.013743f
C524 source.n330 a_n3394_n3288# 0.01335f
C525 source.n331 a_n3394_n3288# 0.024844f
C526 source.n332 a_n3394_n3288# 0.024844f
C527 source.n333 a_n3394_n3288# 0.01335f
C528 source.n334 a_n3394_n3288# 0.014135f
C529 source.n335 a_n3394_n3288# 0.031555f
C530 source.n336 a_n3394_n3288# 0.031555f
C531 source.n337 a_n3394_n3288# 0.014135f
C532 source.n338 a_n3394_n3288# 0.01335f
C533 source.n339 a_n3394_n3288# 0.024844f
C534 source.n340 a_n3394_n3288# 0.024844f
C535 source.n341 a_n3394_n3288# 0.01335f
C536 source.n342 a_n3394_n3288# 0.014135f
C537 source.n343 a_n3394_n3288# 0.031555f
C538 source.n344 a_n3394_n3288# 0.064754f
C539 source.n345 a_n3394_n3288# 0.014135f
C540 source.n346 a_n3394_n3288# 0.01335f
C541 source.n347 a_n3394_n3288# 0.053353f
C542 source.n348 a_n3394_n3288# 0.035737f
C543 source.n349 a_n3394_n3288# 1.44571f
C544 source.t19 a_n3394_n3288# 0.23559f
C545 source.t8 a_n3394_n3288# 0.23559f
C546 source.n350 a_n3394_n3288# 2.01712f
C547 source.n351 a_n3394_n3288# 0.396174f
C548 source.t2 a_n3394_n3288# 0.23559f
C549 source.t21 a_n3394_n3288# 0.23559f
C550 source.n352 a_n3394_n3288# 2.01712f
C551 source.n353 a_n3394_n3288# 0.396174f
C552 source.t23 a_n3394_n3288# 0.23559f
C553 source.t10 a_n3394_n3288# 0.23559f
C554 source.n354 a_n3394_n3288# 2.01712f
C555 source.n355 a_n3394_n3288# 0.396174f
C556 source.t1 a_n3394_n3288# 0.23559f
C557 source.t20 a_n3394_n3288# 0.23559f
C558 source.n356 a_n3394_n3288# 2.01712f
C559 source.n357 a_n3394_n3288# 0.396174f
C560 source.t4 a_n3394_n3288# 0.23559f
C561 source.t3 a_n3394_n3288# 0.23559f
C562 source.n358 a_n3394_n3288# 2.01712f
C563 source.n359 a_n3394_n3288# 0.396174f
C564 source.n360 a_n3394_n3288# 0.032909f
C565 source.n361 a_n3394_n3288# 0.024844f
C566 source.n362 a_n3394_n3288# 0.01335f
C567 source.n363 a_n3394_n3288# 0.031555f
C568 source.n364 a_n3394_n3288# 0.014135f
C569 source.n365 a_n3394_n3288# 0.024844f
C570 source.n366 a_n3394_n3288# 0.01335f
C571 source.n367 a_n3394_n3288# 0.031555f
C572 source.n368 a_n3394_n3288# 0.014135f
C573 source.n369 a_n3394_n3288# 0.024844f
C574 source.n370 a_n3394_n3288# 0.013743f
C575 source.n371 a_n3394_n3288# 0.031555f
C576 source.n372 a_n3394_n3288# 0.014135f
C577 source.n373 a_n3394_n3288# 0.024844f
C578 source.n374 a_n3394_n3288# 0.01335f
C579 source.n375 a_n3394_n3288# 0.031555f
C580 source.n376 a_n3394_n3288# 0.014135f
C581 source.n377 a_n3394_n3288# 0.024844f
C582 source.n378 a_n3394_n3288# 0.01335f
C583 source.n379 a_n3394_n3288# 0.023666f
C584 source.n380 a_n3394_n3288# 0.022307f
C585 source.t18 a_n3394_n3288# 0.053294f
C586 source.n381 a_n3394_n3288# 0.179123f
C587 source.n382 a_n3394_n3288# 1.25334f
C588 source.n383 a_n3394_n3288# 0.01335f
C589 source.n384 a_n3394_n3288# 0.014135f
C590 source.n385 a_n3394_n3288# 0.031555f
C591 source.n386 a_n3394_n3288# 0.031555f
C592 source.n387 a_n3394_n3288# 0.014135f
C593 source.n388 a_n3394_n3288# 0.01335f
C594 source.n389 a_n3394_n3288# 0.024844f
C595 source.n390 a_n3394_n3288# 0.024844f
C596 source.n391 a_n3394_n3288# 0.01335f
C597 source.n392 a_n3394_n3288# 0.014135f
C598 source.n393 a_n3394_n3288# 0.031555f
C599 source.n394 a_n3394_n3288# 0.031555f
C600 source.n395 a_n3394_n3288# 0.014135f
C601 source.n396 a_n3394_n3288# 0.01335f
C602 source.n397 a_n3394_n3288# 0.024844f
C603 source.n398 a_n3394_n3288# 0.024844f
C604 source.n399 a_n3394_n3288# 0.01335f
C605 source.n400 a_n3394_n3288# 0.01335f
C606 source.n401 a_n3394_n3288# 0.014135f
C607 source.n402 a_n3394_n3288# 0.031555f
C608 source.n403 a_n3394_n3288# 0.031555f
C609 source.n404 a_n3394_n3288# 0.031555f
C610 source.n405 a_n3394_n3288# 0.013743f
C611 source.n406 a_n3394_n3288# 0.01335f
C612 source.n407 a_n3394_n3288# 0.024844f
C613 source.n408 a_n3394_n3288# 0.024844f
C614 source.n409 a_n3394_n3288# 0.01335f
C615 source.n410 a_n3394_n3288# 0.014135f
C616 source.n411 a_n3394_n3288# 0.031555f
C617 source.n412 a_n3394_n3288# 0.031555f
C618 source.n413 a_n3394_n3288# 0.014135f
C619 source.n414 a_n3394_n3288# 0.01335f
C620 source.n415 a_n3394_n3288# 0.024844f
C621 source.n416 a_n3394_n3288# 0.024844f
C622 source.n417 a_n3394_n3288# 0.01335f
C623 source.n418 a_n3394_n3288# 0.014135f
C624 source.n419 a_n3394_n3288# 0.031555f
C625 source.n420 a_n3394_n3288# 0.064754f
C626 source.n421 a_n3394_n3288# 0.014135f
C627 source.n422 a_n3394_n3288# 0.01335f
C628 source.n423 a_n3394_n3288# 0.053353f
C629 source.n424 a_n3394_n3288# 0.035737f
C630 source.n425 a_n3394_n3288# 0.127617f
C631 source.n426 a_n3394_n3288# 0.032909f
C632 source.n427 a_n3394_n3288# 0.024844f
C633 source.n428 a_n3394_n3288# 0.01335f
C634 source.n429 a_n3394_n3288# 0.031555f
C635 source.n430 a_n3394_n3288# 0.014135f
C636 source.n431 a_n3394_n3288# 0.024844f
C637 source.n432 a_n3394_n3288# 0.01335f
C638 source.n433 a_n3394_n3288# 0.031555f
C639 source.n434 a_n3394_n3288# 0.014135f
C640 source.n435 a_n3394_n3288# 0.024844f
C641 source.n436 a_n3394_n3288# 0.013743f
C642 source.n437 a_n3394_n3288# 0.031555f
C643 source.n438 a_n3394_n3288# 0.014135f
C644 source.n439 a_n3394_n3288# 0.024844f
C645 source.n440 a_n3394_n3288# 0.01335f
C646 source.n441 a_n3394_n3288# 0.031555f
C647 source.n442 a_n3394_n3288# 0.014135f
C648 source.n443 a_n3394_n3288# 0.024844f
C649 source.n444 a_n3394_n3288# 0.01335f
C650 source.n445 a_n3394_n3288# 0.023666f
C651 source.n446 a_n3394_n3288# 0.022307f
C652 source.t45 a_n3394_n3288# 0.053294f
C653 source.n447 a_n3394_n3288# 0.179123f
C654 source.n448 a_n3394_n3288# 1.25334f
C655 source.n449 a_n3394_n3288# 0.01335f
C656 source.n450 a_n3394_n3288# 0.014135f
C657 source.n451 a_n3394_n3288# 0.031555f
C658 source.n452 a_n3394_n3288# 0.031555f
C659 source.n453 a_n3394_n3288# 0.014135f
C660 source.n454 a_n3394_n3288# 0.01335f
C661 source.n455 a_n3394_n3288# 0.024844f
C662 source.n456 a_n3394_n3288# 0.024844f
C663 source.n457 a_n3394_n3288# 0.01335f
C664 source.n458 a_n3394_n3288# 0.014135f
C665 source.n459 a_n3394_n3288# 0.031555f
C666 source.n460 a_n3394_n3288# 0.031555f
C667 source.n461 a_n3394_n3288# 0.014135f
C668 source.n462 a_n3394_n3288# 0.01335f
C669 source.n463 a_n3394_n3288# 0.024844f
C670 source.n464 a_n3394_n3288# 0.024844f
C671 source.n465 a_n3394_n3288# 0.01335f
C672 source.n466 a_n3394_n3288# 0.01335f
C673 source.n467 a_n3394_n3288# 0.014135f
C674 source.n468 a_n3394_n3288# 0.031555f
C675 source.n469 a_n3394_n3288# 0.031555f
C676 source.n470 a_n3394_n3288# 0.031555f
C677 source.n471 a_n3394_n3288# 0.013743f
C678 source.n472 a_n3394_n3288# 0.01335f
C679 source.n473 a_n3394_n3288# 0.024844f
C680 source.n474 a_n3394_n3288# 0.024844f
C681 source.n475 a_n3394_n3288# 0.01335f
C682 source.n476 a_n3394_n3288# 0.014135f
C683 source.n477 a_n3394_n3288# 0.031555f
C684 source.n478 a_n3394_n3288# 0.031555f
C685 source.n479 a_n3394_n3288# 0.014135f
C686 source.n480 a_n3394_n3288# 0.01335f
C687 source.n481 a_n3394_n3288# 0.024844f
C688 source.n482 a_n3394_n3288# 0.024844f
C689 source.n483 a_n3394_n3288# 0.01335f
C690 source.n484 a_n3394_n3288# 0.014135f
C691 source.n485 a_n3394_n3288# 0.031555f
C692 source.n486 a_n3394_n3288# 0.064754f
C693 source.n487 a_n3394_n3288# 0.014135f
C694 source.n488 a_n3394_n3288# 0.01335f
C695 source.n489 a_n3394_n3288# 0.053353f
C696 source.n490 a_n3394_n3288# 0.035737f
C697 source.n491 a_n3394_n3288# 0.127617f
C698 source.t43 a_n3394_n3288# 0.23559f
C699 source.t28 a_n3394_n3288# 0.23559f
C700 source.n492 a_n3394_n3288# 2.01712f
C701 source.n493 a_n3394_n3288# 0.396174f
C702 source.t27 a_n3394_n3288# 0.23559f
C703 source.t24 a_n3394_n3288# 0.23559f
C704 source.n494 a_n3394_n3288# 2.01712f
C705 source.n495 a_n3394_n3288# 0.396174f
C706 source.t31 a_n3394_n3288# 0.23559f
C707 source.t30 a_n3394_n3288# 0.23559f
C708 source.n496 a_n3394_n3288# 2.01712f
C709 source.n497 a_n3394_n3288# 0.396174f
C710 source.t35 a_n3394_n3288# 0.23559f
C711 source.t36 a_n3394_n3288# 0.23559f
C712 source.n498 a_n3394_n3288# 2.01712f
C713 source.n499 a_n3394_n3288# 0.396174f
C714 source.t41 a_n3394_n3288# 0.23559f
C715 source.t47 a_n3394_n3288# 0.23559f
C716 source.n500 a_n3394_n3288# 2.01712f
C717 source.n501 a_n3394_n3288# 0.396174f
C718 source.n502 a_n3394_n3288# 0.032909f
C719 source.n503 a_n3394_n3288# 0.024844f
C720 source.n504 a_n3394_n3288# 0.01335f
C721 source.n505 a_n3394_n3288# 0.031555f
C722 source.n506 a_n3394_n3288# 0.014135f
C723 source.n507 a_n3394_n3288# 0.024844f
C724 source.n508 a_n3394_n3288# 0.01335f
C725 source.n509 a_n3394_n3288# 0.031555f
C726 source.n510 a_n3394_n3288# 0.014135f
C727 source.n511 a_n3394_n3288# 0.024844f
C728 source.n512 a_n3394_n3288# 0.013743f
C729 source.n513 a_n3394_n3288# 0.031555f
C730 source.n514 a_n3394_n3288# 0.014135f
C731 source.n515 a_n3394_n3288# 0.024844f
C732 source.n516 a_n3394_n3288# 0.01335f
C733 source.n517 a_n3394_n3288# 0.031555f
C734 source.n518 a_n3394_n3288# 0.014135f
C735 source.n519 a_n3394_n3288# 0.024844f
C736 source.n520 a_n3394_n3288# 0.01335f
C737 source.n521 a_n3394_n3288# 0.023666f
C738 source.n522 a_n3394_n3288# 0.022307f
C739 source.t46 a_n3394_n3288# 0.053294f
C740 source.n523 a_n3394_n3288# 0.179123f
C741 source.n524 a_n3394_n3288# 1.25334f
C742 source.n525 a_n3394_n3288# 0.01335f
C743 source.n526 a_n3394_n3288# 0.014135f
C744 source.n527 a_n3394_n3288# 0.031555f
C745 source.n528 a_n3394_n3288# 0.031555f
C746 source.n529 a_n3394_n3288# 0.014135f
C747 source.n530 a_n3394_n3288# 0.01335f
C748 source.n531 a_n3394_n3288# 0.024844f
C749 source.n532 a_n3394_n3288# 0.024844f
C750 source.n533 a_n3394_n3288# 0.01335f
C751 source.n534 a_n3394_n3288# 0.014135f
C752 source.n535 a_n3394_n3288# 0.031555f
C753 source.n536 a_n3394_n3288# 0.031555f
C754 source.n537 a_n3394_n3288# 0.014135f
C755 source.n538 a_n3394_n3288# 0.01335f
C756 source.n539 a_n3394_n3288# 0.024844f
C757 source.n540 a_n3394_n3288# 0.024844f
C758 source.n541 a_n3394_n3288# 0.01335f
C759 source.n542 a_n3394_n3288# 0.01335f
C760 source.n543 a_n3394_n3288# 0.014135f
C761 source.n544 a_n3394_n3288# 0.031555f
C762 source.n545 a_n3394_n3288# 0.031555f
C763 source.n546 a_n3394_n3288# 0.031555f
C764 source.n547 a_n3394_n3288# 0.013743f
C765 source.n548 a_n3394_n3288# 0.01335f
C766 source.n549 a_n3394_n3288# 0.024844f
C767 source.n550 a_n3394_n3288# 0.024844f
C768 source.n551 a_n3394_n3288# 0.01335f
C769 source.n552 a_n3394_n3288# 0.014135f
C770 source.n553 a_n3394_n3288# 0.031555f
C771 source.n554 a_n3394_n3288# 0.031555f
C772 source.n555 a_n3394_n3288# 0.014135f
C773 source.n556 a_n3394_n3288# 0.01335f
C774 source.n557 a_n3394_n3288# 0.024844f
C775 source.n558 a_n3394_n3288# 0.024844f
C776 source.n559 a_n3394_n3288# 0.01335f
C777 source.n560 a_n3394_n3288# 0.014135f
C778 source.n561 a_n3394_n3288# 0.031555f
C779 source.n562 a_n3394_n3288# 0.064754f
C780 source.n563 a_n3394_n3288# 0.014135f
C781 source.n564 a_n3394_n3288# 0.01335f
C782 source.n565 a_n3394_n3288# 0.053353f
C783 source.n566 a_n3394_n3288# 0.035737f
C784 source.n567 a_n3394_n3288# 0.289676f
C785 source.n568 a_n3394_n3288# 1.57432f
C786 drain_right.t19 a_n3394_n3288# 0.257652f
C787 drain_right.t3 a_n3394_n3288# 0.257652f
C788 drain_right.n0 a_n3394_n3288# 2.2985f
C789 drain_right.t12 a_n3394_n3288# 0.257652f
C790 drain_right.t17 a_n3394_n3288# 0.257652f
C791 drain_right.n1 a_n3394_n3288# 2.2927f
C792 drain_right.n2 a_n3394_n3288# 0.772162f
C793 drain_right.t20 a_n3394_n3288# 0.257652f
C794 drain_right.t11 a_n3394_n3288# 0.257652f
C795 drain_right.n3 a_n3394_n3288# 2.2927f
C796 drain_right.n4 a_n3394_n3288# 0.341413f
C797 drain_right.t15 a_n3394_n3288# 0.257652f
C798 drain_right.t14 a_n3394_n3288# 0.257652f
C799 drain_right.n5 a_n3394_n3288# 2.2985f
C800 drain_right.t0 a_n3394_n3288# 0.257652f
C801 drain_right.t23 a_n3394_n3288# 0.257652f
C802 drain_right.n6 a_n3394_n3288# 2.2927f
C803 drain_right.n7 a_n3394_n3288# 0.772162f
C804 drain_right.t10 a_n3394_n3288# 0.257652f
C805 drain_right.t7 a_n3394_n3288# 0.257652f
C806 drain_right.n8 a_n3394_n3288# 2.2927f
C807 drain_right.n9 a_n3394_n3288# 0.341413f
C808 drain_right.n10 a_n3394_n3288# 1.73801f
C809 drain_right.t18 a_n3394_n3288# 0.257652f
C810 drain_right.t6 a_n3394_n3288# 0.257652f
C811 drain_right.n11 a_n3394_n3288# 2.2985f
C812 drain_right.t16 a_n3394_n3288# 0.257652f
C813 drain_right.t1 a_n3394_n3288# 0.257652f
C814 drain_right.n12 a_n3394_n3288# 2.29271f
C815 drain_right.n13 a_n3394_n3288# 0.772152f
C816 drain_right.t21 a_n3394_n3288# 0.257652f
C817 drain_right.t8 a_n3394_n3288# 0.257652f
C818 drain_right.n14 a_n3394_n3288# 2.29271f
C819 drain_right.n15 a_n3394_n3288# 0.383497f
C820 drain_right.t13 a_n3394_n3288# 0.257652f
C821 drain_right.t9 a_n3394_n3288# 0.257652f
C822 drain_right.n16 a_n3394_n3288# 2.29271f
C823 drain_right.n17 a_n3394_n3288# 0.383497f
C824 drain_right.t4 a_n3394_n3288# 0.257652f
C825 drain_right.t22 a_n3394_n3288# 0.257652f
C826 drain_right.n18 a_n3394_n3288# 2.29271f
C827 drain_right.n19 a_n3394_n3288# 0.383497f
C828 drain_right.t5 a_n3394_n3288# 0.257652f
C829 drain_right.t2 a_n3394_n3288# 0.257652f
C830 drain_right.n20 a_n3394_n3288# 2.29271f
C831 drain_right.n21 a_n3394_n3288# 0.623822f
C832 minus.n0 a_n3394_n3288# 0.039092f
C833 minus.n1 a_n3394_n3288# 0.008871f
C834 minus.t5 a_n3394_n3288# 0.936365f
C835 minus.n2 a_n3394_n3288# 0.039092f
C836 minus.n3 a_n3394_n3288# 0.008871f
C837 minus.t7 a_n3394_n3288# 0.936365f
C838 minus.n4 a_n3394_n3288# 0.039092f
C839 minus.n5 a_n3394_n3288# 0.008871f
C840 minus.t8 a_n3394_n3288# 0.936365f
C841 minus.n6 a_n3394_n3288# 0.039092f
C842 minus.n7 a_n3394_n3288# 0.008871f
C843 minus.t9 a_n3394_n3288# 0.936365f
C844 minus.n8 a_n3394_n3288# 0.039092f
C845 minus.n9 a_n3394_n3288# 0.008871f
C846 minus.t10 a_n3394_n3288# 0.936365f
C847 minus.t13 a_n3394_n3288# 0.956262f
C848 minus.t3 a_n3394_n3288# 0.936365f
C849 minus.n10 a_n3394_n3288# 0.38144f
C850 minus.n11 a_n3394_n3288# 0.355625f
C851 minus.n12 a_n3394_n3288# 0.168294f
C852 minus.n13 a_n3394_n3288# 0.039092f
C853 minus.n14 a_n3394_n3288# 0.37344f
C854 minus.n15 a_n3394_n3288# 0.008871f
C855 minus.t21 a_n3394_n3288# 0.936365f
C856 minus.n16 a_n3394_n3288# 0.37344f
C857 minus.n17 a_n3394_n3288# 0.039092f
C858 minus.n18 a_n3394_n3288# 0.039092f
C859 minus.n19 a_n3394_n3288# 0.039092f
C860 minus.n20 a_n3394_n3288# 0.37344f
C861 minus.n21 a_n3394_n3288# 0.008871f
C862 minus.t22 a_n3394_n3288# 0.936365f
C863 minus.n22 a_n3394_n3288# 0.37344f
C864 minus.n23 a_n3394_n3288# 0.039092f
C865 minus.n24 a_n3394_n3288# 0.039092f
C866 minus.n25 a_n3394_n3288# 0.039092f
C867 minus.n26 a_n3394_n3288# 0.37344f
C868 minus.n27 a_n3394_n3288# 0.008871f
C869 minus.t18 a_n3394_n3288# 0.936365f
C870 minus.n28 a_n3394_n3288# 0.37344f
C871 minus.n29 a_n3394_n3288# 0.039092f
C872 minus.n30 a_n3394_n3288# 0.039092f
C873 minus.n31 a_n3394_n3288# 0.039092f
C874 minus.n32 a_n3394_n3288# 0.37344f
C875 minus.n33 a_n3394_n3288# 0.008871f
C876 minus.t15 a_n3394_n3288# 0.936365f
C877 minus.n34 a_n3394_n3288# 0.37344f
C878 minus.n35 a_n3394_n3288# 0.039092f
C879 minus.n36 a_n3394_n3288# 0.039092f
C880 minus.n37 a_n3394_n3288# 0.039092f
C881 minus.n38 a_n3394_n3288# 0.37344f
C882 minus.n39 a_n3394_n3288# 0.008871f
C883 minus.t14 a_n3394_n3288# 0.936365f
C884 minus.n40 a_n3394_n3288# 0.373802f
C885 minus.n41 a_n3394_n3288# 1.74534f
C886 minus.n42 a_n3394_n3288# 0.039092f
C887 minus.n43 a_n3394_n3288# 0.008871f
C888 minus.n44 a_n3394_n3288# 0.039092f
C889 minus.n45 a_n3394_n3288# 0.008871f
C890 minus.n46 a_n3394_n3288# 0.039092f
C891 minus.n47 a_n3394_n3288# 0.008871f
C892 minus.n48 a_n3394_n3288# 0.039092f
C893 minus.n49 a_n3394_n3288# 0.008871f
C894 minus.n50 a_n3394_n3288# 0.039092f
C895 minus.n51 a_n3394_n3288# 0.008871f
C896 minus.t2 a_n3394_n3288# 0.956262f
C897 minus.t4 a_n3394_n3288# 0.936365f
C898 minus.n52 a_n3394_n3288# 0.38144f
C899 minus.n53 a_n3394_n3288# 0.355625f
C900 minus.n54 a_n3394_n3288# 0.168294f
C901 minus.n55 a_n3394_n3288# 0.039092f
C902 minus.t19 a_n3394_n3288# 0.936365f
C903 minus.n56 a_n3394_n3288# 0.37344f
C904 minus.n57 a_n3394_n3288# 0.008871f
C905 minus.t20 a_n3394_n3288# 0.936365f
C906 minus.n58 a_n3394_n3288# 0.37344f
C907 minus.n59 a_n3394_n3288# 0.039092f
C908 minus.n60 a_n3394_n3288# 0.039092f
C909 minus.n61 a_n3394_n3288# 0.039092f
C910 minus.t23 a_n3394_n3288# 0.936365f
C911 minus.n62 a_n3394_n3288# 0.37344f
C912 minus.n63 a_n3394_n3288# 0.008871f
C913 minus.t16 a_n3394_n3288# 0.936365f
C914 minus.n64 a_n3394_n3288# 0.37344f
C915 minus.n65 a_n3394_n3288# 0.039092f
C916 minus.n66 a_n3394_n3288# 0.039092f
C917 minus.n67 a_n3394_n3288# 0.039092f
C918 minus.t17 a_n3394_n3288# 0.936365f
C919 minus.n68 a_n3394_n3288# 0.37344f
C920 minus.n69 a_n3394_n3288# 0.008871f
C921 minus.t12 a_n3394_n3288# 0.936365f
C922 minus.n70 a_n3394_n3288# 0.37344f
C923 minus.n71 a_n3394_n3288# 0.039092f
C924 minus.n72 a_n3394_n3288# 0.039092f
C925 minus.n73 a_n3394_n3288# 0.039092f
C926 minus.t11 a_n3394_n3288# 0.936365f
C927 minus.n74 a_n3394_n3288# 0.37344f
C928 minus.n75 a_n3394_n3288# 0.008871f
C929 minus.t6 a_n3394_n3288# 0.936365f
C930 minus.n76 a_n3394_n3288# 0.37344f
C931 minus.n77 a_n3394_n3288# 0.039092f
C932 minus.n78 a_n3394_n3288# 0.039092f
C933 minus.n79 a_n3394_n3288# 0.039092f
C934 minus.t0 a_n3394_n3288# 0.936365f
C935 minus.n80 a_n3394_n3288# 0.37344f
C936 minus.n81 a_n3394_n3288# 0.008871f
C937 minus.t1 a_n3394_n3288# 0.936365f
C938 minus.n82 a_n3394_n3288# 0.373802f
C939 minus.n83 a_n3394_n3288# 0.271881f
C940 minus.n84 a_n3394_n3288# 2.07956f
.ends

