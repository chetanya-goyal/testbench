* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t37 minus.t0 drain_right.t11 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X1 source.t12 plus.t0 drain_left.t19 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X2 drain_left.t18 plus.t1 source.t15 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X3 source.t36 minus.t1 drain_right.t1 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X4 drain_right.t2 minus.t2 source.t35 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X5 drain_right.t16 minus.t3 source.t34 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X6 drain_right.t12 minus.t4 source.t33 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X7 drain_left.t17 plus.t2 source.t3 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X8 source.t7 plus.t3 drain_left.t16 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X9 drain_right.t3 minus.t5 source.t32 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X10 source.t31 minus.t6 drain_right.t7 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X11 source.t2 plus.t4 drain_left.t15 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X12 drain_right.t17 minus.t7 source.t30 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X13 source.t29 minus.t8 drain_right.t4 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X14 a_n2102_n1288# a_n2102_n1288# a_n2102_n1288# a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.3
X15 a_n2102_n1288# a_n2102_n1288# a_n2102_n1288# a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X16 drain_left.t14 plus.t5 source.t0 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X17 source.t17 plus.t6 drain_left.t13 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X18 drain_left.t12 plus.t7 source.t16 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X19 drain_right.t13 minus.t9 source.t28 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X20 a_n2102_n1288# a_n2102_n1288# a_n2102_n1288# a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X21 source.t27 minus.t10 drain_right.t0 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X22 source.t9 plus.t8 drain_left.t11 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X23 source.t26 minus.t11 drain_right.t5 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X24 source.t8 plus.t9 drain_left.t10 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X25 a_n2102_n1288# a_n2102_n1288# a_n2102_n1288# a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X26 source.t38 plus.t10 drain_left.t9 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X27 source.t25 minus.t12 drain_right.t18 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X28 drain_right.t14 minus.t13 source.t24 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X29 drain_left.t8 plus.t11 source.t39 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X30 drain_right.t19 minus.t14 source.t23 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X31 drain_right.t8 minus.t15 source.t22 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X32 drain_left.t7 plus.t12 source.t4 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X33 drain_left.t6 plus.t13 source.t6 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X34 source.t1 plus.t14 drain_left.t5 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X35 source.t21 minus.t16 drain_right.t9 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X36 source.t11 plus.t15 drain_left.t4 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X37 drain_left.t3 plus.t16 source.t14 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X38 drain_right.t10 minus.t17 source.t20 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X39 source.t19 minus.t18 drain_right.t6 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X40 source.t18 minus.t19 drain_right.t15 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X41 drain_left.t2 plus.t17 source.t5 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X42 source.t10 plus.t18 drain_left.t1 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X43 drain_left.t0 plus.t19 source.t13 a_n2102_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
R0 minus.n27 minus.t8 314.031
R1 minus.n7 minus.t13 314.031
R2 minus.n56 minus.t9 314.031
R3 minus.n35 minus.t0 314.031
R4 minus.n26 minus.t3 265.101
R5 minus.n24 minus.t19 265.101
R6 minus.n3 minus.t7 265.101
R7 minus.n18 minus.t1 265.101
R8 minus.n16 minus.t17 265.101
R9 minus.n4 minus.t11 265.101
R10 minus.n10 minus.t2 265.101
R11 minus.n6 minus.t18 265.101
R12 minus.n55 minus.t12 265.101
R13 minus.n53 minus.t5 265.101
R14 minus.n47 minus.t6 265.101
R15 minus.n46 minus.t14 265.101
R16 minus.n44 minus.t16 265.101
R17 minus.n32 minus.t4 265.101
R18 minus.n38 minus.t10 265.101
R19 minus.n34 minus.t15 265.101
R20 minus.n8 minus.n7 161.489
R21 minus.n36 minus.n35 161.489
R22 minus.n28 minus.n27 161.3
R23 minus.n25 minus.n0 161.3
R24 minus.n23 minus.n22 161.3
R25 minus.n21 minus.n1 161.3
R26 minus.n20 minus.n19 161.3
R27 minus.n17 minus.n2 161.3
R28 minus.n15 minus.n14 161.3
R29 minus.n13 minus.n12 161.3
R30 minus.n11 minus.n5 161.3
R31 minus.n9 minus.n8 161.3
R32 minus.n57 minus.n56 161.3
R33 minus.n54 minus.n29 161.3
R34 minus.n52 minus.n51 161.3
R35 minus.n50 minus.n30 161.3
R36 minus.n49 minus.n48 161.3
R37 minus.n45 minus.n31 161.3
R38 minus.n43 minus.n42 161.3
R39 minus.n41 minus.n40 161.3
R40 minus.n39 minus.n33 161.3
R41 minus.n37 minus.n36 161.3
R42 minus.n23 minus.n1 73.0308
R43 minus.n12 minus.n11 73.0308
R44 minus.n40 minus.n39 73.0308
R45 minus.n52 minus.n30 73.0308
R46 minus.n19 minus.n3 64.9975
R47 minus.n15 minus.n4 64.9975
R48 minus.n43 minus.n32 64.9975
R49 minus.n48 minus.n47 64.9975
R50 minus.n25 minus.n24 62.0763
R51 minus.n10 minus.n9 62.0763
R52 minus.n38 minus.n37 62.0763
R53 minus.n54 minus.n53 62.0763
R54 minus.n18 minus.n17 46.0096
R55 minus.n17 minus.n16 46.0096
R56 minus.n45 minus.n44 46.0096
R57 minus.n46 minus.n45 46.0096
R58 minus.n27 minus.n26 43.0884
R59 minus.n7 minus.n6 43.0884
R60 minus.n35 minus.n34 43.0884
R61 minus.n56 minus.n55 43.0884
R62 minus.n26 minus.n25 29.9429
R63 minus.n9 minus.n6 29.9429
R64 minus.n37 minus.n34 29.9429
R65 minus.n55 minus.n54 29.9429
R66 minus.n58 minus.n28 29.5232
R67 minus.n19 minus.n18 27.0217
R68 minus.n16 minus.n15 27.0217
R69 minus.n44 minus.n43 27.0217
R70 minus.n48 minus.n46 27.0217
R71 minus.n24 minus.n23 10.955
R72 minus.n11 minus.n10 10.955
R73 minus.n39 minus.n38 10.955
R74 minus.n53 minus.n52 10.955
R75 minus.n3 minus.n1 8.03383
R76 minus.n12 minus.n4 8.03383
R77 minus.n40 minus.n32 8.03383
R78 minus.n47 minus.n30 8.03383
R79 minus.n58 minus.n57 6.51565
R80 minus.n28 minus.n0 0.189894
R81 minus.n22 minus.n0 0.189894
R82 minus.n22 minus.n21 0.189894
R83 minus.n21 minus.n20 0.189894
R84 minus.n20 minus.n2 0.189894
R85 minus.n14 minus.n2 0.189894
R86 minus.n14 minus.n13 0.189894
R87 minus.n13 minus.n5 0.189894
R88 minus.n8 minus.n5 0.189894
R89 minus.n36 minus.n33 0.189894
R90 minus.n41 minus.n33 0.189894
R91 minus.n42 minus.n41 0.189894
R92 minus.n42 minus.n31 0.189894
R93 minus.n49 minus.n31 0.189894
R94 minus.n50 minus.n49 0.189894
R95 minus.n51 minus.n50 0.189894
R96 minus.n51 minus.n29 0.189894
R97 minus.n57 minus.n29 0.189894
R98 minus minus.n58 0.188
R99 drain_right.n10 drain_right.n8 101.338
R100 drain_right.n6 drain_right.n4 101.338
R101 drain_right.n2 drain_right.n0 101.338
R102 drain_right.n10 drain_right.n9 100.796
R103 drain_right.n12 drain_right.n11 100.796
R104 drain_right.n14 drain_right.n13 100.796
R105 drain_right.n16 drain_right.n15 100.796
R106 drain_right.n7 drain_right.n3 100.796
R107 drain_right.n6 drain_right.n5 100.796
R108 drain_right.n2 drain_right.n1 100.796
R109 drain_right drain_right.n7 23.5829
R110 drain_right.n3 drain_right.t9 9.9005
R111 drain_right.n3 drain_right.t19 9.9005
R112 drain_right.n4 drain_right.t18 9.9005
R113 drain_right.n4 drain_right.t13 9.9005
R114 drain_right.n5 drain_right.t7 9.9005
R115 drain_right.n5 drain_right.t3 9.9005
R116 drain_right.n1 drain_right.t0 9.9005
R117 drain_right.n1 drain_right.t12 9.9005
R118 drain_right.n0 drain_right.t11 9.9005
R119 drain_right.n0 drain_right.t8 9.9005
R120 drain_right.n8 drain_right.t6 9.9005
R121 drain_right.n8 drain_right.t14 9.9005
R122 drain_right.n9 drain_right.t5 9.9005
R123 drain_right.n9 drain_right.t2 9.9005
R124 drain_right.n11 drain_right.t1 9.9005
R125 drain_right.n11 drain_right.t10 9.9005
R126 drain_right.n13 drain_right.t15 9.9005
R127 drain_right.n13 drain_right.t17 9.9005
R128 drain_right.n15 drain_right.t4 9.9005
R129 drain_right.n15 drain_right.t16 9.9005
R130 drain_right drain_right.n16 6.19632
R131 drain_right.n16 drain_right.n14 0.543603
R132 drain_right.n14 drain_right.n12 0.543603
R133 drain_right.n12 drain_right.n10 0.543603
R134 drain_right.n7 drain_right.n6 0.488257
R135 drain_right.n7 drain_right.n2 0.488257
R136 source.n90 source.n88 289.615
R137 source.n74 source.n72 289.615
R138 source.n66 source.n64 289.615
R139 source.n50 source.n48 289.615
R140 source.n2 source.n0 289.615
R141 source.n18 source.n16 289.615
R142 source.n26 source.n24 289.615
R143 source.n42 source.n40 289.615
R144 source.n91 source.n90 185
R145 source.n75 source.n74 185
R146 source.n67 source.n66 185
R147 source.n51 source.n50 185
R148 source.n3 source.n2 185
R149 source.n19 source.n18 185
R150 source.n27 source.n26 185
R151 source.n43 source.n42 185
R152 source.t28 source.n89 167.117
R153 source.t37 source.n73 167.117
R154 source.t5 source.n65 167.117
R155 source.t2 source.n49 167.117
R156 source.t14 source.n1 167.117
R157 source.t7 source.n17 167.117
R158 source.t24 source.n25 167.117
R159 source.t29 source.n41 167.117
R160 source.n9 source.n8 84.1169
R161 source.n11 source.n10 84.1169
R162 source.n13 source.n12 84.1169
R163 source.n15 source.n14 84.1169
R164 source.n33 source.n32 84.1169
R165 source.n35 source.n34 84.1169
R166 source.n37 source.n36 84.1169
R167 source.n39 source.n38 84.1169
R168 source.n87 source.n86 84.1168
R169 source.n85 source.n84 84.1168
R170 source.n83 source.n82 84.1168
R171 source.n81 source.n80 84.1168
R172 source.n63 source.n62 84.1168
R173 source.n61 source.n60 84.1168
R174 source.n59 source.n58 84.1168
R175 source.n57 source.n56 84.1168
R176 source.n90 source.t28 52.3082
R177 source.n74 source.t37 52.3082
R178 source.n66 source.t5 52.3082
R179 source.n50 source.t2 52.3082
R180 source.n2 source.t14 52.3082
R181 source.n18 source.t7 52.3082
R182 source.n26 source.t24 52.3082
R183 source.n42 source.t29 52.3082
R184 source.n95 source.n94 31.4096
R185 source.n79 source.n78 31.4096
R186 source.n71 source.n70 31.4096
R187 source.n55 source.n54 31.4096
R188 source.n7 source.n6 31.4096
R189 source.n23 source.n22 31.4096
R190 source.n31 source.n30 31.4096
R191 source.n47 source.n46 31.4096
R192 source.n55 source.n47 14.2551
R193 source.n86 source.t32 9.9005
R194 source.n86 source.t25 9.9005
R195 source.n84 source.t23 9.9005
R196 source.n84 source.t31 9.9005
R197 source.n82 source.t33 9.9005
R198 source.n82 source.t21 9.9005
R199 source.n80 source.t22 9.9005
R200 source.n80 source.t27 9.9005
R201 source.n62 source.t0 9.9005
R202 source.n62 source.t9 9.9005
R203 source.n60 source.t4 9.9005
R204 source.n60 source.t12 9.9005
R205 source.n58 source.t3 9.9005
R206 source.n58 source.t8 9.9005
R207 source.n56 source.t6 9.9005
R208 source.n56 source.t11 9.9005
R209 source.n8 source.t15 9.9005
R210 source.n8 source.t38 9.9005
R211 source.n10 source.t39 9.9005
R212 source.n10 source.t10 9.9005
R213 source.n12 source.t13 9.9005
R214 source.n12 source.t17 9.9005
R215 source.n14 source.t16 9.9005
R216 source.n14 source.t1 9.9005
R217 source.n32 source.t35 9.9005
R218 source.n32 source.t19 9.9005
R219 source.n34 source.t20 9.9005
R220 source.n34 source.t26 9.9005
R221 source.n36 source.t30 9.9005
R222 source.n36 source.t36 9.9005
R223 source.n38 source.t34 9.9005
R224 source.n38 source.t18 9.9005
R225 source.n91 source.n89 9.71174
R226 source.n75 source.n73 9.71174
R227 source.n67 source.n65 9.71174
R228 source.n51 source.n49 9.71174
R229 source.n3 source.n1 9.71174
R230 source.n19 source.n17 9.71174
R231 source.n27 source.n25 9.71174
R232 source.n43 source.n41 9.71174
R233 source.n94 source.n93 9.45567
R234 source.n78 source.n77 9.45567
R235 source.n70 source.n69 9.45567
R236 source.n54 source.n53 9.45567
R237 source.n6 source.n5 9.45567
R238 source.n22 source.n21 9.45567
R239 source.n30 source.n29 9.45567
R240 source.n46 source.n45 9.45567
R241 source.n93 source.n92 9.3005
R242 source.n77 source.n76 9.3005
R243 source.n69 source.n68 9.3005
R244 source.n53 source.n52 9.3005
R245 source.n5 source.n4 9.3005
R246 source.n21 source.n20 9.3005
R247 source.n29 source.n28 9.3005
R248 source.n45 source.n44 9.3005
R249 source.n96 source.n7 8.72059
R250 source.n94 source.n88 8.14595
R251 source.n78 source.n72 8.14595
R252 source.n70 source.n64 8.14595
R253 source.n54 source.n48 8.14595
R254 source.n6 source.n0 8.14595
R255 source.n22 source.n16 8.14595
R256 source.n30 source.n24 8.14595
R257 source.n46 source.n40 8.14595
R258 source.n92 source.n91 7.3702
R259 source.n76 source.n75 7.3702
R260 source.n68 source.n67 7.3702
R261 source.n52 source.n51 7.3702
R262 source.n4 source.n3 7.3702
R263 source.n20 source.n19 7.3702
R264 source.n28 source.n27 7.3702
R265 source.n44 source.n43 7.3702
R266 source.n92 source.n88 5.81868
R267 source.n76 source.n72 5.81868
R268 source.n68 source.n64 5.81868
R269 source.n52 source.n48 5.81868
R270 source.n4 source.n0 5.81868
R271 source.n20 source.n16 5.81868
R272 source.n28 source.n24 5.81868
R273 source.n44 source.n40 5.81868
R274 source.n96 source.n95 5.53498
R275 source.n93 source.n89 3.44771
R276 source.n77 source.n73 3.44771
R277 source.n69 source.n65 3.44771
R278 source.n53 source.n49 3.44771
R279 source.n5 source.n1 3.44771
R280 source.n21 source.n17 3.44771
R281 source.n29 source.n25 3.44771
R282 source.n45 source.n41 3.44771
R283 source.n47 source.n39 0.543603
R284 source.n39 source.n37 0.543603
R285 source.n37 source.n35 0.543603
R286 source.n35 source.n33 0.543603
R287 source.n33 source.n31 0.543603
R288 source.n23 source.n15 0.543603
R289 source.n15 source.n13 0.543603
R290 source.n13 source.n11 0.543603
R291 source.n11 source.n9 0.543603
R292 source.n9 source.n7 0.543603
R293 source.n57 source.n55 0.543603
R294 source.n59 source.n57 0.543603
R295 source.n61 source.n59 0.543603
R296 source.n63 source.n61 0.543603
R297 source.n71 source.n63 0.543603
R298 source.n81 source.n79 0.543603
R299 source.n83 source.n81 0.543603
R300 source.n85 source.n83 0.543603
R301 source.n87 source.n85 0.543603
R302 source.n95 source.n87 0.543603
R303 source.n31 source.n23 0.470328
R304 source.n79 source.n71 0.470328
R305 source source.n96 0.188
R306 plus.n6 plus.t3 314.031
R307 plus.n27 plus.t16 314.031
R308 plus.n36 plus.t17 314.031
R309 plus.n56 plus.t4 314.031
R310 plus.n5 plus.t7 265.101
R311 plus.n9 plus.t14 265.101
R312 plus.n3 plus.t19 265.101
R313 plus.n15 plus.t6 265.101
R314 plus.n17 plus.t11 265.101
R315 plus.n18 plus.t18 265.101
R316 plus.n24 plus.t1 265.101
R317 plus.n26 plus.t10 265.101
R318 plus.n35 plus.t8 265.101
R319 plus.n39 plus.t5 265.101
R320 plus.n33 plus.t0 265.101
R321 plus.n45 plus.t12 265.101
R322 plus.n47 plus.t9 265.101
R323 plus.n32 plus.t2 265.101
R324 plus.n53 plus.t15 265.101
R325 plus.n55 plus.t13 265.101
R326 plus.n7 plus.n6 161.489
R327 plus.n37 plus.n36 161.489
R328 plus.n8 plus.n7 161.3
R329 plus.n10 plus.n4 161.3
R330 plus.n12 plus.n11 161.3
R331 plus.n14 plus.n13 161.3
R332 plus.n16 plus.n2 161.3
R333 plus.n20 plus.n19 161.3
R334 plus.n21 plus.n1 161.3
R335 plus.n23 plus.n22 161.3
R336 plus.n25 plus.n0 161.3
R337 plus.n28 plus.n27 161.3
R338 plus.n38 plus.n37 161.3
R339 plus.n40 plus.n34 161.3
R340 plus.n42 plus.n41 161.3
R341 plus.n44 plus.n43 161.3
R342 plus.n46 plus.n31 161.3
R343 plus.n49 plus.n48 161.3
R344 plus.n50 plus.n30 161.3
R345 plus.n52 plus.n51 161.3
R346 plus.n54 plus.n29 161.3
R347 plus.n57 plus.n56 161.3
R348 plus.n11 plus.n10 73.0308
R349 plus.n23 plus.n1 73.0308
R350 plus.n52 plus.n30 73.0308
R351 plus.n41 plus.n40 73.0308
R352 plus.n14 plus.n3 64.9975
R353 plus.n19 plus.n18 64.9975
R354 plus.n48 plus.n32 64.9975
R355 plus.n44 plus.n33 64.9975
R356 plus.n9 plus.n8 62.0763
R357 plus.n25 plus.n24 62.0763
R358 plus.n54 plus.n53 62.0763
R359 plus.n39 plus.n38 62.0763
R360 plus.n16 plus.n15 46.0096
R361 plus.n17 plus.n16 46.0096
R362 plus.n47 plus.n46 46.0096
R363 plus.n46 plus.n45 46.0096
R364 plus.n6 plus.n5 43.0884
R365 plus.n27 plus.n26 43.0884
R366 plus.n56 plus.n55 43.0884
R367 plus.n36 plus.n35 43.0884
R368 plus.n8 plus.n5 29.9429
R369 plus.n26 plus.n25 29.9429
R370 plus.n55 plus.n54 29.9429
R371 plus.n38 plus.n35 29.9429
R372 plus plus.n57 27.1922
R373 plus.n15 plus.n14 27.0217
R374 plus.n19 plus.n17 27.0217
R375 plus.n48 plus.n47 27.0217
R376 plus.n45 plus.n44 27.0217
R377 plus.n10 plus.n9 10.955
R378 plus.n24 plus.n23 10.955
R379 plus.n53 plus.n52 10.955
R380 plus.n40 plus.n39 10.955
R381 plus plus.n28 8.37171
R382 plus.n11 plus.n3 8.03383
R383 plus.n18 plus.n1 8.03383
R384 plus.n32 plus.n30 8.03383
R385 plus.n41 plus.n33 8.03383
R386 plus.n7 plus.n4 0.189894
R387 plus.n12 plus.n4 0.189894
R388 plus.n13 plus.n12 0.189894
R389 plus.n13 plus.n2 0.189894
R390 plus.n20 plus.n2 0.189894
R391 plus.n21 plus.n20 0.189894
R392 plus.n22 plus.n21 0.189894
R393 plus.n22 plus.n0 0.189894
R394 plus.n28 plus.n0 0.189894
R395 plus.n57 plus.n29 0.189894
R396 plus.n51 plus.n29 0.189894
R397 plus.n51 plus.n50 0.189894
R398 plus.n50 plus.n49 0.189894
R399 plus.n49 plus.n31 0.189894
R400 plus.n43 plus.n31 0.189894
R401 plus.n43 plus.n42 0.189894
R402 plus.n42 plus.n34 0.189894
R403 plus.n37 plus.n34 0.189894
R404 drain_left.n10 drain_left.n8 101.338
R405 drain_left.n6 drain_left.n4 101.338
R406 drain_left.n2 drain_left.n0 101.338
R407 drain_left.n16 drain_left.n15 100.796
R408 drain_left.n14 drain_left.n13 100.796
R409 drain_left.n12 drain_left.n11 100.796
R410 drain_left.n10 drain_left.n9 100.796
R411 drain_left.n7 drain_left.n3 100.796
R412 drain_left.n6 drain_left.n5 100.796
R413 drain_left.n2 drain_left.n1 100.796
R414 drain_left drain_left.n7 24.1361
R415 drain_left.n3 drain_left.t10 9.9005
R416 drain_left.n3 drain_left.t7 9.9005
R417 drain_left.n4 drain_left.t11 9.9005
R418 drain_left.n4 drain_left.t2 9.9005
R419 drain_left.n5 drain_left.t19 9.9005
R420 drain_left.n5 drain_left.t14 9.9005
R421 drain_left.n1 drain_left.t4 9.9005
R422 drain_left.n1 drain_left.t17 9.9005
R423 drain_left.n0 drain_left.t15 9.9005
R424 drain_left.n0 drain_left.t6 9.9005
R425 drain_left.n15 drain_left.t9 9.9005
R426 drain_left.n15 drain_left.t3 9.9005
R427 drain_left.n13 drain_left.t1 9.9005
R428 drain_left.n13 drain_left.t18 9.9005
R429 drain_left.n11 drain_left.t13 9.9005
R430 drain_left.n11 drain_left.t8 9.9005
R431 drain_left.n9 drain_left.t5 9.9005
R432 drain_left.n9 drain_left.t0 9.9005
R433 drain_left.n8 drain_left.t16 9.9005
R434 drain_left.n8 drain_left.t12 9.9005
R435 drain_left drain_left.n16 6.19632
R436 drain_left.n12 drain_left.n10 0.543603
R437 drain_left.n14 drain_left.n12 0.543603
R438 drain_left.n16 drain_left.n14 0.543603
R439 drain_left.n7 drain_left.n6 0.488257
R440 drain_left.n7 drain_left.n2 0.488257
C0 drain_right minus 1.70016f
C1 drain_left plus 1.90608f
C2 source drain_left 9.0008f
C3 minus plus 3.93063f
C4 source minus 1.97467f
C5 drain_right plus 0.367499f
C6 drain_left minus 0.177738f
C7 source drain_right 9.001241f
C8 drain_left drain_right 1.10857f
C9 source plus 1.98863f
C10 drain_right a_n2102_n1288# 4.30942f
C11 drain_left a_n2102_n1288# 4.59561f
C12 source a_n2102_n1288# 3.228544f
C13 minus a_n2102_n1288# 7.431102f
C14 plus a_n2102_n1288# 8.015919f
C15 drain_left.t15 a_n2102_n1288# 0.041867f
C16 drain_left.t6 a_n2102_n1288# 0.041867f
C17 drain_left.n0 a_n2102_n1288# 0.26466f
C18 drain_left.t4 a_n2102_n1288# 0.041867f
C19 drain_left.t17 a_n2102_n1288# 0.041867f
C20 drain_left.n1 a_n2102_n1288# 0.263019f
C21 drain_left.n2 a_n2102_n1288# 0.596501f
C22 drain_left.t10 a_n2102_n1288# 0.041867f
C23 drain_left.t7 a_n2102_n1288# 0.041867f
C24 drain_left.n3 a_n2102_n1288# 0.263019f
C25 drain_left.t11 a_n2102_n1288# 0.041867f
C26 drain_left.t2 a_n2102_n1288# 0.041867f
C27 drain_left.n4 a_n2102_n1288# 0.26466f
C28 drain_left.t19 a_n2102_n1288# 0.041867f
C29 drain_left.t14 a_n2102_n1288# 0.041867f
C30 drain_left.n5 a_n2102_n1288# 0.263019f
C31 drain_left.n6 a_n2102_n1288# 0.596501f
C32 drain_left.n7 a_n2102_n1288# 1.07488f
C33 drain_left.t16 a_n2102_n1288# 0.041867f
C34 drain_left.t12 a_n2102_n1288# 0.041867f
C35 drain_left.n8 a_n2102_n1288# 0.264661f
C36 drain_left.t5 a_n2102_n1288# 0.041867f
C37 drain_left.t0 a_n2102_n1288# 0.041867f
C38 drain_left.n9 a_n2102_n1288# 0.26302f
C39 drain_left.n10 a_n2102_n1288# 0.599964f
C40 drain_left.t13 a_n2102_n1288# 0.041867f
C41 drain_left.t8 a_n2102_n1288# 0.041867f
C42 drain_left.n11 a_n2102_n1288# 0.26302f
C43 drain_left.n12 a_n2102_n1288# 0.295468f
C44 drain_left.t1 a_n2102_n1288# 0.041867f
C45 drain_left.t18 a_n2102_n1288# 0.041867f
C46 drain_left.n13 a_n2102_n1288# 0.26302f
C47 drain_left.n14 a_n2102_n1288# 0.295468f
C48 drain_left.t9 a_n2102_n1288# 0.041867f
C49 drain_left.t3 a_n2102_n1288# 0.041867f
C50 drain_left.n15 a_n2102_n1288# 0.26302f
C51 drain_left.n16 a_n2102_n1288# 0.515961f
C52 plus.n0 a_n2102_n1288# 0.025759f
C53 plus.t10 a_n2102_n1288# 0.045479f
C54 plus.t1 a_n2102_n1288# 0.045479f
C55 plus.n1 a_n2102_n1288# 0.009419f
C56 plus.n2 a_n2102_n1288# 0.025759f
C57 plus.t11 a_n2102_n1288# 0.045479f
C58 plus.t6 a_n2102_n1288# 0.045479f
C59 plus.t19 a_n2102_n1288# 0.045479f
C60 plus.n3 a_n2102_n1288# 0.031763f
C61 plus.n4 a_n2102_n1288# 0.025759f
C62 plus.t14 a_n2102_n1288# 0.045479f
C63 plus.t7 a_n2102_n1288# 0.045479f
C64 plus.n5 a_n2102_n1288# 0.031763f
C65 plus.t3 a_n2102_n1288# 0.050762f
C66 plus.n6 a_n2102_n1288# 0.039272f
C67 plus.n7 a_n2102_n1288# 0.058943f
C68 plus.n8 a_n2102_n1288# 0.01061f
C69 plus.n9 a_n2102_n1288# 0.031763f
C70 plus.n10 a_n2102_n1288# 0.009736f
C71 plus.n11 a_n2102_n1288# 0.009419f
C72 plus.n12 a_n2102_n1288# 0.025759f
C73 plus.n13 a_n2102_n1288# 0.025759f
C74 plus.n14 a_n2102_n1288# 0.01061f
C75 plus.n15 a_n2102_n1288# 0.031763f
C76 plus.n16 a_n2102_n1288# 0.01061f
C77 plus.n17 a_n2102_n1288# 0.031763f
C78 plus.t18 a_n2102_n1288# 0.045479f
C79 plus.n18 a_n2102_n1288# 0.031763f
C80 plus.n19 a_n2102_n1288# 0.01061f
C81 plus.n20 a_n2102_n1288# 0.025759f
C82 plus.n21 a_n2102_n1288# 0.025759f
C83 plus.n22 a_n2102_n1288# 0.025759f
C84 plus.n23 a_n2102_n1288# 0.009736f
C85 plus.n24 a_n2102_n1288# 0.031763f
C86 plus.n25 a_n2102_n1288# 0.01061f
C87 plus.n26 a_n2102_n1288# 0.031763f
C88 plus.t16 a_n2102_n1288# 0.050762f
C89 plus.n27 a_n2102_n1288# 0.039233f
C90 plus.n28 a_n2102_n1288# 0.185147f
C91 plus.n29 a_n2102_n1288# 0.025759f
C92 plus.t4 a_n2102_n1288# 0.050762f
C93 plus.t13 a_n2102_n1288# 0.045479f
C94 plus.t15 a_n2102_n1288# 0.045479f
C95 plus.n30 a_n2102_n1288# 0.009419f
C96 plus.n31 a_n2102_n1288# 0.025759f
C97 plus.t2 a_n2102_n1288# 0.045479f
C98 plus.n32 a_n2102_n1288# 0.031763f
C99 plus.t9 a_n2102_n1288# 0.045479f
C100 plus.t12 a_n2102_n1288# 0.045479f
C101 plus.t0 a_n2102_n1288# 0.045479f
C102 plus.n33 a_n2102_n1288# 0.031763f
C103 plus.n34 a_n2102_n1288# 0.025759f
C104 plus.t5 a_n2102_n1288# 0.045479f
C105 plus.t8 a_n2102_n1288# 0.045479f
C106 plus.n35 a_n2102_n1288# 0.031763f
C107 plus.t17 a_n2102_n1288# 0.050762f
C108 plus.n36 a_n2102_n1288# 0.039272f
C109 plus.n37 a_n2102_n1288# 0.058943f
C110 plus.n38 a_n2102_n1288# 0.01061f
C111 plus.n39 a_n2102_n1288# 0.031763f
C112 plus.n40 a_n2102_n1288# 0.009736f
C113 plus.n41 a_n2102_n1288# 0.009419f
C114 plus.n42 a_n2102_n1288# 0.025759f
C115 plus.n43 a_n2102_n1288# 0.025759f
C116 plus.n44 a_n2102_n1288# 0.01061f
C117 plus.n45 a_n2102_n1288# 0.031763f
C118 plus.n46 a_n2102_n1288# 0.01061f
C119 plus.n47 a_n2102_n1288# 0.031763f
C120 plus.n48 a_n2102_n1288# 0.01061f
C121 plus.n49 a_n2102_n1288# 0.025759f
C122 plus.n50 a_n2102_n1288# 0.025759f
C123 plus.n51 a_n2102_n1288# 0.025759f
C124 plus.n52 a_n2102_n1288# 0.009736f
C125 plus.n53 a_n2102_n1288# 0.031763f
C126 plus.n54 a_n2102_n1288# 0.01061f
C127 plus.n55 a_n2102_n1288# 0.031763f
C128 plus.n56 a_n2102_n1288# 0.039233f
C129 plus.n57 a_n2102_n1288# 0.621654f
C130 source.n0 a_n2102_n1288# 0.041033f
C131 source.n1 a_n2102_n1288# 0.090791f
C132 source.t14 a_n2102_n1288# 0.068134f
C133 source.n2 a_n2102_n1288# 0.071056f
C134 source.n3 a_n2102_n1288# 0.022906f
C135 source.n4 a_n2102_n1288# 0.015107f
C136 source.n5 a_n2102_n1288# 0.200125f
C137 source.n6 a_n2102_n1288# 0.044982f
C138 source.n7 a_n2102_n1288# 0.424464f
C139 source.t15 a_n2102_n1288# 0.044432f
C140 source.t38 a_n2102_n1288# 0.044432f
C141 source.n8 a_n2102_n1288# 0.237532f
C142 source.n9 a_n2102_n1288# 0.316964f
C143 source.t39 a_n2102_n1288# 0.044432f
C144 source.t10 a_n2102_n1288# 0.044432f
C145 source.n10 a_n2102_n1288# 0.237532f
C146 source.n11 a_n2102_n1288# 0.316964f
C147 source.t13 a_n2102_n1288# 0.044432f
C148 source.t17 a_n2102_n1288# 0.044432f
C149 source.n12 a_n2102_n1288# 0.237532f
C150 source.n13 a_n2102_n1288# 0.316964f
C151 source.t16 a_n2102_n1288# 0.044432f
C152 source.t1 a_n2102_n1288# 0.044432f
C153 source.n14 a_n2102_n1288# 0.237532f
C154 source.n15 a_n2102_n1288# 0.316964f
C155 source.n16 a_n2102_n1288# 0.041033f
C156 source.n17 a_n2102_n1288# 0.090791f
C157 source.t7 a_n2102_n1288# 0.068134f
C158 source.n18 a_n2102_n1288# 0.071056f
C159 source.n19 a_n2102_n1288# 0.022906f
C160 source.n20 a_n2102_n1288# 0.015107f
C161 source.n21 a_n2102_n1288# 0.200125f
C162 source.n22 a_n2102_n1288# 0.044982f
C163 source.n23 a_n2102_n1288# 0.114903f
C164 source.n24 a_n2102_n1288# 0.041033f
C165 source.n25 a_n2102_n1288# 0.090791f
C166 source.t24 a_n2102_n1288# 0.068134f
C167 source.n26 a_n2102_n1288# 0.071056f
C168 source.n27 a_n2102_n1288# 0.022906f
C169 source.n28 a_n2102_n1288# 0.015107f
C170 source.n29 a_n2102_n1288# 0.200125f
C171 source.n30 a_n2102_n1288# 0.044982f
C172 source.n31 a_n2102_n1288# 0.114903f
C173 source.t35 a_n2102_n1288# 0.044432f
C174 source.t19 a_n2102_n1288# 0.044432f
C175 source.n32 a_n2102_n1288# 0.237532f
C176 source.n33 a_n2102_n1288# 0.316964f
C177 source.t20 a_n2102_n1288# 0.044432f
C178 source.t26 a_n2102_n1288# 0.044432f
C179 source.n34 a_n2102_n1288# 0.237532f
C180 source.n35 a_n2102_n1288# 0.316964f
C181 source.t30 a_n2102_n1288# 0.044432f
C182 source.t36 a_n2102_n1288# 0.044432f
C183 source.n36 a_n2102_n1288# 0.237532f
C184 source.n37 a_n2102_n1288# 0.316964f
C185 source.t34 a_n2102_n1288# 0.044432f
C186 source.t18 a_n2102_n1288# 0.044432f
C187 source.n38 a_n2102_n1288# 0.237532f
C188 source.n39 a_n2102_n1288# 0.316964f
C189 source.n40 a_n2102_n1288# 0.041033f
C190 source.n41 a_n2102_n1288# 0.090791f
C191 source.t29 a_n2102_n1288# 0.068134f
C192 source.n42 a_n2102_n1288# 0.071056f
C193 source.n43 a_n2102_n1288# 0.022906f
C194 source.n44 a_n2102_n1288# 0.015107f
C195 source.n45 a_n2102_n1288# 0.200125f
C196 source.n46 a_n2102_n1288# 0.044982f
C197 source.n47 a_n2102_n1288# 0.686565f
C198 source.n48 a_n2102_n1288# 0.041033f
C199 source.n49 a_n2102_n1288# 0.090791f
C200 source.t2 a_n2102_n1288# 0.068134f
C201 source.n50 a_n2102_n1288# 0.071056f
C202 source.n51 a_n2102_n1288# 0.022906f
C203 source.n52 a_n2102_n1288# 0.015107f
C204 source.n53 a_n2102_n1288# 0.200125f
C205 source.n54 a_n2102_n1288# 0.044982f
C206 source.n55 a_n2102_n1288# 0.686565f
C207 source.t6 a_n2102_n1288# 0.044432f
C208 source.t11 a_n2102_n1288# 0.044432f
C209 source.n56 a_n2102_n1288# 0.23753f
C210 source.n57 a_n2102_n1288# 0.316965f
C211 source.t3 a_n2102_n1288# 0.044432f
C212 source.t8 a_n2102_n1288# 0.044432f
C213 source.n58 a_n2102_n1288# 0.23753f
C214 source.n59 a_n2102_n1288# 0.316965f
C215 source.t4 a_n2102_n1288# 0.044432f
C216 source.t12 a_n2102_n1288# 0.044432f
C217 source.n60 a_n2102_n1288# 0.23753f
C218 source.n61 a_n2102_n1288# 0.316965f
C219 source.t0 a_n2102_n1288# 0.044432f
C220 source.t9 a_n2102_n1288# 0.044432f
C221 source.n62 a_n2102_n1288# 0.23753f
C222 source.n63 a_n2102_n1288# 0.316965f
C223 source.n64 a_n2102_n1288# 0.041033f
C224 source.n65 a_n2102_n1288# 0.090791f
C225 source.t5 a_n2102_n1288# 0.068134f
C226 source.n66 a_n2102_n1288# 0.071056f
C227 source.n67 a_n2102_n1288# 0.022906f
C228 source.n68 a_n2102_n1288# 0.015107f
C229 source.n69 a_n2102_n1288# 0.200125f
C230 source.n70 a_n2102_n1288# 0.044982f
C231 source.n71 a_n2102_n1288# 0.114903f
C232 source.n72 a_n2102_n1288# 0.041033f
C233 source.n73 a_n2102_n1288# 0.090791f
C234 source.t37 a_n2102_n1288# 0.068134f
C235 source.n74 a_n2102_n1288# 0.071056f
C236 source.n75 a_n2102_n1288# 0.022906f
C237 source.n76 a_n2102_n1288# 0.015107f
C238 source.n77 a_n2102_n1288# 0.200125f
C239 source.n78 a_n2102_n1288# 0.044982f
C240 source.n79 a_n2102_n1288# 0.114903f
C241 source.t22 a_n2102_n1288# 0.044432f
C242 source.t27 a_n2102_n1288# 0.044432f
C243 source.n80 a_n2102_n1288# 0.23753f
C244 source.n81 a_n2102_n1288# 0.316965f
C245 source.t33 a_n2102_n1288# 0.044432f
C246 source.t21 a_n2102_n1288# 0.044432f
C247 source.n82 a_n2102_n1288# 0.23753f
C248 source.n83 a_n2102_n1288# 0.316965f
C249 source.t23 a_n2102_n1288# 0.044432f
C250 source.t31 a_n2102_n1288# 0.044432f
C251 source.n84 a_n2102_n1288# 0.23753f
C252 source.n85 a_n2102_n1288# 0.316965f
C253 source.t32 a_n2102_n1288# 0.044432f
C254 source.t25 a_n2102_n1288# 0.044432f
C255 source.n86 a_n2102_n1288# 0.23753f
C256 source.n87 a_n2102_n1288# 0.316965f
C257 source.n88 a_n2102_n1288# 0.041033f
C258 source.n89 a_n2102_n1288# 0.090791f
C259 source.t28 a_n2102_n1288# 0.068134f
C260 source.n90 a_n2102_n1288# 0.071056f
C261 source.n91 a_n2102_n1288# 0.022906f
C262 source.n92 a_n2102_n1288# 0.015107f
C263 source.n93 a_n2102_n1288# 0.200125f
C264 source.n94 a_n2102_n1288# 0.044982f
C265 source.n95 a_n2102_n1288# 0.273601f
C266 source.n96 a_n2102_n1288# 0.69506f
C267 drain_right.t11 a_n2102_n1288# 0.042354f
C268 drain_right.t8 a_n2102_n1288# 0.042354f
C269 drain_right.n0 a_n2102_n1288# 0.267742f
C270 drain_right.t0 a_n2102_n1288# 0.042354f
C271 drain_right.t12 a_n2102_n1288# 0.042354f
C272 drain_right.n1 a_n2102_n1288# 0.266083f
C273 drain_right.n2 a_n2102_n1288# 0.60345f
C274 drain_right.t9 a_n2102_n1288# 0.042354f
C275 drain_right.t19 a_n2102_n1288# 0.042354f
C276 drain_right.n3 a_n2102_n1288# 0.266083f
C277 drain_right.t18 a_n2102_n1288# 0.042354f
C278 drain_right.t13 a_n2102_n1288# 0.042354f
C279 drain_right.n4 a_n2102_n1288# 0.267742f
C280 drain_right.t7 a_n2102_n1288# 0.042354f
C281 drain_right.t3 a_n2102_n1288# 0.042354f
C282 drain_right.n5 a_n2102_n1288# 0.266083f
C283 drain_right.n6 a_n2102_n1288# 0.60345f
C284 drain_right.n7 a_n2102_n1288# 1.03504f
C285 drain_right.t6 a_n2102_n1288# 0.042354f
C286 drain_right.t14 a_n2102_n1288# 0.042354f
C287 drain_right.n8 a_n2102_n1288# 0.267744f
C288 drain_right.t5 a_n2102_n1288# 0.042354f
C289 drain_right.t2 a_n2102_n1288# 0.042354f
C290 drain_right.n9 a_n2102_n1288# 0.266084f
C291 drain_right.n10 a_n2102_n1288# 0.606953f
C292 drain_right.t1 a_n2102_n1288# 0.042354f
C293 drain_right.t10 a_n2102_n1288# 0.042354f
C294 drain_right.n11 a_n2102_n1288# 0.266084f
C295 drain_right.n12 a_n2102_n1288# 0.298909f
C296 drain_right.t15 a_n2102_n1288# 0.042354f
C297 drain_right.t17 a_n2102_n1288# 0.042354f
C298 drain_right.n13 a_n2102_n1288# 0.266084f
C299 drain_right.n14 a_n2102_n1288# 0.298909f
C300 drain_right.t4 a_n2102_n1288# 0.042354f
C301 drain_right.t16 a_n2102_n1288# 0.042354f
C302 drain_right.n15 a_n2102_n1288# 0.266084f
C303 drain_right.n16 a_n2102_n1288# 0.521971f
C304 minus.n0 a_n2102_n1288# 0.025419f
C305 minus.t8 a_n2102_n1288# 0.050093f
C306 minus.t3 a_n2102_n1288# 0.044879f
C307 minus.t19 a_n2102_n1288# 0.044879f
C308 minus.n1 a_n2102_n1288# 0.009294f
C309 minus.n2 a_n2102_n1288# 0.025419f
C310 minus.t7 a_n2102_n1288# 0.044879f
C311 minus.n3 a_n2102_n1288# 0.031344f
C312 minus.t1 a_n2102_n1288# 0.044879f
C313 minus.t17 a_n2102_n1288# 0.044879f
C314 minus.t11 a_n2102_n1288# 0.044879f
C315 minus.n4 a_n2102_n1288# 0.031344f
C316 minus.n5 a_n2102_n1288# 0.025419f
C317 minus.t2 a_n2102_n1288# 0.044879f
C318 minus.t18 a_n2102_n1288# 0.044879f
C319 minus.n6 a_n2102_n1288# 0.031344f
C320 minus.t13 a_n2102_n1288# 0.050093f
C321 minus.n7 a_n2102_n1288# 0.038755f
C322 minus.n8 a_n2102_n1288# 0.058166f
C323 minus.n9 a_n2102_n1288# 0.01047f
C324 minus.n10 a_n2102_n1288# 0.031344f
C325 minus.n11 a_n2102_n1288# 0.009608f
C326 minus.n12 a_n2102_n1288# 0.009294f
C327 minus.n13 a_n2102_n1288# 0.025419f
C328 minus.n14 a_n2102_n1288# 0.025419f
C329 minus.n15 a_n2102_n1288# 0.01047f
C330 minus.n16 a_n2102_n1288# 0.031344f
C331 minus.n17 a_n2102_n1288# 0.01047f
C332 minus.n18 a_n2102_n1288# 0.031344f
C333 minus.n19 a_n2102_n1288# 0.01047f
C334 minus.n20 a_n2102_n1288# 0.025419f
C335 minus.n21 a_n2102_n1288# 0.025419f
C336 minus.n22 a_n2102_n1288# 0.025419f
C337 minus.n23 a_n2102_n1288# 0.009608f
C338 minus.n24 a_n2102_n1288# 0.031344f
C339 minus.n25 a_n2102_n1288# 0.01047f
C340 minus.n26 a_n2102_n1288# 0.031344f
C341 minus.n27 a_n2102_n1288# 0.038716f
C342 minus.n28 a_n2102_n1288# 0.643723f
C343 minus.n29 a_n2102_n1288# 0.025419f
C344 minus.t12 a_n2102_n1288# 0.044879f
C345 minus.t5 a_n2102_n1288# 0.044879f
C346 minus.n30 a_n2102_n1288# 0.009294f
C347 minus.n31 a_n2102_n1288# 0.025419f
C348 minus.t14 a_n2102_n1288# 0.044879f
C349 minus.t16 a_n2102_n1288# 0.044879f
C350 minus.t4 a_n2102_n1288# 0.044879f
C351 minus.n32 a_n2102_n1288# 0.031344f
C352 minus.n33 a_n2102_n1288# 0.025419f
C353 minus.t10 a_n2102_n1288# 0.044879f
C354 minus.t15 a_n2102_n1288# 0.044879f
C355 minus.n34 a_n2102_n1288# 0.031344f
C356 minus.t0 a_n2102_n1288# 0.050093f
C357 minus.n35 a_n2102_n1288# 0.038755f
C358 minus.n36 a_n2102_n1288# 0.058166f
C359 minus.n37 a_n2102_n1288# 0.01047f
C360 minus.n38 a_n2102_n1288# 0.031344f
C361 minus.n39 a_n2102_n1288# 0.009608f
C362 minus.n40 a_n2102_n1288# 0.009294f
C363 minus.n41 a_n2102_n1288# 0.025419f
C364 minus.n42 a_n2102_n1288# 0.025419f
C365 minus.n43 a_n2102_n1288# 0.01047f
C366 minus.n44 a_n2102_n1288# 0.031344f
C367 minus.n45 a_n2102_n1288# 0.01047f
C368 minus.n46 a_n2102_n1288# 0.031344f
C369 minus.t6 a_n2102_n1288# 0.044879f
C370 minus.n47 a_n2102_n1288# 0.031344f
C371 minus.n48 a_n2102_n1288# 0.01047f
C372 minus.n49 a_n2102_n1288# 0.025419f
C373 minus.n50 a_n2102_n1288# 0.025419f
C374 minus.n51 a_n2102_n1288# 0.025419f
C375 minus.n52 a_n2102_n1288# 0.009608f
C376 minus.n53 a_n2102_n1288# 0.031344f
C377 minus.n54 a_n2102_n1288# 0.01047f
C378 minus.n55 a_n2102_n1288# 0.031344f
C379 minus.t9 a_n2102_n1288# 0.050093f
C380 minus.n56 a_n2102_n1288# 0.038716f
C381 minus.n57 a_n2102_n1288# 0.167121f
C382 minus.n58 a_n2102_n1288# 0.794233f
.ends

