* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right.t13 minus.t0 source.t21 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X1 drain_right.t12 minus.t1 source.t24 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.2
X2 source.t12 minus.t2 drain_right.t11 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X3 drain_right.t10 minus.t3 source.t22 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X4 drain_left.t13 plus.t0 source.t8 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X5 drain_left.t12 plus.t1 source.t10 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.2
X6 source.t7 plus.t2 drain_left.t11 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X7 a_n1564_n1088# a_n1564_n1088# a_n1564_n1088# a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.2
X8 a_n1564_n1088# a_n1564_n1088# a_n1564_n1088# a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.2
X9 source.t15 minus.t4 drain_right.t9 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X10 drain_right.t8 minus.t5 source.t13 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.2
X11 source.t11 minus.t6 drain_right.t7 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X12 source.t14 minus.t7 drain_right.t6 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X13 source.t25 plus.t3 drain_left.t10 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X14 a_n1564_n1088# a_n1564_n1088# a_n1564_n1088# a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.2
X15 source.t26 plus.t4 drain_left.t9 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X16 drain_left.t8 plus.t5 source.t27 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.2
X17 drain_right.t5 minus.t8 source.t20 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.2
X18 drain_left.t7 plus.t6 source.t4 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.2
X19 drain_right.t4 minus.t9 source.t18 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.2
X20 drain_right.t3 minus.t10 source.t17 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X21 drain_left.t6 plus.t7 source.t3 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.2
X22 drain_right.t2 minus.t11 source.t23 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X23 a_n1564_n1088# a_n1564_n1088# a_n1564_n1088# a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.2
X24 source.t16 minus.t12 drain_right.t1 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X25 source.t6 plus.t8 drain_left.t5 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X26 drain_left.t4 plus.t9 source.t9 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X27 source.t1 plus.t10 drain_left.t3 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X28 source.t5 plus.t11 drain_left.t2 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X29 source.t19 minus.t13 drain_right.t0 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X30 drain_left.t1 plus.t12 source.t0 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X31 drain_left.t0 plus.t13 source.t2 a_n1564_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
R0 minus.n14 minus.t1 326.812
R1 minus.n3 minus.t9 326.812
R2 minus.n30 minus.t5 326.812
R3 minus.n19 minus.t8 326.812
R4 minus.n13 minus.t4 277.151
R5 minus.n11 minus.t10 277.151
R6 minus.n1 minus.t13 277.151
R7 minus.n6 minus.t0 277.151
R8 minus.n4 minus.t6 277.151
R9 minus.n29 minus.t2 277.151
R10 minus.n27 minus.t11 277.151
R11 minus.n17 minus.t7 277.151
R12 minus.n22 minus.t3 277.151
R13 minus.n20 minus.t12 277.151
R14 minus.n3 minus.n2 161.489
R15 minus.n19 minus.n18 161.489
R16 minus.n15 minus.n14 161.3
R17 minus.n12 minus.n0 161.3
R18 minus.n10 minus.n9 161.3
R19 minus.n8 minus.n7 161.3
R20 minus.n5 minus.n2 161.3
R21 minus.n31 minus.n30 161.3
R22 minus.n28 minus.n16 161.3
R23 minus.n26 minus.n25 161.3
R24 minus.n24 minus.n23 161.3
R25 minus.n21 minus.n18 161.3
R26 minus.n13 minus.n12 45.2793
R27 minus.n5 minus.n4 45.2793
R28 minus.n21 minus.n20 45.2793
R29 minus.n29 minus.n28 45.2793
R30 minus.n11 minus.n10 40.8975
R31 minus.n7 minus.n6 40.8975
R32 minus.n23 minus.n22 40.8975
R33 minus.n27 minus.n26 40.8975
R34 minus.n10 minus.n1 36.5157
R35 minus.n7 minus.n1 36.5157
R36 minus.n23 minus.n17 36.5157
R37 minus.n26 minus.n17 36.5157
R38 minus.n12 minus.n11 32.1338
R39 minus.n6 minus.n5 32.1338
R40 minus.n22 minus.n21 32.1338
R41 minus.n28 minus.n27 32.1338
R42 minus.n14 minus.n13 27.752
R43 minus.n4 minus.n3 27.752
R44 minus.n20 minus.n19 27.752
R45 minus.n30 minus.n29 27.752
R46 minus.n32 minus.n15 26.6728
R47 minus.n32 minus.n31 6.46073
R48 minus.n15 minus.n0 0.189894
R49 minus.n9 minus.n0 0.189894
R50 minus.n9 minus.n8 0.189894
R51 minus.n8 minus.n2 0.189894
R52 minus.n24 minus.n18 0.189894
R53 minus.n25 minus.n24 0.189894
R54 minus.n25 minus.n16 0.189894
R55 minus.n31 minus.n16 0.189894
R56 minus minus.n32 0.188
R57 source.n0 source.t10 243.255
R58 source.n7 source.t18 243.255
R59 source.n27 source.t13 243.254
R60 source.n20 source.t4 243.254
R61 source.n2 source.n1 223.454
R62 source.n4 source.n3 223.454
R63 source.n6 source.n5 223.454
R64 source.n9 source.n8 223.454
R65 source.n11 source.n10 223.454
R66 source.n13 source.n12 223.454
R67 source.n26 source.n25 223.453
R68 source.n24 source.n23 223.453
R69 source.n22 source.n21 223.453
R70 source.n19 source.n18 223.453
R71 source.n17 source.n16 223.453
R72 source.n15 source.n14 223.453
R73 source.n25 source.t23 19.8005
R74 source.n25 source.t12 19.8005
R75 source.n23 source.t22 19.8005
R76 source.n23 source.t14 19.8005
R77 source.n21 source.t20 19.8005
R78 source.n21 source.t16 19.8005
R79 source.n18 source.t8 19.8005
R80 source.n18 source.t5 19.8005
R81 source.n16 source.t0 19.8005
R82 source.n16 source.t6 19.8005
R83 source.n14 source.t3 19.8005
R84 source.n14 source.t25 19.8005
R85 source.n1 source.t9 19.8005
R86 source.n1 source.t26 19.8005
R87 source.n3 source.t2 19.8005
R88 source.n3 source.t1 19.8005
R89 source.n5 source.t27 19.8005
R90 source.n5 source.t7 19.8005
R91 source.n8 source.t21 19.8005
R92 source.n8 source.t11 19.8005
R93 source.n10 source.t17 19.8005
R94 source.n10 source.t19 19.8005
R95 source.n12 source.t24 19.8005
R96 source.n12 source.t15 19.8005
R97 source.n15 source.n13 13.8682
R98 source.n28 source.n0 7.91991
R99 source.n28 source.n27 5.49188
R100 source.n7 source.n6 0.698776
R101 source.n22 source.n20 0.698776
R102 source.n13 source.n11 0.457397
R103 source.n11 source.n9 0.457397
R104 source.n9 source.n7 0.457397
R105 source.n6 source.n4 0.457397
R106 source.n4 source.n2 0.457397
R107 source.n2 source.n0 0.457397
R108 source.n17 source.n15 0.457397
R109 source.n19 source.n17 0.457397
R110 source.n20 source.n19 0.457397
R111 source.n24 source.n22 0.457397
R112 source.n26 source.n24 0.457397
R113 source.n27 source.n26 0.457397
R114 source source.n28 0.188
R115 drain_right.n1 drain_right.t5 260.389
R116 drain_right.n11 drain_right.t12 259.933
R117 drain_right.n8 drain_right.n6 240.589
R118 drain_right.n4 drain_right.n2 240.589
R119 drain_right.n8 drain_right.n7 240.132
R120 drain_right.n10 drain_right.n9 240.132
R121 drain_right.n4 drain_right.n3 240.131
R122 drain_right.n1 drain_right.n0 240.131
R123 drain_right drain_right.n5 21.1077
R124 drain_right.n2 drain_right.t11 19.8005
R125 drain_right.n2 drain_right.t8 19.8005
R126 drain_right.n3 drain_right.t6 19.8005
R127 drain_right.n3 drain_right.t2 19.8005
R128 drain_right.n0 drain_right.t1 19.8005
R129 drain_right.n0 drain_right.t10 19.8005
R130 drain_right.n6 drain_right.t7 19.8005
R131 drain_right.n6 drain_right.t4 19.8005
R132 drain_right.n7 drain_right.t0 19.8005
R133 drain_right.n7 drain_right.t13 19.8005
R134 drain_right.n9 drain_right.t9 19.8005
R135 drain_right.n9 drain_right.t3 19.8005
R136 drain_right drain_right.n11 5.88166
R137 drain_right.n11 drain_right.n10 0.457397
R138 drain_right.n10 drain_right.n8 0.457397
R139 drain_right.n5 drain_right.n1 0.287826
R140 drain_right.n5 drain_right.n4 0.0593781
R141 plus.n3 plus.t5 326.812
R142 plus.n14 plus.t1 326.812
R143 plus.n19 plus.t6 326.812
R144 plus.n30 plus.t7 326.812
R145 plus.n4 plus.t2 277.151
R146 plus.n6 plus.t13 277.151
R147 plus.n1 plus.t10 277.151
R148 plus.n11 plus.t9 277.151
R149 plus.n13 plus.t4 277.151
R150 plus.n20 plus.t11 277.151
R151 plus.n22 plus.t0 277.151
R152 plus.n17 plus.t8 277.151
R153 plus.n27 plus.t12 277.151
R154 plus.n29 plus.t3 277.151
R155 plus.n3 plus.n2 161.489
R156 plus.n19 plus.n18 161.489
R157 plus.n5 plus.n2 161.3
R158 plus.n8 plus.n7 161.3
R159 plus.n10 plus.n9 161.3
R160 plus.n12 plus.n0 161.3
R161 plus.n15 plus.n14 161.3
R162 plus.n21 plus.n18 161.3
R163 plus.n24 plus.n23 161.3
R164 plus.n26 plus.n25 161.3
R165 plus.n28 plus.n16 161.3
R166 plus.n31 plus.n30 161.3
R167 plus.n5 plus.n4 45.2793
R168 plus.n13 plus.n12 45.2793
R169 plus.n29 plus.n28 45.2793
R170 plus.n21 plus.n20 45.2793
R171 plus.n7 plus.n6 40.8975
R172 plus.n11 plus.n10 40.8975
R173 plus.n27 plus.n26 40.8975
R174 plus.n23 plus.n22 40.8975
R175 plus.n7 plus.n1 36.5157
R176 plus.n10 plus.n1 36.5157
R177 plus.n26 plus.n17 36.5157
R178 plus.n23 plus.n17 36.5157
R179 plus.n6 plus.n5 32.1338
R180 plus.n12 plus.n11 32.1338
R181 plus.n28 plus.n27 32.1338
R182 plus.n22 plus.n21 32.1338
R183 plus.n4 plus.n3 27.752
R184 plus.n14 plus.n13 27.752
R185 plus.n30 plus.n29 27.752
R186 plus.n20 plus.n19 27.752
R187 plus plus.n31 24.7206
R188 plus plus.n15 7.938
R189 plus.n8 plus.n2 0.189894
R190 plus.n9 plus.n8 0.189894
R191 plus.n9 plus.n0 0.189894
R192 plus.n15 plus.n0 0.189894
R193 plus.n31 plus.n16 0.189894
R194 plus.n25 plus.n16 0.189894
R195 plus.n25 plus.n24 0.189894
R196 plus.n24 plus.n18 0.189894
R197 drain_left.n7 drain_left.t8 260.389
R198 drain_left.n1 drain_left.t6 260.389
R199 drain_left.n4 drain_left.n2 240.589
R200 drain_left.n11 drain_left.n10 240.132
R201 drain_left.n9 drain_left.n8 240.132
R202 drain_left.n7 drain_left.n6 240.132
R203 drain_left.n4 drain_left.n3 240.131
R204 drain_left.n1 drain_left.n0 240.131
R205 drain_left drain_left.n5 21.6609
R206 drain_left.n2 drain_left.t2 19.8005
R207 drain_left.n2 drain_left.t7 19.8005
R208 drain_left.n3 drain_left.t5 19.8005
R209 drain_left.n3 drain_left.t13 19.8005
R210 drain_left.n0 drain_left.t10 19.8005
R211 drain_left.n0 drain_left.t1 19.8005
R212 drain_left.n10 drain_left.t9 19.8005
R213 drain_left.n10 drain_left.t12 19.8005
R214 drain_left.n8 drain_left.t3 19.8005
R215 drain_left.n8 drain_left.t4 19.8005
R216 drain_left.n6 drain_left.t11 19.8005
R217 drain_left.n6 drain_left.t0 19.8005
R218 drain_left drain_left.n11 6.11011
R219 drain_left.n9 drain_left.n7 0.457397
R220 drain_left.n11 drain_left.n9 0.457397
R221 drain_left.n5 drain_left.n1 0.287826
R222 drain_left.n5 drain_left.n4 0.0593781
C0 drain_right drain_left 0.79079f
C1 drain_right minus 0.751013f
C2 drain_left minus 0.17873f
C3 drain_right source 5.119f
C4 drain_left source 5.12134f
C5 source minus 0.942045f
C6 drain_right plus 0.312711f
C7 drain_left plus 0.900745f
C8 plus minus 3.07747f
C9 plus source 0.955967f
C10 drain_right a_n1564_n1088# 3.52064f
C11 drain_left a_n1564_n1088# 3.74526f
C12 source a_n1564_n1088# 2.091053f
C13 minus a_n1564_n1088# 5.154123f
C14 plus a_n1564_n1088# 5.869838f
C15 drain_left.t6 a_n1564_n1088# 0.128553f
C16 drain_left.t10 a_n1564_n1088# 0.020715f
C17 drain_left.t1 a_n1564_n1088# 0.020715f
C18 drain_left.n0 a_n1564_n1088# 0.080491f
C19 drain_left.n1 a_n1564_n1088# 0.489188f
C20 drain_left.t2 a_n1564_n1088# 0.020715f
C21 drain_left.t7 a_n1564_n1088# 0.020715f
C22 drain_left.n2 a_n1564_n1088# 0.081006f
C23 drain_left.t5 a_n1564_n1088# 0.020715f
C24 drain_left.t13 a_n1564_n1088# 0.020715f
C25 drain_left.n3 a_n1564_n1088# 0.080491f
C26 drain_left.n4 a_n1564_n1088# 0.507742f
C27 drain_left.n5 a_n1564_n1088# 0.621295f
C28 drain_left.t8 a_n1564_n1088# 0.128553f
C29 drain_left.t11 a_n1564_n1088# 0.020715f
C30 drain_left.t0 a_n1564_n1088# 0.020715f
C31 drain_left.n6 a_n1564_n1088# 0.080491f
C32 drain_left.n7 a_n1564_n1088# 0.501395f
C33 drain_left.t3 a_n1564_n1088# 0.020715f
C34 drain_left.t4 a_n1564_n1088# 0.020715f
C35 drain_left.n8 a_n1564_n1088# 0.080491f
C36 drain_left.n9 a_n1564_n1088# 0.260498f
C37 drain_left.t9 a_n1564_n1088# 0.020715f
C38 drain_left.t12 a_n1564_n1088# 0.020715f
C39 drain_left.n10 a_n1564_n1088# 0.080491f
C40 drain_left.n11 a_n1564_n1088# 0.475031f
C41 plus.n0 a_n1564_n1088# 0.036024f
C42 plus.t4 a_n1564_n1088# 0.02221f
C43 plus.t9 a_n1564_n1088# 0.02221f
C44 plus.t10 a_n1564_n1088# 0.02221f
C45 plus.n1 a_n1564_n1088# 0.026585f
C46 plus.n2 a_n1564_n1088# 0.080435f
C47 plus.t13 a_n1564_n1088# 0.02221f
C48 plus.t2 a_n1564_n1088# 0.02221f
C49 plus.t5 a_n1564_n1088# 0.026385f
C50 plus.n3 a_n1564_n1088# 0.035967f
C51 plus.n4 a_n1564_n1088# 0.026585f
C52 plus.n5 a_n1564_n1088# 0.012617f
C53 plus.n6 a_n1564_n1088# 0.026585f
C54 plus.n7 a_n1564_n1088# 0.012617f
C55 plus.n8 a_n1564_n1088# 0.036024f
C56 plus.n9 a_n1564_n1088# 0.036024f
C57 plus.n10 a_n1564_n1088# 0.012617f
C58 plus.n11 a_n1564_n1088# 0.026585f
C59 plus.n12 a_n1564_n1088# 0.012617f
C60 plus.n13 a_n1564_n1088# 0.026585f
C61 plus.t1 a_n1564_n1088# 0.026385f
C62 plus.n14 a_n1564_n1088# 0.035915f
C63 plus.n15 a_n1564_n1088# 0.243461f
C64 plus.n16 a_n1564_n1088# 0.036024f
C65 plus.t7 a_n1564_n1088# 0.026385f
C66 plus.t3 a_n1564_n1088# 0.02221f
C67 plus.t12 a_n1564_n1088# 0.02221f
C68 plus.t8 a_n1564_n1088# 0.02221f
C69 plus.n17 a_n1564_n1088# 0.026585f
C70 plus.n18 a_n1564_n1088# 0.080435f
C71 plus.t0 a_n1564_n1088# 0.02221f
C72 plus.t11 a_n1564_n1088# 0.02221f
C73 plus.t6 a_n1564_n1088# 0.026385f
C74 plus.n19 a_n1564_n1088# 0.035967f
C75 plus.n20 a_n1564_n1088# 0.026585f
C76 plus.n21 a_n1564_n1088# 0.012617f
C77 plus.n22 a_n1564_n1088# 0.026585f
C78 plus.n23 a_n1564_n1088# 0.012617f
C79 plus.n24 a_n1564_n1088# 0.036024f
C80 plus.n25 a_n1564_n1088# 0.036024f
C81 plus.n26 a_n1564_n1088# 0.012617f
C82 plus.n27 a_n1564_n1088# 0.026585f
C83 plus.n28 a_n1564_n1088# 0.012617f
C84 plus.n29 a_n1564_n1088# 0.026585f
C85 plus.n30 a_n1564_n1088# 0.035915f
C86 plus.n31 a_n1564_n1088# 0.740096f
C87 drain_right.t5 a_n1564_n1088# 0.13119f
C88 drain_right.t1 a_n1564_n1088# 0.02114f
C89 drain_right.t10 a_n1564_n1088# 0.02114f
C90 drain_right.n0 a_n1564_n1088# 0.082143f
C91 drain_right.n1 a_n1564_n1088# 0.499226f
C92 drain_right.t11 a_n1564_n1088# 0.02114f
C93 drain_right.t8 a_n1564_n1088# 0.02114f
C94 drain_right.n2 a_n1564_n1088# 0.082668f
C95 drain_right.t6 a_n1564_n1088# 0.02114f
C96 drain_right.t2 a_n1564_n1088# 0.02114f
C97 drain_right.n3 a_n1564_n1088# 0.082143f
C98 drain_right.n4 a_n1564_n1088# 0.518161f
C99 drain_right.n5 a_n1564_n1088# 0.582244f
C100 drain_right.t7 a_n1564_n1088# 0.02114f
C101 drain_right.t4 a_n1564_n1088# 0.02114f
C102 drain_right.n6 a_n1564_n1088# 0.082668f
C103 drain_right.t0 a_n1564_n1088# 0.02114f
C104 drain_right.t13 a_n1564_n1088# 0.02114f
C105 drain_right.n7 a_n1564_n1088# 0.082143f
C106 drain_right.n8 a_n1564_n1088# 0.541936f
C107 drain_right.t9 a_n1564_n1088# 0.02114f
C108 drain_right.t3 a_n1564_n1088# 0.02114f
C109 drain_right.n9 a_n1564_n1088# 0.082143f
C110 drain_right.n10 a_n1564_n1088# 0.265843f
C111 drain_right.t12 a_n1564_n1088# 0.130758f
C112 drain_right.n11 a_n1564_n1088# 0.463702f
C113 source.t10 a_n1564_n1088# 0.154609f
C114 source.n0 a_n1564_n1088# 0.646354f
C115 source.t9 a_n1564_n1088# 0.027778f
C116 source.t26 a_n1564_n1088# 0.027778f
C117 source.n1 a_n1564_n1088# 0.090089f
C118 source.n2 a_n1564_n1088# 0.319395f
C119 source.t2 a_n1564_n1088# 0.027778f
C120 source.t1 a_n1564_n1088# 0.027778f
C121 source.n3 a_n1564_n1088# 0.090089f
C122 source.n4 a_n1564_n1088# 0.319395f
C123 source.t27 a_n1564_n1088# 0.027778f
C124 source.t7 a_n1564_n1088# 0.027778f
C125 source.n5 a_n1564_n1088# 0.090089f
C126 source.n6 a_n1564_n1088# 0.346735f
C127 source.t18 a_n1564_n1088# 0.154609f
C128 source.n7 a_n1564_n1088# 0.357973f
C129 source.t21 a_n1564_n1088# 0.027778f
C130 source.t11 a_n1564_n1088# 0.027778f
C131 source.n8 a_n1564_n1088# 0.090089f
C132 source.n9 a_n1564_n1088# 0.319395f
C133 source.t17 a_n1564_n1088# 0.027778f
C134 source.t19 a_n1564_n1088# 0.027778f
C135 source.n10 a_n1564_n1088# 0.090089f
C136 source.n11 a_n1564_n1088# 0.319395f
C137 source.t24 a_n1564_n1088# 0.027778f
C138 source.t15 a_n1564_n1088# 0.027778f
C139 source.n12 a_n1564_n1088# 0.090089f
C140 source.n13 a_n1564_n1088# 0.966524f
C141 source.t3 a_n1564_n1088# 0.027778f
C142 source.t25 a_n1564_n1088# 0.027778f
C143 source.n14 a_n1564_n1088# 0.090089f
C144 source.n15 a_n1564_n1088# 0.966524f
C145 source.t0 a_n1564_n1088# 0.027778f
C146 source.t6 a_n1564_n1088# 0.027778f
C147 source.n16 a_n1564_n1088# 0.090089f
C148 source.n17 a_n1564_n1088# 0.319395f
C149 source.t8 a_n1564_n1088# 0.027778f
C150 source.t5 a_n1564_n1088# 0.027778f
C151 source.n18 a_n1564_n1088# 0.090089f
C152 source.n19 a_n1564_n1088# 0.319395f
C153 source.t4 a_n1564_n1088# 0.154609f
C154 source.n20 a_n1564_n1088# 0.357974f
C155 source.t20 a_n1564_n1088# 0.027778f
C156 source.t16 a_n1564_n1088# 0.027778f
C157 source.n21 a_n1564_n1088# 0.090089f
C158 source.n22 a_n1564_n1088# 0.346735f
C159 source.t22 a_n1564_n1088# 0.027778f
C160 source.t14 a_n1564_n1088# 0.027778f
C161 source.n23 a_n1564_n1088# 0.090089f
C162 source.n24 a_n1564_n1088# 0.319395f
C163 source.t23 a_n1564_n1088# 0.027778f
C164 source.t12 a_n1564_n1088# 0.027778f
C165 source.n25 a_n1564_n1088# 0.090089f
C166 source.n26 a_n1564_n1088# 0.319395f
C167 source.t13 a_n1564_n1088# 0.154609f
C168 source.n27 a_n1564_n1088# 0.522703f
C169 source.n28 a_n1564_n1088# 0.707969f
C170 minus.n0 a_n1564_n1088# 0.035197f
C171 minus.t1 a_n1564_n1088# 0.025779f
C172 minus.t4 a_n1564_n1088# 0.0217f
C173 minus.t10 a_n1564_n1088# 0.0217f
C174 minus.t13 a_n1564_n1088# 0.0217f
C175 minus.n1 a_n1564_n1088# 0.025975f
C176 minus.n2 a_n1564_n1088# 0.078589f
C177 minus.t0 a_n1564_n1088# 0.0217f
C178 minus.t6 a_n1564_n1088# 0.0217f
C179 minus.t9 a_n1564_n1088# 0.025779f
C180 minus.n3 a_n1564_n1088# 0.035142f
C181 minus.n4 a_n1564_n1088# 0.025975f
C182 minus.n5 a_n1564_n1088# 0.012327f
C183 minus.n6 a_n1564_n1088# 0.025975f
C184 minus.n7 a_n1564_n1088# 0.012327f
C185 minus.n8 a_n1564_n1088# 0.035197f
C186 minus.n9 a_n1564_n1088# 0.035197f
C187 minus.n10 a_n1564_n1088# 0.012327f
C188 minus.n11 a_n1564_n1088# 0.025975f
C189 minus.n12 a_n1564_n1088# 0.012327f
C190 minus.n13 a_n1564_n1088# 0.025975f
C191 minus.n14 a_n1564_n1088# 0.035091f
C192 minus.n15 a_n1564_n1088# 0.74292f
C193 minus.n16 a_n1564_n1088# 0.035197f
C194 minus.t2 a_n1564_n1088# 0.0217f
C195 minus.t11 a_n1564_n1088# 0.0217f
C196 minus.t7 a_n1564_n1088# 0.0217f
C197 minus.n17 a_n1564_n1088# 0.025975f
C198 minus.n18 a_n1564_n1088# 0.078589f
C199 minus.t3 a_n1564_n1088# 0.0217f
C200 minus.t12 a_n1564_n1088# 0.0217f
C201 minus.t8 a_n1564_n1088# 0.025779f
C202 minus.n19 a_n1564_n1088# 0.035142f
C203 minus.n20 a_n1564_n1088# 0.025975f
C204 minus.n21 a_n1564_n1088# 0.012327f
C205 minus.n22 a_n1564_n1088# 0.025975f
C206 minus.n23 a_n1564_n1088# 0.012327f
C207 minus.n24 a_n1564_n1088# 0.035197f
C208 minus.n25 a_n1564_n1088# 0.035197f
C209 minus.n26 a_n1564_n1088# 0.012327f
C210 minus.n27 a_n1564_n1088# 0.025975f
C211 minus.n28 a_n1564_n1088# 0.012327f
C212 minus.n29 a_n1564_n1088# 0.025975f
C213 minus.t5 a_n1564_n1088# 0.025779f
C214 minus.n30 a_n1564_n1088# 0.035091f
C215 minus.n31 a_n1564_n1088# 0.226845f
C216 minus.n32 a_n1564_n1088# 0.919819f
.ends

