* NGSPICE file created from diffpair69.ext - technology: sky130A

.subckt diffpair69 minus drain_right drain_left source plus
X0 a_n3394_n1088# a_n3394_n1088# a_n3394_n1088# a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.7
X1 drain_left.t23 plus.t0 source.t30 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X2 source.t26 plus.t1 drain_left.t22 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X3 source.t21 plus.t2 drain_left.t21 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X4 source.t2 minus.t0 drain_right.t23 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X5 drain_left.t20 plus.t3 source.t14 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X6 source.t10 plus.t4 drain_left.t19 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X7 drain_left.t18 plus.t5 source.t24 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X8 source.t19 plus.t6 drain_left.t17 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X9 source.t31 plus.t7 drain_left.t16 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X10 drain_right.t22 minus.t1 source.t7 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X11 drain_right.t21 minus.t2 source.t37 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X12 source.t42 minus.t3 drain_right.t20 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X13 drain_right.t19 minus.t4 source.t0 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X14 a_n3394_n1088# a_n3394_n1088# a_n3394_n1088# a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X15 source.t27 plus.t8 drain_left.t15 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X16 drain_right.t18 minus.t5 source.t46 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X17 drain_right.t17 minus.t6 source.t1 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X18 drain_right.t16 minus.t7 source.t36 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X19 source.t41 minus.t8 drain_right.t15 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X20 drain_left.t14 plus.t9 source.t28 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X21 drain_right.t14 minus.t9 source.t9 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X22 source.t35 minus.t10 drain_right.t13 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X23 source.t23 plus.t10 drain_left.t13 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X24 drain_right.t12 minus.t11 source.t40 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X25 drain_left.t12 plus.t11 source.t29 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X26 drain_left.t11 plus.t12 source.t25 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X27 a_n3394_n1088# a_n3394_n1088# a_n3394_n1088# a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X28 source.t22 plus.t13 drain_left.t10 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X29 drain_left.t9 plus.t14 source.t12 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X30 source.t18 plus.t15 drain_left.t8 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X31 drain_right.t11 minus.t12 source.t8 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X32 a_n3394_n1088# a_n3394_n1088# a_n3394_n1088# a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X33 drain_left.t7 plus.t16 source.t20 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X34 drain_left.t6 plus.t17 source.t32 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X35 source.t47 minus.t13 drain_right.t10 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X36 source.t43 minus.t14 drain_right.t9 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X37 drain_right.t8 minus.t15 source.t6 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X38 drain_right.t7 minus.t16 source.t39 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X39 source.t45 minus.t17 drain_right.t6 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X40 source.t4 minus.t18 drain_right.t5 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X41 drain_left.t5 plus.t18 source.t13 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X42 source.t44 minus.t19 drain_right.t4 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X43 source.t5 minus.t20 drain_right.t3 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X44 source.t15 plus.t19 drain_left.t4 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X45 source.t34 minus.t21 drain_right.t2 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X46 source.t38 minus.t22 drain_right.t1 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X47 drain_right.t0 minus.t23 source.t3 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X48 drain_left.t3 plus.t20 source.t11 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X49 source.t17 plus.t21 drain_left.t2 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X50 source.t33 plus.t22 drain_left.t1 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X51 drain_left.t0 plus.t23 source.t16 a_n3394_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
R0 plus.n13 plus.n12 161.3
R1 plus.n14 plus.n9 161.3
R2 plus.n16 plus.n15 161.3
R3 plus.n17 plus.n8 161.3
R4 plus.n19 plus.n18 161.3
R5 plus.n20 plus.n7 161.3
R6 plus.n22 plus.n21 161.3
R7 plus.n23 plus.n6 161.3
R8 plus.n25 plus.n24 161.3
R9 plus.n26 plus.n5 161.3
R10 plus.n28 plus.n27 161.3
R11 plus.n29 plus.n4 161.3
R12 plus.n31 plus.n30 161.3
R13 plus.n32 plus.n3 161.3
R14 plus.n34 plus.n33 161.3
R15 plus.n35 plus.n2 161.3
R16 plus.n37 plus.n36 161.3
R17 plus.n38 plus.n1 161.3
R18 plus.n39 plus.n0 161.3
R19 plus.n41 plus.n40 161.3
R20 plus.n55 plus.n54 161.3
R21 plus.n56 plus.n51 161.3
R22 plus.n58 plus.n57 161.3
R23 plus.n59 plus.n50 161.3
R24 plus.n61 plus.n60 161.3
R25 plus.n62 plus.n49 161.3
R26 plus.n64 plus.n63 161.3
R27 plus.n65 plus.n48 161.3
R28 plus.n67 plus.n66 161.3
R29 plus.n68 plus.n47 161.3
R30 plus.n70 plus.n69 161.3
R31 plus.n71 plus.n46 161.3
R32 plus.n73 plus.n72 161.3
R33 plus.n74 plus.n45 161.3
R34 plus.n76 plus.n75 161.3
R35 plus.n77 plus.n44 161.3
R36 plus.n79 plus.n78 161.3
R37 plus.n80 plus.n43 161.3
R38 plus.n81 plus.n42 161.3
R39 plus.n83 plus.n82 161.3
R40 plus.n11 plus.t7 116.906
R41 plus.n53 plus.t11 116.906
R42 plus.n40 plus.t0 90.5476
R43 plus.n38 plus.t13 90.5476
R44 plus.n2 plus.t3 90.5476
R45 plus.n32 plus.t21 90.5476
R46 plus.n4 plus.t9 90.5476
R47 plus.n26 plus.t1 90.5476
R48 plus.n6 plus.t14 90.5476
R49 plus.n20 plus.t6 90.5476
R50 plus.n8 plus.t12 90.5476
R51 plus.n14 plus.t2 90.5476
R52 plus.n10 plus.t17 90.5476
R53 plus.n82 plus.t19 90.5476
R54 plus.n80 plus.t20 90.5476
R55 plus.n44 plus.t15 90.5476
R56 plus.n74 plus.t16 90.5476
R57 plus.n46 plus.t8 90.5476
R58 plus.n68 plus.t5 90.5476
R59 plus.n48 plus.t4 90.5476
R60 plus.n62 plus.t23 90.5476
R61 plus.n50 plus.t22 90.5476
R62 plus.n56 plus.t18 90.5476
R63 plus.n52 plus.t10 90.5476
R64 plus.n40 plus.n39 46.0096
R65 plus.n82 plus.n81 46.0096
R66 plus.n12 plus.n11 45.0871
R67 plus.n54 plus.n53 45.0871
R68 plus.n38 plus.n37 41.6278
R69 plus.n13 plus.n10 41.6278
R70 plus.n80 plus.n79 41.6278
R71 plus.n55 plus.n52 41.6278
R72 plus.n33 plus.n2 37.246
R73 plus.n15 plus.n14 37.246
R74 plus.n75 plus.n44 37.246
R75 plus.n57 plus.n56 37.246
R76 plus.n32 plus.n31 32.8641
R77 plus.n19 plus.n8 32.8641
R78 plus.n74 plus.n73 32.8641
R79 plus.n61 plus.n50 32.8641
R80 plus plus.n83 31.8702
R81 plus.n27 plus.n4 28.4823
R82 plus.n21 plus.n20 28.4823
R83 plus.n69 plus.n46 28.4823
R84 plus.n63 plus.n62 28.4823
R85 plus.n25 plus.n6 24.1005
R86 plus.n26 plus.n25 24.1005
R87 plus.n68 plus.n67 24.1005
R88 plus.n67 plus.n48 24.1005
R89 plus.n27 plus.n26 19.7187
R90 plus.n21 plus.n6 19.7187
R91 plus.n69 plus.n68 19.7187
R92 plus.n63 plus.n48 19.7187
R93 plus.n31 plus.n4 15.3369
R94 plus.n20 plus.n19 15.3369
R95 plus.n73 plus.n46 15.3369
R96 plus.n62 plus.n61 15.3369
R97 plus.n11 plus.n10 14.1472
R98 plus.n53 plus.n52 14.1472
R99 plus.n33 plus.n32 10.955
R100 plus.n15 plus.n8 10.955
R101 plus.n75 plus.n74 10.955
R102 plus.n57 plus.n50 10.955
R103 plus plus.n41 8.1558
R104 plus.n37 plus.n2 6.57323
R105 plus.n14 plus.n13 6.57323
R106 plus.n79 plus.n44 6.57323
R107 plus.n56 plus.n55 6.57323
R108 plus.n39 plus.n38 2.19141
R109 plus.n81 plus.n80 2.19141
R110 plus.n12 plus.n9 0.189894
R111 plus.n16 plus.n9 0.189894
R112 plus.n17 plus.n16 0.189894
R113 plus.n18 plus.n17 0.189894
R114 plus.n18 plus.n7 0.189894
R115 plus.n22 plus.n7 0.189894
R116 plus.n23 plus.n22 0.189894
R117 plus.n24 plus.n23 0.189894
R118 plus.n24 plus.n5 0.189894
R119 plus.n28 plus.n5 0.189894
R120 plus.n29 plus.n28 0.189894
R121 plus.n30 plus.n29 0.189894
R122 plus.n30 plus.n3 0.189894
R123 plus.n34 plus.n3 0.189894
R124 plus.n35 plus.n34 0.189894
R125 plus.n36 plus.n35 0.189894
R126 plus.n36 plus.n1 0.189894
R127 plus.n1 plus.n0 0.189894
R128 plus.n41 plus.n0 0.189894
R129 plus.n83 plus.n42 0.189894
R130 plus.n43 plus.n42 0.189894
R131 plus.n78 plus.n43 0.189894
R132 plus.n78 plus.n77 0.189894
R133 plus.n77 plus.n76 0.189894
R134 plus.n76 plus.n45 0.189894
R135 plus.n72 plus.n45 0.189894
R136 plus.n72 plus.n71 0.189894
R137 plus.n71 plus.n70 0.189894
R138 plus.n70 plus.n47 0.189894
R139 plus.n66 plus.n47 0.189894
R140 plus.n66 plus.n65 0.189894
R141 plus.n65 plus.n64 0.189894
R142 plus.n64 plus.n49 0.189894
R143 plus.n60 plus.n49 0.189894
R144 plus.n60 plus.n59 0.189894
R145 plus.n59 plus.n58 0.189894
R146 plus.n58 plus.n51 0.189894
R147 plus.n54 plus.n51 0.189894
R148 source.n0 source.t30 243.255
R149 source.n11 source.t31 243.255
R150 source.n12 source.t8 243.255
R151 source.n23 source.t47 243.255
R152 source.n47 source.t6 243.254
R153 source.n36 source.t42 243.254
R154 source.n35 source.t29 243.254
R155 source.n24 source.t15 243.254
R156 source.n2 source.n1 223.454
R157 source.n4 source.n3 223.454
R158 source.n6 source.n5 223.454
R159 source.n8 source.n7 223.454
R160 source.n10 source.n9 223.454
R161 source.n14 source.n13 223.454
R162 source.n16 source.n15 223.454
R163 source.n18 source.n17 223.454
R164 source.n20 source.n19 223.454
R165 source.n22 source.n21 223.454
R166 source.n46 source.n45 223.453
R167 source.n44 source.n43 223.453
R168 source.n42 source.n41 223.453
R169 source.n40 source.n39 223.453
R170 source.n38 source.n37 223.453
R171 source.n34 source.n33 223.453
R172 source.n32 source.n31 223.453
R173 source.n30 source.n29 223.453
R174 source.n28 source.n27 223.453
R175 source.n26 source.n25 223.453
R176 source.n45 source.t9 19.8005
R177 source.n45 source.t4 19.8005
R178 source.n43 source.t3 19.8005
R179 source.n43 source.t5 19.8005
R180 source.n41 source.t39 19.8005
R181 source.n41 source.t43 19.8005
R182 source.n39 source.t36 19.8005
R183 source.n39 source.t35 19.8005
R184 source.n37 source.t37 19.8005
R185 source.n37 source.t41 19.8005
R186 source.n33 source.t13 19.8005
R187 source.n33 source.t23 19.8005
R188 source.n31 source.t16 19.8005
R189 source.n31 source.t33 19.8005
R190 source.n29 source.t24 19.8005
R191 source.n29 source.t10 19.8005
R192 source.n27 source.t20 19.8005
R193 source.n27 source.t27 19.8005
R194 source.n25 source.t11 19.8005
R195 source.n25 source.t18 19.8005
R196 source.n1 source.t14 19.8005
R197 source.n1 source.t22 19.8005
R198 source.n3 source.t28 19.8005
R199 source.n3 source.t17 19.8005
R200 source.n5 source.t12 19.8005
R201 source.n5 source.t26 19.8005
R202 source.n7 source.t25 19.8005
R203 source.n7 source.t19 19.8005
R204 source.n9 source.t32 19.8005
R205 source.n9 source.t21 19.8005
R206 source.n13 source.t40 19.8005
R207 source.n13 source.t2 19.8005
R208 source.n15 source.t1 19.8005
R209 source.n15 source.t34 19.8005
R210 source.n17 source.t46 19.8005
R211 source.n17 source.t38 19.8005
R212 source.n19 source.t0 19.8005
R213 source.n19 source.t44 19.8005
R214 source.n21 source.t7 19.8005
R215 source.n21 source.t45 19.8005
R216 source.n24 source.n23 13.8423
R217 source.n48 source.n0 8.13543
R218 source.n48 source.n47 5.7074
R219 source.n23 source.n22 0.888431
R220 source.n22 source.n20 0.888431
R221 source.n20 source.n18 0.888431
R222 source.n18 source.n16 0.888431
R223 source.n16 source.n14 0.888431
R224 source.n14 source.n12 0.888431
R225 source.n11 source.n10 0.888431
R226 source.n10 source.n8 0.888431
R227 source.n8 source.n6 0.888431
R228 source.n6 source.n4 0.888431
R229 source.n4 source.n2 0.888431
R230 source.n2 source.n0 0.888431
R231 source.n26 source.n24 0.888431
R232 source.n28 source.n26 0.888431
R233 source.n30 source.n28 0.888431
R234 source.n32 source.n30 0.888431
R235 source.n34 source.n32 0.888431
R236 source.n35 source.n34 0.888431
R237 source.n38 source.n36 0.888431
R238 source.n40 source.n38 0.888431
R239 source.n42 source.n40 0.888431
R240 source.n44 source.n42 0.888431
R241 source.n46 source.n44 0.888431
R242 source.n47 source.n46 0.888431
R243 source.n12 source.n11 0.470328
R244 source.n36 source.n35 0.470328
R245 source source.n48 0.188
R246 drain_left.n13 drain_left.n11 241.02
R247 drain_left.n7 drain_left.n5 241.019
R248 drain_left.n2 drain_left.n0 241.019
R249 drain_left.n21 drain_left.n20 240.132
R250 drain_left.n19 drain_left.n18 240.132
R251 drain_left.n17 drain_left.n16 240.132
R252 drain_left.n15 drain_left.n14 240.132
R253 drain_left.n13 drain_left.n12 240.132
R254 drain_left.n7 drain_left.n6 240.131
R255 drain_left.n9 drain_left.n8 240.131
R256 drain_left.n4 drain_left.n3 240.131
R257 drain_left.n2 drain_left.n1 240.131
R258 drain_left drain_left.n10 27.4691
R259 drain_left.n5 drain_left.t13 19.8005
R260 drain_left.n5 drain_left.t12 19.8005
R261 drain_left.n6 drain_left.t1 19.8005
R262 drain_left.n6 drain_left.t5 19.8005
R263 drain_left.n8 drain_left.t19 19.8005
R264 drain_left.n8 drain_left.t0 19.8005
R265 drain_left.n3 drain_left.t15 19.8005
R266 drain_left.n3 drain_left.t18 19.8005
R267 drain_left.n1 drain_left.t8 19.8005
R268 drain_left.n1 drain_left.t7 19.8005
R269 drain_left.n0 drain_left.t4 19.8005
R270 drain_left.n0 drain_left.t3 19.8005
R271 drain_left.n20 drain_left.t10 19.8005
R272 drain_left.n20 drain_left.t23 19.8005
R273 drain_left.n18 drain_left.t2 19.8005
R274 drain_left.n18 drain_left.t20 19.8005
R275 drain_left.n16 drain_left.t22 19.8005
R276 drain_left.n16 drain_left.t14 19.8005
R277 drain_left.n14 drain_left.t17 19.8005
R278 drain_left.n14 drain_left.t9 19.8005
R279 drain_left.n12 drain_left.t21 19.8005
R280 drain_left.n12 drain_left.t11 19.8005
R281 drain_left.n11 drain_left.t16 19.8005
R282 drain_left.n11 drain_left.t6 19.8005
R283 drain_left drain_left.n21 6.54115
R284 drain_left.n9 drain_left.n7 0.888431
R285 drain_left.n4 drain_left.n2 0.888431
R286 drain_left.n15 drain_left.n13 0.888431
R287 drain_left.n17 drain_left.n15 0.888431
R288 drain_left.n19 drain_left.n17 0.888431
R289 drain_left.n21 drain_left.n19 0.888431
R290 drain_left.n10 drain_left.n9 0.389119
R291 drain_left.n10 drain_left.n4 0.389119
R292 minus.n41 minus.n40 161.3
R293 minus.n39 minus.n0 161.3
R294 minus.n38 minus.n37 161.3
R295 minus.n36 minus.n1 161.3
R296 minus.n35 minus.n34 161.3
R297 minus.n33 minus.n2 161.3
R298 minus.n32 minus.n31 161.3
R299 minus.n30 minus.n3 161.3
R300 minus.n29 minus.n28 161.3
R301 minus.n27 minus.n4 161.3
R302 minus.n26 minus.n25 161.3
R303 minus.n24 minus.n5 161.3
R304 minus.n23 minus.n22 161.3
R305 minus.n21 minus.n6 161.3
R306 minus.n20 minus.n19 161.3
R307 minus.n18 minus.n7 161.3
R308 minus.n17 minus.n16 161.3
R309 minus.n15 minus.n8 161.3
R310 minus.n14 minus.n13 161.3
R311 minus.n12 minus.n9 161.3
R312 minus.n83 minus.n82 161.3
R313 minus.n81 minus.n42 161.3
R314 minus.n80 minus.n79 161.3
R315 minus.n78 minus.n43 161.3
R316 minus.n77 minus.n76 161.3
R317 minus.n75 minus.n44 161.3
R318 minus.n74 minus.n73 161.3
R319 minus.n72 minus.n45 161.3
R320 minus.n71 minus.n70 161.3
R321 minus.n69 minus.n46 161.3
R322 minus.n68 minus.n67 161.3
R323 minus.n66 minus.n47 161.3
R324 minus.n65 minus.n64 161.3
R325 minus.n63 minus.n48 161.3
R326 minus.n62 minus.n61 161.3
R327 minus.n60 minus.n49 161.3
R328 minus.n59 minus.n58 161.3
R329 minus.n57 minus.n50 161.3
R330 minus.n56 minus.n55 161.3
R331 minus.n54 minus.n51 161.3
R332 minus.n11 minus.t12 116.906
R333 minus.n53 minus.t3 116.906
R334 minus.n10 minus.t0 90.5476
R335 minus.n14 minus.t11 90.5476
R336 minus.n16 minus.t21 90.5476
R337 minus.n20 minus.t6 90.5476
R338 minus.n22 minus.t22 90.5476
R339 minus.n26 minus.t5 90.5476
R340 minus.n28 minus.t19 90.5476
R341 minus.n32 minus.t4 90.5476
R342 minus.n34 minus.t17 90.5476
R343 minus.n38 minus.t1 90.5476
R344 minus.n40 minus.t13 90.5476
R345 minus.n52 minus.t2 90.5476
R346 minus.n56 minus.t8 90.5476
R347 minus.n58 minus.t7 90.5476
R348 minus.n62 minus.t10 90.5476
R349 minus.n64 minus.t16 90.5476
R350 minus.n68 minus.t14 90.5476
R351 minus.n70 minus.t23 90.5476
R352 minus.n74 minus.t20 90.5476
R353 minus.n76 minus.t9 90.5476
R354 minus.n80 minus.t18 90.5476
R355 minus.n82 minus.t15 90.5476
R356 minus.n40 minus.n39 46.0096
R357 minus.n82 minus.n81 46.0096
R358 minus.n12 minus.n11 45.0871
R359 minus.n54 minus.n53 45.0871
R360 minus.n10 minus.n9 41.6278
R361 minus.n38 minus.n1 41.6278
R362 minus.n52 minus.n51 41.6278
R363 minus.n80 minus.n43 41.6278
R364 minus.n15 minus.n14 37.246
R365 minus.n34 minus.n33 37.246
R366 minus.n57 minus.n56 37.246
R367 minus.n76 minus.n75 37.246
R368 minus.n84 minus.n41 33.8225
R369 minus.n16 minus.n7 32.8641
R370 minus.n32 minus.n3 32.8641
R371 minus.n58 minus.n49 32.8641
R372 minus.n74 minus.n45 32.8641
R373 minus.n21 minus.n20 28.4823
R374 minus.n28 minus.n27 28.4823
R375 minus.n63 minus.n62 28.4823
R376 minus.n70 minus.n69 28.4823
R377 minus.n26 minus.n5 24.1005
R378 minus.n22 minus.n5 24.1005
R379 minus.n64 minus.n47 24.1005
R380 minus.n68 minus.n47 24.1005
R381 minus.n22 minus.n21 19.7187
R382 minus.n27 minus.n26 19.7187
R383 minus.n64 minus.n63 19.7187
R384 minus.n69 minus.n68 19.7187
R385 minus.n20 minus.n7 15.3369
R386 minus.n28 minus.n3 15.3369
R387 minus.n62 minus.n49 15.3369
R388 minus.n70 minus.n45 15.3369
R389 minus.n11 minus.n10 14.1472
R390 minus.n53 minus.n52 14.1472
R391 minus.n16 minus.n15 10.955
R392 minus.n33 minus.n32 10.955
R393 minus.n58 minus.n57 10.955
R394 minus.n75 minus.n74 10.955
R395 minus.n84 minus.n83 6.67853
R396 minus.n14 minus.n9 6.57323
R397 minus.n34 minus.n1 6.57323
R398 minus.n56 minus.n51 6.57323
R399 minus.n76 minus.n43 6.57323
R400 minus.n39 minus.n38 2.19141
R401 minus.n81 minus.n80 2.19141
R402 minus.n41 minus.n0 0.189894
R403 minus.n37 minus.n0 0.189894
R404 minus.n37 minus.n36 0.189894
R405 minus.n36 minus.n35 0.189894
R406 minus.n35 minus.n2 0.189894
R407 minus.n31 minus.n2 0.189894
R408 minus.n31 minus.n30 0.189894
R409 minus.n30 minus.n29 0.189894
R410 minus.n29 minus.n4 0.189894
R411 minus.n25 minus.n4 0.189894
R412 minus.n25 minus.n24 0.189894
R413 minus.n24 minus.n23 0.189894
R414 minus.n23 minus.n6 0.189894
R415 minus.n19 minus.n6 0.189894
R416 minus.n19 minus.n18 0.189894
R417 minus.n18 minus.n17 0.189894
R418 minus.n17 minus.n8 0.189894
R419 minus.n13 minus.n8 0.189894
R420 minus.n13 minus.n12 0.189894
R421 minus.n55 minus.n54 0.189894
R422 minus.n55 minus.n50 0.189894
R423 minus.n59 minus.n50 0.189894
R424 minus.n60 minus.n59 0.189894
R425 minus.n61 minus.n60 0.189894
R426 minus.n61 minus.n48 0.189894
R427 minus.n65 minus.n48 0.189894
R428 minus.n66 minus.n65 0.189894
R429 minus.n67 minus.n66 0.189894
R430 minus.n67 minus.n46 0.189894
R431 minus.n71 minus.n46 0.189894
R432 minus.n72 minus.n71 0.189894
R433 minus.n73 minus.n72 0.189894
R434 minus.n73 minus.n44 0.189894
R435 minus.n77 minus.n44 0.189894
R436 minus.n78 minus.n77 0.189894
R437 minus.n79 minus.n78 0.189894
R438 minus.n79 minus.n42 0.189894
R439 minus.n83 minus.n42 0.189894
R440 minus minus.n84 0.188
R441 drain_right.n13 drain_right.n11 241.02
R442 drain_right.n7 drain_right.n5 241.019
R443 drain_right.n2 drain_right.n0 241.019
R444 drain_right.n13 drain_right.n12 240.132
R445 drain_right.n15 drain_right.n14 240.132
R446 drain_right.n17 drain_right.n16 240.132
R447 drain_right.n19 drain_right.n18 240.132
R448 drain_right.n21 drain_right.n20 240.132
R449 drain_right.n7 drain_right.n6 240.131
R450 drain_right.n9 drain_right.n8 240.131
R451 drain_right.n4 drain_right.n3 240.131
R452 drain_right.n2 drain_right.n1 240.131
R453 drain_right drain_right.n10 26.9159
R454 drain_right.n5 drain_right.t5 19.8005
R455 drain_right.n5 drain_right.t8 19.8005
R456 drain_right.n6 drain_right.t3 19.8005
R457 drain_right.n6 drain_right.t14 19.8005
R458 drain_right.n8 drain_right.t9 19.8005
R459 drain_right.n8 drain_right.t0 19.8005
R460 drain_right.n3 drain_right.t13 19.8005
R461 drain_right.n3 drain_right.t7 19.8005
R462 drain_right.n1 drain_right.t15 19.8005
R463 drain_right.n1 drain_right.t16 19.8005
R464 drain_right.n0 drain_right.t20 19.8005
R465 drain_right.n0 drain_right.t21 19.8005
R466 drain_right.n11 drain_right.t23 19.8005
R467 drain_right.n11 drain_right.t11 19.8005
R468 drain_right.n12 drain_right.t2 19.8005
R469 drain_right.n12 drain_right.t12 19.8005
R470 drain_right.n14 drain_right.t1 19.8005
R471 drain_right.n14 drain_right.t17 19.8005
R472 drain_right.n16 drain_right.t4 19.8005
R473 drain_right.n16 drain_right.t18 19.8005
R474 drain_right.n18 drain_right.t6 19.8005
R475 drain_right.n18 drain_right.t19 19.8005
R476 drain_right.n20 drain_right.t10 19.8005
R477 drain_right.n20 drain_right.t22 19.8005
R478 drain_right drain_right.n21 6.54115
R479 drain_right.n9 drain_right.n7 0.888431
R480 drain_right.n4 drain_right.n2 0.888431
R481 drain_right.n21 drain_right.n19 0.888431
R482 drain_right.n19 drain_right.n17 0.888431
R483 drain_right.n17 drain_right.n15 0.888431
R484 drain_right.n15 drain_right.n13 0.888431
R485 drain_right.n10 drain_right.n9 0.389119
R486 drain_right.n10 drain_right.n4 0.389119
C0 drain_left plus 2.31018f
C1 source minus 2.9706f
C2 drain_right plus 0.507807f
C3 drain_left minus 0.181981f
C4 drain_right minus 1.97005f
C5 drain_left source 6.71879f
C6 drain_right source 6.72135f
C7 minus plus 5.35389f
C8 drain_right drain_left 1.87049f
C9 source plus 2.98446f
C10 drain_right a_n3394_n1088# 5.35695f
C11 drain_left a_n3394_n1088# 6.26671f
C12 source a_n3394_n1088# 3.060339f
C13 minus a_n3394_n1088# 12.80733f
C14 plus a_n3394_n1088# 14.275311f
C15 drain_right.t20 a_n3394_n1088# 0.016395f
C16 drain_right.t21 a_n3394_n1088# 0.016395f
C17 drain_right.n0 a_n3394_n1088# 0.064707f
C18 drain_right.t15 a_n3394_n1088# 0.016395f
C19 drain_right.t16 a_n3394_n1088# 0.016395f
C20 drain_right.n1 a_n3394_n1088# 0.063704f
C21 drain_right.n2 a_n3394_n1088# 0.53495f
C22 drain_right.t13 a_n3394_n1088# 0.016395f
C23 drain_right.t7 a_n3394_n1088# 0.016395f
C24 drain_right.n3 a_n3394_n1088# 0.063704f
C25 drain_right.n4 a_n3394_n1088# 0.231657f
C26 drain_right.t5 a_n3394_n1088# 0.016395f
C27 drain_right.t8 a_n3394_n1088# 0.016395f
C28 drain_right.n5 a_n3394_n1088# 0.064707f
C29 drain_right.t3 a_n3394_n1088# 0.016395f
C30 drain_right.t14 a_n3394_n1088# 0.016395f
C31 drain_right.n6 a_n3394_n1088# 0.063704f
C32 drain_right.n7 a_n3394_n1088# 0.53495f
C33 drain_right.t9 a_n3394_n1088# 0.016395f
C34 drain_right.t0 a_n3394_n1088# 0.016395f
C35 drain_right.n8 a_n3394_n1088# 0.063704f
C36 drain_right.n9 a_n3394_n1088# 0.231657f
C37 drain_right.n10 a_n3394_n1088# 0.853489f
C38 drain_right.t23 a_n3394_n1088# 0.016395f
C39 drain_right.t11 a_n3394_n1088# 0.016395f
C40 drain_right.n11 a_n3394_n1088# 0.064707f
C41 drain_right.t2 a_n3394_n1088# 0.016395f
C42 drain_right.t12 a_n3394_n1088# 0.016395f
C43 drain_right.n12 a_n3394_n1088# 0.063704f
C44 drain_right.n13 a_n3394_n1088# 0.53495f
C45 drain_right.t1 a_n3394_n1088# 0.016395f
C46 drain_right.t17 a_n3394_n1088# 0.016395f
C47 drain_right.n14 a_n3394_n1088# 0.063704f
C48 drain_right.n15 a_n3394_n1088# 0.263798f
C49 drain_right.t4 a_n3394_n1088# 0.016395f
C50 drain_right.t18 a_n3394_n1088# 0.016395f
C51 drain_right.n16 a_n3394_n1088# 0.063704f
C52 drain_right.n17 a_n3394_n1088# 0.263798f
C53 drain_right.t6 a_n3394_n1088# 0.016395f
C54 drain_right.t19 a_n3394_n1088# 0.016395f
C55 drain_right.n18 a_n3394_n1088# 0.063704f
C56 drain_right.n19 a_n3394_n1088# 0.263798f
C57 drain_right.t10 a_n3394_n1088# 0.016395f
C58 drain_right.t22 a_n3394_n1088# 0.016395f
C59 drain_right.n20 a_n3394_n1088# 0.063704f
C60 drain_right.n21 a_n3394_n1088# 0.447302f
C61 minus.n0 a_n3394_n1088# 0.034766f
C62 minus.n1 a_n3394_n1088# 0.007889f
C63 minus.t1 a_n3394_n1088# 0.082525f
C64 minus.n2 a_n3394_n1088# 0.034766f
C65 minus.n3 a_n3394_n1088# 0.007889f
C66 minus.t4 a_n3394_n1088# 0.082525f
C67 minus.n4 a_n3394_n1088# 0.034766f
C68 minus.n5 a_n3394_n1088# 0.007889f
C69 minus.t5 a_n3394_n1088# 0.082525f
C70 minus.n6 a_n3394_n1088# 0.034766f
C71 minus.n7 a_n3394_n1088# 0.007889f
C72 minus.t6 a_n3394_n1088# 0.082525f
C73 minus.n8 a_n3394_n1088# 0.034766f
C74 minus.n9 a_n3394_n1088# 0.007889f
C75 minus.t11 a_n3394_n1088# 0.082525f
C76 minus.t12 a_n3394_n1088# 0.10116f
C77 minus.t0 a_n3394_n1088# 0.082525f
C78 minus.n10 a_n3394_n1088# 0.089156f
C79 minus.n11 a_n3394_n1088# 0.065257f
C80 minus.n12 a_n3394_n1088# 0.149671f
C81 minus.n13 a_n3394_n1088# 0.034766f
C82 minus.n14 a_n3394_n1088# 0.082041f
C83 minus.n15 a_n3394_n1088# 0.007889f
C84 minus.t21 a_n3394_n1088# 0.082525f
C85 minus.n16 a_n3394_n1088# 0.082041f
C86 minus.n17 a_n3394_n1088# 0.034766f
C87 minus.n18 a_n3394_n1088# 0.034766f
C88 minus.n19 a_n3394_n1088# 0.034766f
C89 minus.n20 a_n3394_n1088# 0.082041f
C90 minus.n21 a_n3394_n1088# 0.007889f
C91 minus.t22 a_n3394_n1088# 0.082525f
C92 minus.n22 a_n3394_n1088# 0.082041f
C93 minus.n23 a_n3394_n1088# 0.034766f
C94 minus.n24 a_n3394_n1088# 0.034766f
C95 minus.n25 a_n3394_n1088# 0.034766f
C96 minus.n26 a_n3394_n1088# 0.082041f
C97 minus.n27 a_n3394_n1088# 0.007889f
C98 minus.t19 a_n3394_n1088# 0.082525f
C99 minus.n28 a_n3394_n1088# 0.082041f
C100 minus.n29 a_n3394_n1088# 0.034766f
C101 minus.n30 a_n3394_n1088# 0.034766f
C102 minus.n31 a_n3394_n1088# 0.034766f
C103 minus.n32 a_n3394_n1088# 0.082041f
C104 minus.n33 a_n3394_n1088# 0.007889f
C105 minus.t17 a_n3394_n1088# 0.082525f
C106 minus.n34 a_n3394_n1088# 0.082041f
C107 minus.n35 a_n3394_n1088# 0.034766f
C108 minus.n36 a_n3394_n1088# 0.034766f
C109 minus.n37 a_n3394_n1088# 0.034766f
C110 minus.n38 a_n3394_n1088# 0.082041f
C111 minus.n39 a_n3394_n1088# 0.007889f
C112 minus.t13 a_n3394_n1088# 0.082525f
C113 minus.n40 a_n3394_n1088# 0.082363f
C114 minus.n41 a_n3394_n1088# 1.10853f
C115 minus.n42 a_n3394_n1088# 0.034766f
C116 minus.n43 a_n3394_n1088# 0.007889f
C117 minus.n44 a_n3394_n1088# 0.034766f
C118 minus.n45 a_n3394_n1088# 0.007889f
C119 minus.n46 a_n3394_n1088# 0.034766f
C120 minus.n47 a_n3394_n1088# 0.007889f
C121 minus.n48 a_n3394_n1088# 0.034766f
C122 minus.n49 a_n3394_n1088# 0.007889f
C123 minus.n50 a_n3394_n1088# 0.034766f
C124 minus.n51 a_n3394_n1088# 0.007889f
C125 minus.t3 a_n3394_n1088# 0.10116f
C126 minus.t2 a_n3394_n1088# 0.082525f
C127 minus.n52 a_n3394_n1088# 0.089156f
C128 minus.n53 a_n3394_n1088# 0.065257f
C129 minus.n54 a_n3394_n1088# 0.149671f
C130 minus.n55 a_n3394_n1088# 0.034766f
C131 minus.t8 a_n3394_n1088# 0.082525f
C132 minus.n56 a_n3394_n1088# 0.082041f
C133 minus.n57 a_n3394_n1088# 0.007889f
C134 minus.t7 a_n3394_n1088# 0.082525f
C135 minus.n58 a_n3394_n1088# 0.082041f
C136 minus.n59 a_n3394_n1088# 0.034766f
C137 minus.n60 a_n3394_n1088# 0.034766f
C138 minus.n61 a_n3394_n1088# 0.034766f
C139 minus.t10 a_n3394_n1088# 0.082525f
C140 minus.n62 a_n3394_n1088# 0.082041f
C141 minus.n63 a_n3394_n1088# 0.007889f
C142 minus.t16 a_n3394_n1088# 0.082525f
C143 minus.n64 a_n3394_n1088# 0.082041f
C144 minus.n65 a_n3394_n1088# 0.034766f
C145 minus.n66 a_n3394_n1088# 0.034766f
C146 minus.n67 a_n3394_n1088# 0.034766f
C147 minus.t14 a_n3394_n1088# 0.082525f
C148 minus.n68 a_n3394_n1088# 0.082041f
C149 minus.n69 a_n3394_n1088# 0.007889f
C150 minus.t23 a_n3394_n1088# 0.082525f
C151 minus.n70 a_n3394_n1088# 0.082041f
C152 minus.n71 a_n3394_n1088# 0.034766f
C153 minus.n72 a_n3394_n1088# 0.034766f
C154 minus.n73 a_n3394_n1088# 0.034766f
C155 minus.t20 a_n3394_n1088# 0.082525f
C156 minus.n74 a_n3394_n1088# 0.082041f
C157 minus.n75 a_n3394_n1088# 0.007889f
C158 minus.t9 a_n3394_n1088# 0.082525f
C159 minus.n76 a_n3394_n1088# 0.082041f
C160 minus.n77 a_n3394_n1088# 0.034766f
C161 minus.n78 a_n3394_n1088# 0.034766f
C162 minus.n79 a_n3394_n1088# 0.034766f
C163 minus.t18 a_n3394_n1088# 0.082525f
C164 minus.n80 a_n3394_n1088# 0.082041f
C165 minus.n81 a_n3394_n1088# 0.007889f
C166 minus.t15 a_n3394_n1088# 0.082525f
C167 minus.n82 a_n3394_n1088# 0.082363f
C168 minus.n83 a_n3394_n1088# 0.241796f
C169 minus.n84 a_n3394_n1088# 1.34998f
C170 drain_left.t4 a_n3394_n1088# 0.021759f
C171 drain_left.t3 a_n3394_n1088# 0.021759f
C172 drain_left.n0 a_n3394_n1088# 0.085879f
C173 drain_left.t8 a_n3394_n1088# 0.021759f
C174 drain_left.t7 a_n3394_n1088# 0.021759f
C175 drain_left.n1 a_n3394_n1088# 0.084549f
C176 drain_left.n2 a_n3394_n1088# 0.709989f
C177 drain_left.t15 a_n3394_n1088# 0.021759f
C178 drain_left.t18 a_n3394_n1088# 0.021759f
C179 drain_left.n3 a_n3394_n1088# 0.084549f
C180 drain_left.n4 a_n3394_n1088# 0.307457f
C181 drain_left.t13 a_n3394_n1088# 0.021759f
C182 drain_left.t12 a_n3394_n1088# 0.021759f
C183 drain_left.n5 a_n3394_n1088# 0.085879f
C184 drain_left.t1 a_n3394_n1088# 0.021759f
C185 drain_left.t5 a_n3394_n1088# 0.021759f
C186 drain_left.n6 a_n3394_n1088# 0.084549f
C187 drain_left.n7 a_n3394_n1088# 0.709989f
C188 drain_left.t19 a_n3394_n1088# 0.021759f
C189 drain_left.t0 a_n3394_n1088# 0.021759f
C190 drain_left.n8 a_n3394_n1088# 0.084549f
C191 drain_left.n9 a_n3394_n1088# 0.307457f
C192 drain_left.n10 a_n3394_n1088# 1.18541f
C193 drain_left.t16 a_n3394_n1088# 0.021759f
C194 drain_left.t6 a_n3394_n1088# 0.021759f
C195 drain_left.n11 a_n3394_n1088# 0.085879f
C196 drain_left.t21 a_n3394_n1088# 0.021759f
C197 drain_left.t11 a_n3394_n1088# 0.021759f
C198 drain_left.n12 a_n3394_n1088# 0.084549f
C199 drain_left.n13 a_n3394_n1088# 0.709989f
C200 drain_left.t17 a_n3394_n1088# 0.021759f
C201 drain_left.t9 a_n3394_n1088# 0.021759f
C202 drain_left.n14 a_n3394_n1088# 0.084549f
C203 drain_left.n15 a_n3394_n1088# 0.350115f
C204 drain_left.t22 a_n3394_n1088# 0.021759f
C205 drain_left.t14 a_n3394_n1088# 0.021759f
C206 drain_left.n16 a_n3394_n1088# 0.084549f
C207 drain_left.n17 a_n3394_n1088# 0.350115f
C208 drain_left.t2 a_n3394_n1088# 0.021759f
C209 drain_left.t20 a_n3394_n1088# 0.021759f
C210 drain_left.n18 a_n3394_n1088# 0.084549f
C211 drain_left.n19 a_n3394_n1088# 0.350115f
C212 drain_left.t10 a_n3394_n1088# 0.021759f
C213 drain_left.t23 a_n3394_n1088# 0.021759f
C214 drain_left.n20 a_n3394_n1088# 0.084549f
C215 drain_left.n21 a_n3394_n1088# 0.593662f
C216 source.t30 a_n3394_n1088# 0.164866f
C217 source.n0 a_n3394_n1088# 0.782286f
C218 source.t14 a_n3394_n1088# 0.029621f
C219 source.t22 a_n3394_n1088# 0.029621f
C220 source.n1 a_n3394_n1088# 0.096066f
C221 source.n2 a_n3394_n1088# 0.444706f
C222 source.t28 a_n3394_n1088# 0.029621f
C223 source.t17 a_n3394_n1088# 0.029621f
C224 source.n3 a_n3394_n1088# 0.096066f
C225 source.n4 a_n3394_n1088# 0.444706f
C226 source.t12 a_n3394_n1088# 0.029621f
C227 source.t26 a_n3394_n1088# 0.029621f
C228 source.n5 a_n3394_n1088# 0.096066f
C229 source.n6 a_n3394_n1088# 0.444706f
C230 source.t25 a_n3394_n1088# 0.029621f
C231 source.t19 a_n3394_n1088# 0.029621f
C232 source.n7 a_n3394_n1088# 0.096066f
C233 source.n8 a_n3394_n1088# 0.444706f
C234 source.t32 a_n3394_n1088# 0.029621f
C235 source.t21 a_n3394_n1088# 0.029621f
C236 source.n9 a_n3394_n1088# 0.096066f
C237 source.n10 a_n3394_n1088# 0.444706f
C238 source.t31 a_n3394_n1088# 0.164866f
C239 source.n11 a_n3394_n1088# 0.406191f
C240 source.t8 a_n3394_n1088# 0.164866f
C241 source.n12 a_n3394_n1088# 0.406191f
C242 source.t40 a_n3394_n1088# 0.029621f
C243 source.t2 a_n3394_n1088# 0.029621f
C244 source.n13 a_n3394_n1088# 0.096066f
C245 source.n14 a_n3394_n1088# 0.444706f
C246 source.t1 a_n3394_n1088# 0.029621f
C247 source.t34 a_n3394_n1088# 0.029621f
C248 source.n15 a_n3394_n1088# 0.096066f
C249 source.n16 a_n3394_n1088# 0.444706f
C250 source.t46 a_n3394_n1088# 0.029621f
C251 source.t38 a_n3394_n1088# 0.029621f
C252 source.n17 a_n3394_n1088# 0.096066f
C253 source.n18 a_n3394_n1088# 0.444706f
C254 source.t0 a_n3394_n1088# 0.029621f
C255 source.t44 a_n3394_n1088# 0.029621f
C256 source.n19 a_n3394_n1088# 0.096066f
C257 source.n20 a_n3394_n1088# 0.444706f
C258 source.t7 a_n3394_n1088# 0.029621f
C259 source.t45 a_n3394_n1088# 0.029621f
C260 source.n21 a_n3394_n1088# 0.096066f
C261 source.n22 a_n3394_n1088# 0.444706f
C262 source.t47 a_n3394_n1088# 0.164866f
C263 source.n23 a_n3394_n1088# 1.09157f
C264 source.t15 a_n3394_n1088# 0.164866f
C265 source.n24 a_n3394_n1088# 1.09157f
C266 source.t11 a_n3394_n1088# 0.029621f
C267 source.t18 a_n3394_n1088# 0.029621f
C268 source.n25 a_n3394_n1088# 0.096065f
C269 source.n26 a_n3394_n1088# 0.444706f
C270 source.t20 a_n3394_n1088# 0.029621f
C271 source.t27 a_n3394_n1088# 0.029621f
C272 source.n27 a_n3394_n1088# 0.096065f
C273 source.n28 a_n3394_n1088# 0.444706f
C274 source.t24 a_n3394_n1088# 0.029621f
C275 source.t10 a_n3394_n1088# 0.029621f
C276 source.n29 a_n3394_n1088# 0.096065f
C277 source.n30 a_n3394_n1088# 0.444706f
C278 source.t16 a_n3394_n1088# 0.029621f
C279 source.t33 a_n3394_n1088# 0.029621f
C280 source.n31 a_n3394_n1088# 0.096065f
C281 source.n32 a_n3394_n1088# 0.444706f
C282 source.t13 a_n3394_n1088# 0.029621f
C283 source.t23 a_n3394_n1088# 0.029621f
C284 source.n33 a_n3394_n1088# 0.096065f
C285 source.n34 a_n3394_n1088# 0.444706f
C286 source.t29 a_n3394_n1088# 0.164866f
C287 source.n35 a_n3394_n1088# 0.406191f
C288 source.t42 a_n3394_n1088# 0.164866f
C289 source.n36 a_n3394_n1088# 0.406191f
C290 source.t37 a_n3394_n1088# 0.029621f
C291 source.t41 a_n3394_n1088# 0.029621f
C292 source.n37 a_n3394_n1088# 0.096065f
C293 source.n38 a_n3394_n1088# 0.444706f
C294 source.t36 a_n3394_n1088# 0.029621f
C295 source.t35 a_n3394_n1088# 0.029621f
C296 source.n39 a_n3394_n1088# 0.096065f
C297 source.n40 a_n3394_n1088# 0.444706f
C298 source.t39 a_n3394_n1088# 0.029621f
C299 source.t43 a_n3394_n1088# 0.029621f
C300 source.n41 a_n3394_n1088# 0.096065f
C301 source.n42 a_n3394_n1088# 0.444706f
C302 source.t3 a_n3394_n1088# 0.029621f
C303 source.t5 a_n3394_n1088# 0.029621f
C304 source.n43 a_n3394_n1088# 0.096065f
C305 source.n44 a_n3394_n1088# 0.444706f
C306 source.t9 a_n3394_n1088# 0.029621f
C307 source.t4 a_n3394_n1088# 0.029621f
C308 source.n45 a_n3394_n1088# 0.096065f
C309 source.n46 a_n3394_n1088# 0.444706f
C310 source.t6 a_n3394_n1088# 0.164866f
C311 source.n47 a_n3394_n1088# 0.650701f
C312 source.n48 a_n3394_n1088# 0.77681f
C313 plus.n0 a_n3394_n1088# 0.04466f
C314 plus.t0 a_n3394_n1088# 0.106008f
C315 plus.t13 a_n3394_n1088# 0.106008f
C316 plus.n1 a_n3394_n1088# 0.04466f
C317 plus.t3 a_n3394_n1088# 0.106008f
C318 plus.n2 a_n3394_n1088# 0.105387f
C319 plus.n3 a_n3394_n1088# 0.04466f
C320 plus.t21 a_n3394_n1088# 0.106008f
C321 plus.t9 a_n3394_n1088# 0.106008f
C322 plus.n4 a_n3394_n1088# 0.105387f
C323 plus.n5 a_n3394_n1088# 0.04466f
C324 plus.t1 a_n3394_n1088# 0.106008f
C325 plus.t14 a_n3394_n1088# 0.106008f
C326 plus.n6 a_n3394_n1088# 0.105387f
C327 plus.n7 a_n3394_n1088# 0.04466f
C328 plus.t6 a_n3394_n1088# 0.106008f
C329 plus.t12 a_n3394_n1088# 0.106008f
C330 plus.n8 a_n3394_n1088# 0.105387f
C331 plus.n9 a_n3394_n1088# 0.04466f
C332 plus.t2 a_n3394_n1088# 0.106008f
C333 plus.t17 a_n3394_n1088# 0.106008f
C334 plus.n10 a_n3394_n1088# 0.114526f
C335 plus.t7 a_n3394_n1088# 0.129946f
C336 plus.n11 a_n3394_n1088# 0.083827f
C337 plus.n12 a_n3394_n1088# 0.192262f
C338 plus.n13 a_n3394_n1088# 0.010134f
C339 plus.n14 a_n3394_n1088# 0.105387f
C340 plus.n15 a_n3394_n1088# 0.010134f
C341 plus.n16 a_n3394_n1088# 0.04466f
C342 plus.n17 a_n3394_n1088# 0.04466f
C343 plus.n18 a_n3394_n1088# 0.04466f
C344 plus.n19 a_n3394_n1088# 0.010134f
C345 plus.n20 a_n3394_n1088# 0.105387f
C346 plus.n21 a_n3394_n1088# 0.010134f
C347 plus.n22 a_n3394_n1088# 0.04466f
C348 plus.n23 a_n3394_n1088# 0.04466f
C349 plus.n24 a_n3394_n1088# 0.04466f
C350 plus.n25 a_n3394_n1088# 0.010134f
C351 plus.n26 a_n3394_n1088# 0.105387f
C352 plus.n27 a_n3394_n1088# 0.010134f
C353 plus.n28 a_n3394_n1088# 0.04466f
C354 plus.n29 a_n3394_n1088# 0.04466f
C355 plus.n30 a_n3394_n1088# 0.04466f
C356 plus.n31 a_n3394_n1088# 0.010134f
C357 plus.n32 a_n3394_n1088# 0.105387f
C358 plus.n33 a_n3394_n1088# 0.010134f
C359 plus.n34 a_n3394_n1088# 0.04466f
C360 plus.n35 a_n3394_n1088# 0.04466f
C361 plus.n36 a_n3394_n1088# 0.04466f
C362 plus.n37 a_n3394_n1088# 0.010134f
C363 plus.n38 a_n3394_n1088# 0.105387f
C364 plus.n39 a_n3394_n1088# 0.010134f
C365 plus.n40 a_n3394_n1088# 0.1058f
C366 plus.n41 a_n3394_n1088# 0.32583f
C367 plus.n42 a_n3394_n1088# 0.04466f
C368 plus.t19 a_n3394_n1088# 0.106008f
C369 plus.n43 a_n3394_n1088# 0.04466f
C370 plus.t20 a_n3394_n1088# 0.106008f
C371 plus.t15 a_n3394_n1088# 0.106008f
C372 plus.n44 a_n3394_n1088# 0.105387f
C373 plus.n45 a_n3394_n1088# 0.04466f
C374 plus.t16 a_n3394_n1088# 0.106008f
C375 plus.t8 a_n3394_n1088# 0.106008f
C376 plus.n46 a_n3394_n1088# 0.105387f
C377 plus.n47 a_n3394_n1088# 0.04466f
C378 plus.t5 a_n3394_n1088# 0.106008f
C379 plus.t4 a_n3394_n1088# 0.106008f
C380 plus.n48 a_n3394_n1088# 0.105387f
C381 plus.n49 a_n3394_n1088# 0.04466f
C382 plus.t23 a_n3394_n1088# 0.106008f
C383 plus.t22 a_n3394_n1088# 0.106008f
C384 plus.n50 a_n3394_n1088# 0.105387f
C385 plus.n51 a_n3394_n1088# 0.04466f
C386 plus.t18 a_n3394_n1088# 0.106008f
C387 plus.t10 a_n3394_n1088# 0.106008f
C388 plus.n52 a_n3394_n1088# 0.114526f
C389 plus.t11 a_n3394_n1088# 0.129946f
C390 plus.n53 a_n3394_n1088# 0.083827f
C391 plus.n54 a_n3394_n1088# 0.192262f
C392 plus.n55 a_n3394_n1088# 0.010134f
C393 plus.n56 a_n3394_n1088# 0.105387f
C394 plus.n57 a_n3394_n1088# 0.010134f
C395 plus.n58 a_n3394_n1088# 0.04466f
C396 plus.n59 a_n3394_n1088# 0.04466f
C397 plus.n60 a_n3394_n1088# 0.04466f
C398 plus.n61 a_n3394_n1088# 0.010134f
C399 plus.n62 a_n3394_n1088# 0.105387f
C400 plus.n63 a_n3394_n1088# 0.010134f
C401 plus.n64 a_n3394_n1088# 0.04466f
C402 plus.n65 a_n3394_n1088# 0.04466f
C403 plus.n66 a_n3394_n1088# 0.04466f
C404 plus.n67 a_n3394_n1088# 0.010134f
C405 plus.n68 a_n3394_n1088# 0.105387f
C406 plus.n69 a_n3394_n1088# 0.010134f
C407 plus.n70 a_n3394_n1088# 0.04466f
C408 plus.n71 a_n3394_n1088# 0.04466f
C409 plus.n72 a_n3394_n1088# 0.04466f
C410 plus.n73 a_n3394_n1088# 0.010134f
C411 plus.n74 a_n3394_n1088# 0.105387f
C412 plus.n75 a_n3394_n1088# 0.010134f
C413 plus.n76 a_n3394_n1088# 0.04466f
C414 plus.n77 a_n3394_n1088# 0.04466f
C415 plus.n78 a_n3394_n1088# 0.04466f
C416 plus.n79 a_n3394_n1088# 0.010134f
C417 plus.n80 a_n3394_n1088# 0.105387f
C418 plus.n81 a_n3394_n1088# 0.010134f
C419 plus.n82 a_n3394_n1088# 0.1058f
C420 plus.n83 a_n3394_n1088# 1.37028f
.ends

