* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right.t5 minus.t0 source.t7 a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X1 a_n1236_n1088# a_n1236_n1088# a_n1236_n1088# a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=3.8 ps=23.6 w=1 l=0.15
X2 a_n1236_n1088# a_n1236_n1088# a_n1236_n1088# a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X3 source.t3 plus.t0 drain_left.t5 a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X4 a_n1236_n1088# a_n1236_n1088# a_n1236_n1088# a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X5 source.t10 minus.t1 drain_right.t4 a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X6 a_n1236_n1088# a_n1236_n1088# a_n1236_n1088# a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X7 drain_left.t4 plus.t1 source.t2 a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X8 source.t6 minus.t2 drain_right.t3 a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X9 drain_right.t2 minus.t3 source.t8 a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X10 drain_right.t1 minus.t4 source.t9 a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
X11 drain_left.t3 plus.t2 source.t0 a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
X12 drain_right.t0 minus.t5 source.t11 a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
X13 drain_left.t2 plus.t3 source.t5 a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.475 ps=2.95 w=1 l=0.15
X14 source.t1 plus.t4 drain_left.t1 a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X15 drain_left.t0 plus.t5 source.t4 a_n1236_n1088# sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.25 ps=1.5 w=1 l=0.15
R0 minus.n2 minus.t5 427.959
R1 minus.n0 minus.t3 427.959
R2 minus.n6 minus.t0 427.959
R3 minus.n4 minus.t4 427.959
R4 minus.n1 minus.t2 369.534
R5 minus.n5 minus.t1 369.534
R6 minus.n3 minus.n0 161.489
R7 minus.n7 minus.n4 161.489
R8 minus.n3 minus.n2 161.3
R9 minus.n7 minus.n6 161.3
R10 minus.n2 minus.n1 36.5157
R11 minus.n1 minus.n0 36.5157
R12 minus.n5 minus.n4 36.5157
R13 minus.n6 minus.n5 36.5157
R14 minus.n8 minus.n3 25.5213
R15 minus.n8 minus.n7 6.55164
R16 minus minus.n8 0.188
R17 source.n0 source.t5 253.454
R18 source.n3 source.t8 253.454
R19 source.n11 source.t7 253.453
R20 source.n8 source.t2 253.453
R21 source.n2 source.n1 223.454
R22 source.n5 source.n4 223.454
R23 source.n10 source.n9 223.453
R24 source.n7 source.n6 223.453
R25 source.n9 source.t9 30.0005
R26 source.n9 source.t10 30.0005
R27 source.n6 source.t4 30.0005
R28 source.n6 source.t3 30.0005
R29 source.n1 source.t0 30.0005
R30 source.n1 source.t1 30.0005
R31 source.n4 source.t11 30.0005
R32 source.n4 source.t6 30.0005
R33 source.n7 source.n5 14.0751
R34 source.n12 source.n0 7.97163
R35 source.n12 source.n11 5.5436
R36 source.n3 source.n2 0.7505
R37 source.n10 source.n8 0.7505
R38 source.n5 source.n3 0.560845
R39 source.n2 source.n0 0.560845
R40 source.n8 source.n7 0.560845
R41 source.n11 source.n10 0.560845
R42 source source.n12 0.188
R43 drain_right.n1 drain_right.t1 270.497
R44 drain_right.n3 drain_right.t0 270.132
R45 drain_right.n3 drain_right.n2 240.694
R46 drain_right.n1 drain_right.n0 240.216
R47 drain_right.n0 drain_right.t4 30.0005
R48 drain_right.n0 drain_right.t5 30.0005
R49 drain_right.n2 drain_right.t3 30.0005
R50 drain_right.n2 drain_right.t2 30.0005
R51 drain_right drain_right.n1 20.0215
R52 drain_right drain_right.n3 5.93339
R53 plus.n0 plus.t2 427.959
R54 plus.n2 plus.t3 427.959
R55 plus.n4 plus.t1 427.959
R56 plus.n6 plus.t5 427.959
R57 plus.n1 plus.t4 369.534
R58 plus.n5 plus.t0 369.534
R59 plus.n3 plus.n0 161.489
R60 plus.n7 plus.n4 161.489
R61 plus.n3 plus.n2 161.3
R62 plus.n7 plus.n6 161.3
R63 plus.n1 plus.n0 36.5157
R64 plus.n2 plus.n1 36.5157
R65 plus.n6 plus.n5 36.5157
R66 plus.n5 plus.n4 36.5157
R67 plus plus.n7 23.5691
R68 plus plus.n3 8.02891
R69 drain_left.n3 drain_left.t3 270.693
R70 drain_left.n1 drain_left.t0 270.497
R71 drain_left.n1 drain_left.n0 240.216
R72 drain_left.n3 drain_left.n2 240.132
R73 drain_left.n0 drain_left.t5 30.0005
R74 drain_left.n0 drain_left.t4 30.0005
R75 drain_left.n2 drain_left.t1 30.0005
R76 drain_left.n2 drain_left.t2 30.0005
R77 drain_left drain_left.n1 20.5747
R78 drain_left drain_left.n3 6.21356
C0 drain_left drain_right 0.571741f
C1 drain_left source 2.72315f
C2 drain_right plus 0.277546f
C3 minus drain_left 0.177869f
C4 source plus 0.540184f
C5 minus plus 2.64701f
C6 source drain_right 2.72054f
C7 minus drain_right 0.429507f
C8 minus source 0.526267f
C9 drain_left plus 0.545125f
C10 drain_right a_n1236_n1088# 2.741291f
C11 drain_left a_n1236_n1088# 2.892856f
C12 source a_n1236_n1088# 1.957489f
C13 minus a_n1236_n1088# 3.622617f
C14 plus a_n1236_n1088# 4.43168f
C15 drain_left.t0 a_n1236_n1088# 0.109142f
C16 drain_left.t5 a_n1236_n1088# 0.023697f
C17 drain_left.t4 a_n1236_n1088# 0.023697f
C18 drain_left.n0 a_n1236_n1088# 0.076955f
C19 drain_left.n1 a_n1236_n1088# 0.788788f
C20 drain_left.t3 a_n1236_n1088# 0.109296f
C21 drain_left.t1 a_n1236_n1088# 0.023697f
C22 drain_left.t2 a_n1236_n1088# 0.023697f
C23 drain_left.n2 a_n1236_n1088# 0.076887f
C24 drain_left.n3 a_n1236_n1088# 0.567517f
C25 plus.t2 a_n1236_n1088# 0.02403f
C26 plus.n0 a_n1236_n1088# 0.043339f
C27 plus.t4 a_n1236_n1088# 0.020104f
C28 plus.n1 a_n1236_n1088# 0.027415f
C29 plus.t3 a_n1236_n1088# 0.02403f
C30 plus.n2 a_n1236_n1088# 0.043273f
C31 plus.n3 a_n1236_n1088# 0.359118f
C32 plus.t1 a_n1236_n1088# 0.02403f
C33 plus.n4 a_n1236_n1088# 0.043339f
C34 plus.t5 a_n1236_n1088# 0.02403f
C35 plus.t0 a_n1236_n1088# 0.020104f
C36 plus.n5 a_n1236_n1088# 0.027415f
C37 plus.n6 a_n1236_n1088# 0.043273f
C38 plus.n7 a_n1236_n1088# 0.887899f
C39 drain_right.t1 a_n1236_n1088# 0.112364f
C40 drain_right.t4 a_n1236_n1088# 0.024397f
C41 drain_right.t5 a_n1236_n1088# 0.024397f
C42 drain_right.n0 a_n1236_n1088# 0.079227f
C43 drain_right.n1 a_n1236_n1088# 0.772536f
C44 drain_right.t3 a_n1236_n1088# 0.024397f
C45 drain_right.t2 a_n1236_n1088# 0.024397f
C46 drain_right.n2 a_n1236_n1088# 0.079679f
C47 drain_right.t0 a_n1236_n1088# 0.112112f
C48 drain_right.n3 a_n1236_n1088# 0.593064f
C49 source.t5 a_n1236_n1088# 0.135898f
C50 source.n0 a_n1236_n1088# 0.519283f
C51 source.t0 a_n1236_n1088# 0.032419f
C52 source.t1 a_n1236_n1088# 0.032419f
C53 source.n1 a_n1236_n1088# 0.091437f
C54 source.n2 a_n1236_n1088# 0.280615f
C55 source.t8 a_n1236_n1088# 0.135898f
C56 source.n3 a_n1236_n1088# 0.294508f
C57 source.t11 a_n1236_n1088# 0.032419f
C58 source.t6 a_n1236_n1088# 0.032419f
C59 source.n4 a_n1236_n1088# 0.091437f
C60 source.n5 a_n1236_n1088# 0.771554f
C61 source.t4 a_n1236_n1088# 0.032419f
C62 source.t3 a_n1236_n1088# 0.032419f
C63 source.n6 a_n1236_n1088# 0.091437f
C64 source.n7 a_n1236_n1088# 0.771554f
C65 source.t2 a_n1236_n1088# 0.135898f
C66 source.n8 a_n1236_n1088# 0.294508f
C67 source.t9 a_n1236_n1088# 0.032419f
C68 source.t10 a_n1236_n1088# 0.032419f
C69 source.n9 a_n1236_n1088# 0.091437f
C70 source.n10 a_n1236_n1088# 0.280615f
C71 source.t7 a_n1236_n1088# 0.135898f
C72 source.n11 a_n1236_n1088# 0.424111f
C73 source.n12 a_n1236_n1088# 0.548982f
C74 minus.t3 a_n1236_n1088# 0.023244f
C75 minus.n0 a_n1236_n1088# 0.041921f
C76 minus.t5 a_n1236_n1088# 0.023244f
C77 minus.t2 a_n1236_n1088# 0.019447f
C78 minus.n1 a_n1236_n1088# 0.026518f
C79 minus.n2 a_n1236_n1088# 0.041858f
C80 minus.n3 a_n1236_n1088# 0.876042f
C81 minus.t4 a_n1236_n1088# 0.023244f
C82 minus.n4 a_n1236_n1088# 0.041921f
C83 minus.t1 a_n1236_n1088# 0.019447f
C84 minus.n5 a_n1236_n1088# 0.026518f
C85 minus.t0 a_n1236_n1088# 0.023244f
C86 minus.n6 a_n1236_n1088# 0.041858f
C87 minus.n7 a_n1236_n1088# 0.333711f
C88 minus.n8 a_n1236_n1088# 1.01017f
.ends

