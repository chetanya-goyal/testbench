* NGSPICE file created from diffpair578.ext - technology: sky130A

.subckt diffpair578 minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t34 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X1 drain_left.t18 plus.t1 source.t36 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X2 drain_right.t19 minus.t0 source.t7 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X3 drain_right.t18 minus.t1 source.t10 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X4 source.t32 plus.t2 drain_left.t17 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X5 source.t31 plus.t3 drain_left.t16 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X6 drain_left.t15 plus.t4 source.t23 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X7 source.t12 minus.t2 drain_right.t17 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X8 source.t16 minus.t3 drain_right.t16 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X9 source.t9 minus.t4 drain_right.t15 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X10 source.t13 minus.t5 drain_right.t14 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X11 drain_left.t14 plus.t5 source.t27 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X12 drain_right.t13 minus.t6 source.t14 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X13 source.t17 minus.t7 drain_right.t12 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X14 drain_right.t11 minus.t8 source.t2 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X15 drain_right.t10 minus.t9 source.t5 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X16 drain_left.t13 plus.t6 source.t22 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X17 source.t30 plus.t7 drain_left.t12 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X18 a_n1882_n4888# a_n1882_n4888# a_n1882_n4888# a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.2
X19 drain_right.t9 minus.t10 source.t1 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X20 drain_right.t8 minus.t11 source.t4 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X21 source.t11 minus.t12 drain_right.t7 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X22 drain_right.t6 minus.t13 source.t15 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X23 source.t8 minus.t14 drain_right.t5 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X24 source.t21 plus.t8 drain_left.t11 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X25 drain_right.t4 minus.t15 source.t6 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X26 drain_right.t3 minus.t16 source.t38 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X27 source.t39 minus.t17 drain_right.t2 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X28 drain_left.t10 plus.t9 source.t28 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X29 source.t33 plus.t10 drain_left.t9 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X30 a_n1882_n4888# a_n1882_n4888# a_n1882_n4888# a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X31 a_n1882_n4888# a_n1882_n4888# a_n1882_n4888# a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X32 source.t26 plus.t11 drain_left.t8 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X33 drain_left.t7 plus.t12 source.t29 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X34 source.t20 plus.t13 drain_left.t6 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X35 source.t3 minus.t18 drain_right.t1 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X36 source.t0 minus.t19 drain_right.t0 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X37 source.t19 plus.t14 drain_left.t5 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X38 source.t35 plus.t15 drain_left.t4 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X39 drain_left.t3 plus.t16 source.t37 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X40 drain_left.t2 plus.t17 source.t24 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X41 source.t18 plus.t18 drain_left.t1 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X42 a_n1882_n4888# a_n1882_n4888# a_n1882_n4888# a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X43 drain_left.t0 plus.t19 source.t25 a_n1882_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
R0 plus.n5 plus.t7 2622.88
R1 plus.n23 plus.t5 2622.88
R2 plus.n30 plus.t0 2622.88
R3 plus.n48 plus.t8 2622.88
R4 plus.n6 plus.t4 2566.65
R5 plus.n8 plus.t18 2566.65
R6 plus.n3 plus.t12 2566.65
R7 plus.n13 plus.t11 2566.65
R8 plus.n15 plus.t6 2566.65
R9 plus.n1 plus.t3 2566.65
R10 plus.n20 plus.t17 2566.65
R11 plus.n22 plus.t10 2566.65
R12 plus.n31 plus.t2 2566.65
R13 plus.n33 plus.t1 2566.65
R14 plus.n28 plus.t14 2566.65
R15 plus.n38 plus.t19 2566.65
R16 plus.n40 plus.t15 2566.65
R17 plus.n26 plus.t16 2566.65
R18 plus.n45 plus.t13 2566.65
R19 plus.n47 plus.t9 2566.65
R20 plus.n5 plus.n4 161.489
R21 plus.n30 plus.n29 161.489
R22 plus.n7 plus.n4 161.3
R23 plus.n10 plus.n9 161.3
R24 plus.n12 plus.n11 161.3
R25 plus.n14 plus.n2 161.3
R26 plus.n17 plus.n16 161.3
R27 plus.n19 plus.n18 161.3
R28 plus.n21 plus.n0 161.3
R29 plus.n24 plus.n23 161.3
R30 plus.n32 plus.n29 161.3
R31 plus.n35 plus.n34 161.3
R32 plus.n37 plus.n36 161.3
R33 plus.n39 plus.n27 161.3
R34 plus.n42 plus.n41 161.3
R35 plus.n44 plus.n43 161.3
R36 plus.n46 plus.n25 161.3
R37 plus.n49 plus.n48 161.3
R38 plus.n7 plus.n6 51.852
R39 plus.n22 plus.n21 51.852
R40 plus.n47 plus.n46 51.852
R41 plus.n32 plus.n31 51.852
R42 plus.n9 plus.n8 47.4702
R43 plus.n20 plus.n19 47.4702
R44 plus.n45 plus.n44 47.4702
R45 plus.n34 plus.n33 47.4702
R46 plus.n12 plus.n3 43.0884
R47 plus.n16 plus.n1 43.0884
R48 plus.n41 plus.n26 43.0884
R49 plus.n37 plus.n28 43.0884
R50 plus.n14 plus.n13 38.7066
R51 plus.n15 plus.n14 38.7066
R52 plus.n40 plus.n39 38.7066
R53 plus.n39 plus.n38 38.7066
R54 plus.n13 plus.n12 34.3247
R55 plus.n16 plus.n15 34.3247
R56 plus.n41 plus.n40 34.3247
R57 plus.n38 plus.n37 34.3247
R58 plus plus.n49 33.1392
R59 plus.n9 plus.n3 29.9429
R60 plus.n19 plus.n1 29.9429
R61 plus.n44 plus.n26 29.9429
R62 plus.n34 plus.n28 29.9429
R63 plus.n8 plus.n7 25.5611
R64 plus.n21 plus.n20 25.5611
R65 plus.n46 plus.n45 25.5611
R66 plus.n33 plus.n32 25.5611
R67 plus.n6 plus.n5 21.1793
R68 plus.n23 plus.n22 21.1793
R69 plus.n48 plus.n47 21.1793
R70 plus.n31 plus.n30 21.1793
R71 plus plus.n24 15.152
R72 plus.n10 plus.n4 0.189894
R73 plus.n11 plus.n10 0.189894
R74 plus.n11 plus.n2 0.189894
R75 plus.n17 plus.n2 0.189894
R76 plus.n18 plus.n17 0.189894
R77 plus.n18 plus.n0 0.189894
R78 plus.n24 plus.n0 0.189894
R79 plus.n49 plus.n25 0.189894
R80 plus.n43 plus.n25 0.189894
R81 plus.n43 plus.n42 0.189894
R82 plus.n42 plus.n27 0.189894
R83 plus.n36 plus.n27 0.189894
R84 plus.n36 plus.n35 0.189894
R85 plus.n35 plus.n29 0.189894
R86 source.n0 source.t27 44.1297
R87 source.n9 source.t30 44.1296
R88 source.n10 source.t6 44.1296
R89 source.n19 source.t17 44.1296
R90 source.n39 source.t14 44.1295
R91 source.n30 source.t9 44.1295
R92 source.n29 source.t34 44.1295
R93 source.n20 source.t21 44.1295
R94 source.n2 source.n1 43.1397
R95 source.n4 source.n3 43.1397
R96 source.n6 source.n5 43.1397
R97 source.n8 source.n7 43.1397
R98 source.n12 source.n11 43.1397
R99 source.n14 source.n13 43.1397
R100 source.n16 source.n15 43.1397
R101 source.n18 source.n17 43.1397
R102 source.n38 source.n37 43.1396
R103 source.n36 source.n35 43.1396
R104 source.n34 source.n33 43.1396
R105 source.n32 source.n31 43.1396
R106 source.n28 source.n27 43.1396
R107 source.n26 source.n25 43.1396
R108 source.n24 source.n23 43.1396
R109 source.n22 source.n21 43.1396
R110 source.n20 source.n19 27.8052
R111 source.n40 source.n0 22.3138
R112 source.n40 source.n39 5.49188
R113 source.n37 source.t1 0.9905
R114 source.n37 source.t11 0.9905
R115 source.n35 source.t4 0.9905
R116 source.n35 source.t8 0.9905
R117 source.n33 source.t2 0.9905
R118 source.n33 source.t39 0.9905
R119 source.n31 source.t5 0.9905
R120 source.n31 source.t12 0.9905
R121 source.n27 source.t36 0.9905
R122 source.n27 source.t32 0.9905
R123 source.n25 source.t25 0.9905
R124 source.n25 source.t19 0.9905
R125 source.n23 source.t37 0.9905
R126 source.n23 source.t35 0.9905
R127 source.n21 source.t28 0.9905
R128 source.n21 source.t20 0.9905
R129 source.n1 source.t24 0.9905
R130 source.n1 source.t33 0.9905
R131 source.n3 source.t22 0.9905
R132 source.n3 source.t31 0.9905
R133 source.n5 source.t29 0.9905
R134 source.n5 source.t26 0.9905
R135 source.n7 source.t23 0.9905
R136 source.n7 source.t18 0.9905
R137 source.n11 source.t7 0.9905
R138 source.n11 source.t13 0.9905
R139 source.n13 source.t38 0.9905
R140 source.n13 source.t3 0.9905
R141 source.n15 source.t10 0.9905
R142 source.n15 source.t16 0.9905
R143 source.n17 source.t15 0.9905
R144 source.n17 source.t0 0.9905
R145 source.n10 source.n9 0.470328
R146 source.n30 source.n29 0.470328
R147 source.n19 source.n18 0.457397
R148 source.n18 source.n16 0.457397
R149 source.n16 source.n14 0.457397
R150 source.n14 source.n12 0.457397
R151 source.n12 source.n10 0.457397
R152 source.n9 source.n8 0.457397
R153 source.n8 source.n6 0.457397
R154 source.n6 source.n4 0.457397
R155 source.n4 source.n2 0.457397
R156 source.n2 source.n0 0.457397
R157 source.n22 source.n20 0.457397
R158 source.n24 source.n22 0.457397
R159 source.n26 source.n24 0.457397
R160 source.n28 source.n26 0.457397
R161 source.n29 source.n28 0.457397
R162 source.n32 source.n30 0.457397
R163 source.n34 source.n32 0.457397
R164 source.n36 source.n34 0.457397
R165 source.n38 source.n36 0.457397
R166 source.n39 source.n38 0.457397
R167 source source.n40 0.188
R168 drain_left.n10 drain_left.n8 60.2753
R169 drain_left.n6 drain_left.n4 60.2753
R170 drain_left.n2 drain_left.n0 60.2753
R171 drain_left.n16 drain_left.n15 59.8185
R172 drain_left.n14 drain_left.n13 59.8185
R173 drain_left.n12 drain_left.n11 59.8185
R174 drain_left.n10 drain_left.n9 59.8185
R175 drain_left.n7 drain_left.n3 59.8184
R176 drain_left.n6 drain_left.n5 59.8184
R177 drain_left.n2 drain_left.n1 59.8184
R178 drain_left drain_left.n7 37.0829
R179 drain_left drain_left.n16 6.11011
R180 drain_left.n3 drain_left.t4 0.9905
R181 drain_left.n3 drain_left.t0 0.9905
R182 drain_left.n4 drain_left.t17 0.9905
R183 drain_left.n4 drain_left.t19 0.9905
R184 drain_left.n5 drain_left.t5 0.9905
R185 drain_left.n5 drain_left.t18 0.9905
R186 drain_left.n1 drain_left.t6 0.9905
R187 drain_left.n1 drain_left.t3 0.9905
R188 drain_left.n0 drain_left.t11 0.9905
R189 drain_left.n0 drain_left.t10 0.9905
R190 drain_left.n15 drain_left.t9 0.9905
R191 drain_left.n15 drain_left.t14 0.9905
R192 drain_left.n13 drain_left.t16 0.9905
R193 drain_left.n13 drain_left.t2 0.9905
R194 drain_left.n11 drain_left.t8 0.9905
R195 drain_left.n11 drain_left.t13 0.9905
R196 drain_left.n9 drain_left.t1 0.9905
R197 drain_left.n9 drain_left.t7 0.9905
R198 drain_left.n8 drain_left.t12 0.9905
R199 drain_left.n8 drain_left.t15 0.9905
R200 drain_left.n12 drain_left.n10 0.457397
R201 drain_left.n14 drain_left.n12 0.457397
R202 drain_left.n16 drain_left.n14 0.457397
R203 drain_left.n7 drain_left.n6 0.402051
R204 drain_left.n7 drain_left.n2 0.402051
R205 minus.n23 minus.t7 2622.88
R206 minus.n5 minus.t15 2622.88
R207 minus.n48 minus.t6 2622.88
R208 minus.n30 minus.t4 2622.88
R209 minus.n22 minus.t13 2566.65
R210 minus.n20 minus.t19 2566.65
R211 minus.n1 minus.t1 2566.65
R212 minus.n15 minus.t3 2566.65
R213 minus.n13 minus.t16 2566.65
R214 minus.n3 minus.t18 2566.65
R215 minus.n8 minus.t0 2566.65
R216 minus.n6 minus.t5 2566.65
R217 minus.n47 minus.t12 2566.65
R218 minus.n45 minus.t10 2566.65
R219 minus.n26 minus.t14 2566.65
R220 minus.n40 minus.t11 2566.65
R221 minus.n38 minus.t17 2566.65
R222 minus.n28 minus.t8 2566.65
R223 minus.n33 minus.t2 2566.65
R224 minus.n31 minus.t9 2566.65
R225 minus.n5 minus.n4 161.489
R226 minus.n30 minus.n29 161.489
R227 minus.n24 minus.n23 161.3
R228 minus.n21 minus.n0 161.3
R229 minus.n19 minus.n18 161.3
R230 minus.n17 minus.n16 161.3
R231 minus.n14 minus.n2 161.3
R232 minus.n12 minus.n11 161.3
R233 minus.n10 minus.n9 161.3
R234 minus.n7 minus.n4 161.3
R235 minus.n49 minus.n48 161.3
R236 minus.n46 minus.n25 161.3
R237 minus.n44 minus.n43 161.3
R238 minus.n42 minus.n41 161.3
R239 minus.n39 minus.n27 161.3
R240 minus.n37 minus.n36 161.3
R241 minus.n35 minus.n34 161.3
R242 minus.n32 minus.n29 161.3
R243 minus.n22 minus.n21 51.852
R244 minus.n7 minus.n6 51.852
R245 minus.n32 minus.n31 51.852
R246 minus.n47 minus.n46 51.852
R247 minus.n20 minus.n19 47.4702
R248 minus.n9 minus.n8 47.4702
R249 minus.n34 minus.n33 47.4702
R250 minus.n45 minus.n44 47.4702
R251 minus.n16 minus.n1 43.0884
R252 minus.n12 minus.n3 43.0884
R253 minus.n37 minus.n28 43.0884
R254 minus.n41 minus.n26 43.0884
R255 minus.n50 minus.n24 42.2884
R256 minus.n15 minus.n14 38.7066
R257 minus.n14 minus.n13 38.7066
R258 minus.n39 minus.n38 38.7066
R259 minus.n40 minus.n39 38.7066
R260 minus.n16 minus.n15 34.3247
R261 minus.n13 minus.n12 34.3247
R262 minus.n38 minus.n37 34.3247
R263 minus.n41 minus.n40 34.3247
R264 minus.n19 minus.n1 29.9429
R265 minus.n9 minus.n3 29.9429
R266 minus.n34 minus.n28 29.9429
R267 minus.n44 minus.n26 29.9429
R268 minus.n21 minus.n20 25.5611
R269 minus.n8 minus.n7 25.5611
R270 minus.n33 minus.n32 25.5611
R271 minus.n46 minus.n45 25.5611
R272 minus.n23 minus.n22 21.1793
R273 minus.n6 minus.n5 21.1793
R274 minus.n31 minus.n30 21.1793
R275 minus.n48 minus.n47 21.1793
R276 minus.n50 minus.n49 6.47777
R277 minus.n24 minus.n0 0.189894
R278 minus.n18 minus.n0 0.189894
R279 minus.n18 minus.n17 0.189894
R280 minus.n17 minus.n2 0.189894
R281 minus.n11 minus.n2 0.189894
R282 minus.n11 minus.n10 0.189894
R283 minus.n10 minus.n4 0.189894
R284 minus.n35 minus.n29 0.189894
R285 minus.n36 minus.n35 0.189894
R286 minus.n36 minus.n27 0.189894
R287 minus.n42 minus.n27 0.189894
R288 minus.n43 minus.n42 0.189894
R289 minus.n43 minus.n25 0.189894
R290 minus.n49 minus.n25 0.189894
R291 minus minus.n50 0.188
R292 drain_right.n10 drain_right.n8 60.2753
R293 drain_right.n6 drain_right.n4 60.2753
R294 drain_right.n2 drain_right.n0 60.2753
R295 drain_right.n10 drain_right.n9 59.8185
R296 drain_right.n12 drain_right.n11 59.8185
R297 drain_right.n14 drain_right.n13 59.8185
R298 drain_right.n16 drain_right.n15 59.8185
R299 drain_right.n7 drain_right.n3 59.8184
R300 drain_right.n6 drain_right.n5 59.8184
R301 drain_right.n2 drain_right.n1 59.8184
R302 drain_right drain_right.n7 36.5296
R303 drain_right drain_right.n16 6.11011
R304 drain_right.n3 drain_right.t2 0.9905
R305 drain_right.n3 drain_right.t8 0.9905
R306 drain_right.n4 drain_right.t7 0.9905
R307 drain_right.n4 drain_right.t13 0.9905
R308 drain_right.n5 drain_right.t5 0.9905
R309 drain_right.n5 drain_right.t9 0.9905
R310 drain_right.n1 drain_right.t17 0.9905
R311 drain_right.n1 drain_right.t11 0.9905
R312 drain_right.n0 drain_right.t15 0.9905
R313 drain_right.n0 drain_right.t10 0.9905
R314 drain_right.n8 drain_right.t14 0.9905
R315 drain_right.n8 drain_right.t4 0.9905
R316 drain_right.n9 drain_right.t1 0.9905
R317 drain_right.n9 drain_right.t19 0.9905
R318 drain_right.n11 drain_right.t16 0.9905
R319 drain_right.n11 drain_right.t3 0.9905
R320 drain_right.n13 drain_right.t0 0.9905
R321 drain_right.n13 drain_right.t18 0.9905
R322 drain_right.n15 drain_right.t12 0.9905
R323 drain_right.n15 drain_right.t6 0.9905
R324 drain_right.n16 drain_right.n14 0.457397
R325 drain_right.n14 drain_right.n12 0.457397
R326 drain_right.n12 drain_right.n10 0.457397
R327 drain_right.n7 drain_right.n6 0.402051
R328 drain_right.n7 drain_right.n2 0.402051
C0 minus plus 6.98315f
C1 source drain_right 73.2134f
C2 source minus 7.78142f
C3 minus drain_right 8.4922f
C4 drain_left plus 8.67526f
C5 drain_left source 73.2134f
C6 drain_left drain_right 0.982035f
C7 source plus 7.79546f
C8 drain_left minus 0.171252f
C9 drain_right plus 0.337271f
C10 drain_right a_n1882_n4888# 8.98437f
C11 drain_left a_n1882_n4888# 9.28558f
C12 source a_n1882_n4888# 12.844003f
C13 minus a_n1882_n4888# 7.850942f
C14 plus a_n1882_n4888# 10.495729f
C15 drain_right.t15 a_n1882_n4888# 0.621598f
C16 drain_right.t10 a_n1882_n4888# 0.621598f
C17 drain_right.n0 a_n1882_n4888# 5.6863f
C18 drain_right.t17 a_n1882_n4888# 0.621598f
C19 drain_right.t11 a_n1882_n4888# 0.621598f
C20 drain_right.n1 a_n1882_n4888# 5.68279f
C21 drain_right.n2 a_n1882_n4888# 0.902976f
C22 drain_right.t2 a_n1882_n4888# 0.621598f
C23 drain_right.t8 a_n1882_n4888# 0.621598f
C24 drain_right.n3 a_n1882_n4888# 5.68279f
C25 drain_right.t7 a_n1882_n4888# 0.621598f
C26 drain_right.t13 a_n1882_n4888# 0.621598f
C27 drain_right.n4 a_n1882_n4888# 5.6863f
C28 drain_right.t5 a_n1882_n4888# 0.621598f
C29 drain_right.t9 a_n1882_n4888# 0.621598f
C30 drain_right.n5 a_n1882_n4888# 5.68279f
C31 drain_right.n6 a_n1882_n4888# 0.902976f
C32 drain_right.n7 a_n1882_n4888# 3.01744f
C33 drain_right.t14 a_n1882_n4888# 0.621598f
C34 drain_right.t4 a_n1882_n4888# 0.621598f
C35 drain_right.n8 a_n1882_n4888# 5.68629f
C36 drain_right.t1 a_n1882_n4888# 0.621598f
C37 drain_right.t19 a_n1882_n4888# 0.621598f
C38 drain_right.n9 a_n1882_n4888# 5.68278f
C39 drain_right.n10 a_n1882_n4888# 0.907736f
C40 drain_right.t16 a_n1882_n4888# 0.621598f
C41 drain_right.t3 a_n1882_n4888# 0.621598f
C42 drain_right.n11 a_n1882_n4888# 5.68278f
C43 drain_right.n12 a_n1882_n4888# 0.447704f
C44 drain_right.t0 a_n1882_n4888# 0.621598f
C45 drain_right.t18 a_n1882_n4888# 0.621598f
C46 drain_right.n13 a_n1882_n4888# 5.68278f
C47 drain_right.n14 a_n1882_n4888# 0.447704f
C48 drain_right.t12 a_n1882_n4888# 0.621598f
C49 drain_right.t6 a_n1882_n4888# 0.621598f
C50 drain_right.n15 a_n1882_n4888# 5.68278f
C51 drain_right.n16 a_n1882_n4888# 0.769584f
C52 minus.n0 a_n1882_n4888# 0.053027f
C53 minus.t7 a_n1882_n4888# 0.602331f
C54 minus.t13 a_n1882_n4888# 0.597397f
C55 minus.t19 a_n1882_n4888# 0.597397f
C56 minus.t1 a_n1882_n4888# 0.597397f
C57 minus.n1 a_n1882_n4888# 0.227367f
C58 minus.n2 a_n1882_n4888# 0.053027f
C59 minus.t3 a_n1882_n4888# 0.597397f
C60 minus.t16 a_n1882_n4888# 0.597397f
C61 minus.t18 a_n1882_n4888# 0.597397f
C62 minus.n3 a_n1882_n4888# 0.227367f
C63 minus.n4 a_n1882_n4888# 0.121339f
C64 minus.t0 a_n1882_n4888# 0.597397f
C65 minus.t5 a_n1882_n4888# 0.597397f
C66 minus.t15 a_n1882_n4888# 0.602331f
C67 minus.n5 a_n1882_n4888# 0.243864f
C68 minus.n6 a_n1882_n4888# 0.227367f
C69 minus.n7 a_n1882_n4888# 0.018572f
C70 minus.n8 a_n1882_n4888# 0.227367f
C71 minus.n9 a_n1882_n4888# 0.018572f
C72 minus.n10 a_n1882_n4888# 0.053027f
C73 minus.n11 a_n1882_n4888# 0.053027f
C74 minus.n12 a_n1882_n4888# 0.018572f
C75 minus.n13 a_n1882_n4888# 0.227367f
C76 minus.n14 a_n1882_n4888# 0.018572f
C77 minus.n15 a_n1882_n4888# 0.227367f
C78 minus.n16 a_n1882_n4888# 0.018572f
C79 minus.n17 a_n1882_n4888# 0.053027f
C80 minus.n18 a_n1882_n4888# 0.053027f
C81 minus.n19 a_n1882_n4888# 0.018572f
C82 minus.n20 a_n1882_n4888# 0.227367f
C83 minus.n21 a_n1882_n4888# 0.018572f
C84 minus.n22 a_n1882_n4888# 0.227367f
C85 minus.n23 a_n1882_n4888# 0.243784f
C86 minus.n24 a_n1882_n4888# 2.37135f
C87 minus.n25 a_n1882_n4888# 0.053027f
C88 minus.t12 a_n1882_n4888# 0.597397f
C89 minus.t10 a_n1882_n4888# 0.597397f
C90 minus.t14 a_n1882_n4888# 0.597397f
C91 minus.n26 a_n1882_n4888# 0.227367f
C92 minus.n27 a_n1882_n4888# 0.053027f
C93 minus.t11 a_n1882_n4888# 0.597397f
C94 minus.t17 a_n1882_n4888# 0.597397f
C95 minus.t8 a_n1882_n4888# 0.597397f
C96 minus.n28 a_n1882_n4888# 0.227367f
C97 minus.n29 a_n1882_n4888# 0.121339f
C98 minus.t2 a_n1882_n4888# 0.597397f
C99 minus.t9 a_n1882_n4888# 0.597397f
C100 minus.t4 a_n1882_n4888# 0.602331f
C101 minus.n30 a_n1882_n4888# 0.243864f
C102 minus.n31 a_n1882_n4888# 0.227367f
C103 minus.n32 a_n1882_n4888# 0.018572f
C104 minus.n33 a_n1882_n4888# 0.227367f
C105 minus.n34 a_n1882_n4888# 0.018572f
C106 minus.n35 a_n1882_n4888# 0.053027f
C107 minus.n36 a_n1882_n4888# 0.053027f
C108 minus.n37 a_n1882_n4888# 0.018572f
C109 minus.n38 a_n1882_n4888# 0.227367f
C110 minus.n39 a_n1882_n4888# 0.018572f
C111 minus.n40 a_n1882_n4888# 0.227367f
C112 minus.n41 a_n1882_n4888# 0.018572f
C113 minus.n42 a_n1882_n4888# 0.053027f
C114 minus.n43 a_n1882_n4888# 0.053027f
C115 minus.n44 a_n1882_n4888# 0.018572f
C116 minus.n45 a_n1882_n4888# 0.227367f
C117 minus.n46 a_n1882_n4888# 0.018572f
C118 minus.n47 a_n1882_n4888# 0.227367f
C119 minus.t6 a_n1882_n4888# 0.602331f
C120 minus.n48 a_n1882_n4888# 0.243784f
C121 minus.n49 a_n1882_n4888# 0.343896f
C122 minus.n50 a_n1882_n4888# 2.83009f
C123 drain_left.t11 a_n1882_n4888# 0.621949f
C124 drain_left.t10 a_n1882_n4888# 0.621949f
C125 drain_left.n0 a_n1882_n4888# 5.6895f
C126 drain_left.t6 a_n1882_n4888# 0.621949f
C127 drain_left.t3 a_n1882_n4888# 0.621949f
C128 drain_left.n1 a_n1882_n4888# 5.68599f
C129 drain_left.n2 a_n1882_n4888# 0.903485f
C130 drain_left.t4 a_n1882_n4888# 0.621949f
C131 drain_left.t0 a_n1882_n4888# 0.621949f
C132 drain_left.n3 a_n1882_n4888# 5.68599f
C133 drain_left.t17 a_n1882_n4888# 0.621949f
C134 drain_left.t19 a_n1882_n4888# 0.621949f
C135 drain_left.n4 a_n1882_n4888# 5.6895f
C136 drain_left.t5 a_n1882_n4888# 0.621949f
C137 drain_left.t18 a_n1882_n4888# 0.621949f
C138 drain_left.n5 a_n1882_n4888# 5.68599f
C139 drain_left.n6 a_n1882_n4888# 0.903485f
C140 drain_left.n7 a_n1882_n4888# 3.10099f
C141 drain_left.t12 a_n1882_n4888# 0.621949f
C142 drain_left.t15 a_n1882_n4888# 0.621949f
C143 drain_left.n8 a_n1882_n4888# 5.6895f
C144 drain_left.t1 a_n1882_n4888# 0.621949f
C145 drain_left.t7 a_n1882_n4888# 0.621949f
C146 drain_left.n9 a_n1882_n4888# 5.68598f
C147 drain_left.n10 a_n1882_n4888# 0.908247f
C148 drain_left.t8 a_n1882_n4888# 0.621949f
C149 drain_left.t13 a_n1882_n4888# 0.621949f
C150 drain_left.n11 a_n1882_n4888# 5.68598f
C151 drain_left.n12 a_n1882_n4888# 0.447956f
C152 drain_left.t16 a_n1882_n4888# 0.621949f
C153 drain_left.t2 a_n1882_n4888# 0.621949f
C154 drain_left.n13 a_n1882_n4888# 5.68598f
C155 drain_left.n14 a_n1882_n4888# 0.447956f
C156 drain_left.t9 a_n1882_n4888# 0.621949f
C157 drain_left.t14 a_n1882_n4888# 0.621949f
C158 drain_left.n15 a_n1882_n4888# 5.68598f
C159 drain_left.n16 a_n1882_n4888# 0.770018f
C160 source.t27 a_n1882_n4888# 6.00904f
C161 source.n0 a_n1882_n4888# 2.54128f
C162 source.t24 a_n1882_n4888# 0.5258f
C163 source.t33 a_n1882_n4888# 0.5258f
C164 source.n1 a_n1882_n4888# 4.70088f
C165 source.n2 a_n1882_n4888# 0.439583f
C166 source.t22 a_n1882_n4888# 0.5258f
C167 source.t31 a_n1882_n4888# 0.5258f
C168 source.n3 a_n1882_n4888# 4.70088f
C169 source.n4 a_n1882_n4888# 0.439583f
C170 source.t29 a_n1882_n4888# 0.5258f
C171 source.t26 a_n1882_n4888# 0.5258f
C172 source.n5 a_n1882_n4888# 4.70088f
C173 source.n6 a_n1882_n4888# 0.439583f
C174 source.t23 a_n1882_n4888# 0.5258f
C175 source.t18 a_n1882_n4888# 0.5258f
C176 source.n7 a_n1882_n4888# 4.70088f
C177 source.n8 a_n1882_n4888# 0.439583f
C178 source.t30 a_n1882_n4888# 6.00906f
C179 source.n9 a_n1882_n4888# 0.566791f
C180 source.t6 a_n1882_n4888# 6.00906f
C181 source.n10 a_n1882_n4888# 0.566791f
C182 source.t7 a_n1882_n4888# 0.5258f
C183 source.t13 a_n1882_n4888# 0.5258f
C184 source.n11 a_n1882_n4888# 4.70088f
C185 source.n12 a_n1882_n4888# 0.439583f
C186 source.t38 a_n1882_n4888# 0.5258f
C187 source.t3 a_n1882_n4888# 0.5258f
C188 source.n13 a_n1882_n4888# 4.70088f
C189 source.n14 a_n1882_n4888# 0.439583f
C190 source.t10 a_n1882_n4888# 0.5258f
C191 source.t16 a_n1882_n4888# 0.5258f
C192 source.n15 a_n1882_n4888# 4.70088f
C193 source.n16 a_n1882_n4888# 0.439583f
C194 source.t15 a_n1882_n4888# 0.5258f
C195 source.t0 a_n1882_n4888# 0.5258f
C196 source.n17 a_n1882_n4888# 4.70088f
C197 source.n18 a_n1882_n4888# 0.439583f
C198 source.t17 a_n1882_n4888# 6.00906f
C199 source.n19 a_n1882_n4888# 3.12693f
C200 source.t21 a_n1882_n4888# 6.00902f
C201 source.n20 a_n1882_n4888# 3.12696f
C202 source.t28 a_n1882_n4888# 0.5258f
C203 source.t20 a_n1882_n4888# 0.5258f
C204 source.n21 a_n1882_n4888# 4.70089f
C205 source.n22 a_n1882_n4888# 0.439574f
C206 source.t37 a_n1882_n4888# 0.5258f
C207 source.t35 a_n1882_n4888# 0.5258f
C208 source.n23 a_n1882_n4888# 4.70089f
C209 source.n24 a_n1882_n4888# 0.439574f
C210 source.t25 a_n1882_n4888# 0.5258f
C211 source.t19 a_n1882_n4888# 0.5258f
C212 source.n25 a_n1882_n4888# 4.70089f
C213 source.n26 a_n1882_n4888# 0.439574f
C214 source.t36 a_n1882_n4888# 0.5258f
C215 source.t32 a_n1882_n4888# 0.5258f
C216 source.n27 a_n1882_n4888# 4.70089f
C217 source.n28 a_n1882_n4888# 0.439574f
C218 source.t34 a_n1882_n4888# 6.00902f
C219 source.n29 a_n1882_n4888# 0.566824f
C220 source.t9 a_n1882_n4888# 6.00902f
C221 source.n30 a_n1882_n4888# 0.566824f
C222 source.t5 a_n1882_n4888# 0.5258f
C223 source.t12 a_n1882_n4888# 0.5258f
C224 source.n31 a_n1882_n4888# 4.70089f
C225 source.n32 a_n1882_n4888# 0.439574f
C226 source.t2 a_n1882_n4888# 0.5258f
C227 source.t39 a_n1882_n4888# 0.5258f
C228 source.n33 a_n1882_n4888# 4.70089f
C229 source.n34 a_n1882_n4888# 0.439574f
C230 source.t4 a_n1882_n4888# 0.5258f
C231 source.t8 a_n1882_n4888# 0.5258f
C232 source.n35 a_n1882_n4888# 4.70089f
C233 source.n36 a_n1882_n4888# 0.439574f
C234 source.t1 a_n1882_n4888# 0.5258f
C235 source.t11 a_n1882_n4888# 0.5258f
C236 source.n37 a_n1882_n4888# 4.70089f
C237 source.n38 a_n1882_n4888# 0.439574f
C238 source.t14 a_n1882_n4888# 6.00902f
C239 source.n39 a_n1882_n4888# 0.747218f
C240 source.n40 a_n1882_n4888# 2.98907f
C241 plus.n0 a_n1882_n4888# 0.053729f
C242 plus.t10 a_n1882_n4888# 0.60531f
C243 plus.t17 a_n1882_n4888# 0.60531f
C244 plus.t3 a_n1882_n4888# 0.60531f
C245 plus.n1 a_n1882_n4888# 0.230379f
C246 plus.n2 a_n1882_n4888# 0.053729f
C247 plus.t6 a_n1882_n4888# 0.60531f
C248 plus.t11 a_n1882_n4888# 0.60531f
C249 plus.t12 a_n1882_n4888# 0.60531f
C250 plus.n3 a_n1882_n4888# 0.230379f
C251 plus.n4 a_n1882_n4888# 0.122947f
C252 plus.t18 a_n1882_n4888# 0.60531f
C253 plus.t4 a_n1882_n4888# 0.60531f
C254 plus.t7 a_n1882_n4888# 0.61031f
C255 plus.n5 a_n1882_n4888# 0.247094f
C256 plus.n6 a_n1882_n4888# 0.230379f
C257 plus.n7 a_n1882_n4888# 0.018818f
C258 plus.n8 a_n1882_n4888# 0.230379f
C259 plus.n9 a_n1882_n4888# 0.018818f
C260 plus.n10 a_n1882_n4888# 0.053729f
C261 plus.n11 a_n1882_n4888# 0.053729f
C262 plus.n12 a_n1882_n4888# 0.018818f
C263 plus.n13 a_n1882_n4888# 0.230379f
C264 plus.n14 a_n1882_n4888# 0.018818f
C265 plus.n15 a_n1882_n4888# 0.230379f
C266 plus.n16 a_n1882_n4888# 0.018818f
C267 plus.n17 a_n1882_n4888# 0.053729f
C268 plus.n18 a_n1882_n4888# 0.053729f
C269 plus.n19 a_n1882_n4888# 0.018818f
C270 plus.n20 a_n1882_n4888# 0.230379f
C271 plus.n21 a_n1882_n4888# 0.018818f
C272 plus.n22 a_n1882_n4888# 0.230379f
C273 plus.t5 a_n1882_n4888# 0.61031f
C274 plus.n23 a_n1882_n4888# 0.247013f
C275 plus.n24 a_n1882_n4888# 0.813095f
C276 plus.n25 a_n1882_n4888# 0.053729f
C277 plus.t8 a_n1882_n4888# 0.61031f
C278 plus.t9 a_n1882_n4888# 0.60531f
C279 plus.t13 a_n1882_n4888# 0.60531f
C280 plus.t16 a_n1882_n4888# 0.60531f
C281 plus.n26 a_n1882_n4888# 0.230379f
C282 plus.n27 a_n1882_n4888# 0.053729f
C283 plus.t15 a_n1882_n4888# 0.60531f
C284 plus.t19 a_n1882_n4888# 0.60531f
C285 plus.t14 a_n1882_n4888# 0.60531f
C286 plus.n28 a_n1882_n4888# 0.230379f
C287 plus.n29 a_n1882_n4888# 0.122947f
C288 plus.t1 a_n1882_n4888# 0.60531f
C289 plus.t2 a_n1882_n4888# 0.60531f
C290 plus.t0 a_n1882_n4888# 0.61031f
C291 plus.n30 a_n1882_n4888# 0.247094f
C292 plus.n31 a_n1882_n4888# 0.230379f
C293 plus.n32 a_n1882_n4888# 0.018818f
C294 plus.n33 a_n1882_n4888# 0.230379f
C295 plus.n34 a_n1882_n4888# 0.018818f
C296 plus.n35 a_n1882_n4888# 0.053729f
C297 plus.n36 a_n1882_n4888# 0.053729f
C298 plus.n37 a_n1882_n4888# 0.018818f
C299 plus.n38 a_n1882_n4888# 0.230379f
C300 plus.n39 a_n1882_n4888# 0.018818f
C301 plus.n40 a_n1882_n4888# 0.230379f
C302 plus.n41 a_n1882_n4888# 0.018818f
C303 plus.n42 a_n1882_n4888# 0.053729f
C304 plus.n43 a_n1882_n4888# 0.053729f
C305 plus.n44 a_n1882_n4888# 0.018818f
C306 plus.n45 a_n1882_n4888# 0.230379f
C307 plus.n46 a_n1882_n4888# 0.018818f
C308 plus.n47 a_n1882_n4888# 0.230379f
C309 plus.n48 a_n1882_n4888# 0.247013f
C310 plus.n49 a_n1882_n4888# 1.90091f
.ends

