* NGSPICE file created from diffpair238.ext - technology: sky130A

.subckt diffpair238 minus drain_right drain_left source plus
X0 source.t37 minus.t0 drain_right.t19 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X1 source.t36 minus.t1 drain_right.t13 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X2 a_n3202_n1488# a_n3202_n1488# a_n3202_n1488# a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.8
X3 drain_left.t19 plus.t0 source.t2 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X4 drain_left.t18 plus.t1 source.t7 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X5 drain_left.t17 plus.t2 source.t14 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X6 a_n3202_n1488# a_n3202_n1488# a_n3202_n1488# a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X7 source.t35 minus.t2 drain_right.t2 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X8 source.t34 minus.t3 drain_right.t3 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X9 source.t33 minus.t4 drain_right.t9 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X10 drain_left.t16 plus.t3 source.t1 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X11 drain_left.t15 plus.t4 source.t8 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X12 source.t32 minus.t5 drain_right.t6 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X13 source.t3 plus.t5 drain_left.t14 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X14 drain_right.t0 minus.t6 source.t31 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X15 drain_right.t7 minus.t7 source.t30 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X16 drain_left.t13 plus.t6 source.t9 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X17 source.t29 minus.t8 drain_right.t4 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X18 drain_right.t8 minus.t9 source.t28 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X19 drain_right.t10 minus.t10 source.t27 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X20 a_n3202_n1488# a_n3202_n1488# a_n3202_n1488# a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X21 drain_right.t5 minus.t11 source.t26 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X22 a_n3202_n1488# a_n3202_n1488# a_n3202_n1488# a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.8
X23 source.t17 plus.t7 drain_left.t12 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X24 source.t25 minus.t12 drain_right.t1 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X25 drain_right.t12 minus.t13 source.t24 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X26 drain_right.t11 minus.t14 source.t23 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X27 source.t13 plus.t8 drain_left.t11 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X28 drain_left.t10 plus.t9 source.t5 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X29 source.t22 minus.t15 drain_right.t14 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X30 drain_right.t15 minus.t16 source.t21 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X31 source.t0 plus.t10 drain_left.t9 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X32 source.t11 plus.t11 drain_left.t8 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X33 drain_right.t16 minus.t17 source.t20 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X34 source.t6 plus.t12 drain_left.t7 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X35 drain_left.t6 plus.t13 source.t4 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X36 drain_left.t5 plus.t14 source.t12 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X37 source.t19 minus.t18 drain_right.t17 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X38 drain_right.t18 minus.t19 source.t18 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.8
X39 source.t38 plus.t15 drain_left.t4 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X40 source.t10 plus.t16 drain_left.t3 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
X41 source.t16 plus.t17 drain_left.t2 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X42 drain_left.t1 plus.t18 source.t15 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.8
X43 source.t39 plus.t19 drain_left.t0 a_n3202_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.8
R0 minus.n29 minus.n28 161.3
R1 minus.n27 minus.n0 161.3
R2 minus.n26 minus.n25 161.3
R3 minus.n24 minus.n1 161.3
R4 minus.n20 minus.n19 161.3
R5 minus.n18 minus.n3 161.3
R6 minus.n17 minus.n16 161.3
R7 minus.n15 minus.n4 161.3
R8 minus.n14 minus.n13 161.3
R9 minus.n9 minus.n6 161.3
R10 minus.n59 minus.n58 161.3
R11 minus.n57 minus.n30 161.3
R12 minus.n56 minus.n55 161.3
R13 minus.n54 minus.n31 161.3
R14 minus.n50 minus.n49 161.3
R15 minus.n48 minus.n33 161.3
R16 minus.n47 minus.n46 161.3
R17 minus.n45 minus.n34 161.3
R18 minus.n44 minus.n43 161.3
R19 minus.n39 minus.n36 161.3
R20 minus.n7 minus.t11 161.269
R21 minus.n37 minus.t3 161.269
R22 minus.n8 minus.t8 139.48
R23 minus.n10 minus.t6 139.48
R24 minus.n5 minus.t15 139.48
R25 minus.n15 minus.t17 139.48
R26 minus.n3 minus.t12 139.48
R27 minus.n21 minus.t10 139.48
R28 minus.n22 minus.t18 139.48
R29 minus.n26 minus.t16 139.48
R30 minus.n28 minus.t5 139.48
R31 minus.n38 minus.t7 139.48
R32 minus.n40 minus.t4 139.48
R33 minus.n35 minus.t9 139.48
R34 minus.n45 minus.t0 139.48
R35 minus.n33 minus.t14 139.48
R36 minus.n51 minus.t1 139.48
R37 minus.n52 minus.t13 139.48
R38 minus.n56 minus.t2 139.48
R39 minus.n58 minus.t19 139.48
R40 minus.n23 minus.n22 80.6037
R41 minus.n21 minus.n2 80.6037
R42 minus.n12 minus.n5 80.6037
R43 minus.n11 minus.n10 80.6037
R44 minus.n53 minus.n52 80.6037
R45 minus.n51 minus.n32 80.6037
R46 minus.n42 minus.n35 80.6037
R47 minus.n41 minus.n40 80.6037
R48 minus.n10 minus.n5 48.2005
R49 minus.n22 minus.n21 48.2005
R50 minus.n40 minus.n35 48.2005
R51 minus.n52 minus.n51 48.2005
R52 minus.n7 minus.n6 44.8565
R53 minus.n37 minus.n36 44.8565
R54 minus.n14 minus.n5 43.0884
R55 minus.n21 minus.n20 43.0884
R56 minus.n44 minus.n35 43.0884
R57 minus.n51 minus.n50 43.0884
R58 minus.n10 minus.n9 40.1672
R59 minus.n22 minus.n1 40.1672
R60 minus.n40 minus.n39 40.1672
R61 minus.n52 minus.n31 40.1672
R62 minus.n60 minus.n29 34.6369
R63 minus.n28 minus.n27 27.0217
R64 minus.n58 minus.n57 27.0217
R65 minus.n16 minus.n3 24.1005
R66 minus.n16 minus.n15 24.1005
R67 minus.n46 minus.n45 24.1005
R68 minus.n46 minus.n33 24.1005
R69 minus.n27 minus.n26 21.1793
R70 minus.n57 minus.n56 21.1793
R71 minus.n8 minus.n7 20.1275
R72 minus.n38 minus.n37 20.1275
R73 minus.n9 minus.n8 8.03383
R74 minus.n26 minus.n1 8.03383
R75 minus.n39 minus.n38 8.03383
R76 minus.n56 minus.n31 8.03383
R77 minus.n60 minus.n59 6.70505
R78 minus.n15 minus.n14 5.11262
R79 minus.n20 minus.n3 5.11262
R80 minus.n45 minus.n44 5.11262
R81 minus.n50 minus.n33 5.11262
R82 minus.n23 minus.n2 0.380177
R83 minus.n12 minus.n11 0.380177
R84 minus.n42 minus.n41 0.380177
R85 minus.n53 minus.n32 0.380177
R86 minus.n24 minus.n23 0.285035
R87 minus.n19 minus.n2 0.285035
R88 minus.n13 minus.n12 0.285035
R89 minus.n11 minus.n6 0.285035
R90 minus.n41 minus.n36 0.285035
R91 minus.n43 minus.n42 0.285035
R92 minus.n49 minus.n32 0.285035
R93 minus.n54 minus.n53 0.285035
R94 minus.n29 minus.n0 0.189894
R95 minus.n25 minus.n0 0.189894
R96 minus.n25 minus.n24 0.189894
R97 minus.n19 minus.n18 0.189894
R98 minus.n18 minus.n17 0.189894
R99 minus.n17 minus.n4 0.189894
R100 minus.n13 minus.n4 0.189894
R101 minus.n43 minus.n34 0.189894
R102 minus.n47 minus.n34 0.189894
R103 minus.n48 minus.n47 0.189894
R104 minus.n49 minus.n48 0.189894
R105 minus.n55 minus.n54 0.189894
R106 minus.n55 minus.n30 0.189894
R107 minus.n59 minus.n30 0.189894
R108 minus minus.n60 0.188
R109 drain_right.n10 drain_right.n8 80.7472
R110 drain_right.n6 drain_right.n4 80.7471
R111 drain_right.n2 drain_right.n0 80.7471
R112 drain_right.n10 drain_right.n9 79.7731
R113 drain_right.n12 drain_right.n11 79.7731
R114 drain_right.n14 drain_right.n13 79.7731
R115 drain_right.n16 drain_right.n15 79.7731
R116 drain_right.n7 drain_right.n3 79.773
R117 drain_right.n6 drain_right.n5 79.773
R118 drain_right.n2 drain_right.n1 79.773
R119 drain_right drain_right.n7 27.7888
R120 drain_right drain_right.n16 6.62735
R121 drain_right.n3 drain_right.t19 6.6005
R122 drain_right.n3 drain_right.t11 6.6005
R123 drain_right.n4 drain_right.t2 6.6005
R124 drain_right.n4 drain_right.t18 6.6005
R125 drain_right.n5 drain_right.t13 6.6005
R126 drain_right.n5 drain_right.t12 6.6005
R127 drain_right.n1 drain_right.t9 6.6005
R128 drain_right.n1 drain_right.t8 6.6005
R129 drain_right.n0 drain_right.t3 6.6005
R130 drain_right.n0 drain_right.t7 6.6005
R131 drain_right.n8 drain_right.t4 6.6005
R132 drain_right.n8 drain_right.t5 6.6005
R133 drain_right.n9 drain_right.t14 6.6005
R134 drain_right.n9 drain_right.t0 6.6005
R135 drain_right.n11 drain_right.t1 6.6005
R136 drain_right.n11 drain_right.t16 6.6005
R137 drain_right.n13 drain_right.t17 6.6005
R138 drain_right.n13 drain_right.t10 6.6005
R139 drain_right.n15 drain_right.t6 6.6005
R140 drain_right.n15 drain_right.t15 6.6005
R141 drain_right.n16 drain_right.n14 0.974638
R142 drain_right.n14 drain_right.n12 0.974638
R143 drain_right.n12 drain_right.n10 0.974638
R144 drain_right.n7 drain_right.n6 0.919292
R145 drain_right.n7 drain_right.n2 0.919292
R146 source.n0 source.t9 69.6943
R147 source.n9 source.t39 69.6943
R148 source.n10 source.t26 69.6943
R149 source.n19 source.t32 69.6943
R150 source.n39 source.t18 69.6942
R151 source.n30 source.t34 69.6942
R152 source.n29 source.t1 69.6942
R153 source.n20 source.t10 69.6942
R154 source.n2 source.n1 63.0943
R155 source.n4 source.n3 63.0943
R156 source.n6 source.n5 63.0943
R157 source.n8 source.n7 63.0943
R158 source.n12 source.n11 63.0943
R159 source.n14 source.n13 63.0943
R160 source.n16 source.n15 63.0943
R161 source.n18 source.n17 63.0943
R162 source.n38 source.n37 63.0942
R163 source.n36 source.n35 63.0942
R164 source.n34 source.n33 63.0942
R165 source.n32 source.n31 63.0942
R166 source.n28 source.n27 63.0942
R167 source.n26 source.n25 63.0942
R168 source.n24 source.n23 63.0942
R169 source.n22 source.n21 63.0942
R170 source.n20 source.n19 15.4437
R171 source.n40 source.n0 9.69368
R172 source.n37 source.t24 6.6005
R173 source.n37 source.t35 6.6005
R174 source.n35 source.t23 6.6005
R175 source.n35 source.t36 6.6005
R176 source.n33 source.t28 6.6005
R177 source.n33 source.t37 6.6005
R178 source.n31 source.t30 6.6005
R179 source.n31 source.t33 6.6005
R180 source.n27 source.t8 6.6005
R181 source.n27 source.t13 6.6005
R182 source.n25 source.t2 6.6005
R183 source.n25 source.t0 6.6005
R184 source.n23 source.t7 6.6005
R185 source.n23 source.t11 6.6005
R186 source.n21 source.t14 6.6005
R187 source.n21 source.t3 6.6005
R188 source.n1 source.t5 6.6005
R189 source.n1 source.t17 6.6005
R190 source.n3 source.t4 6.6005
R191 source.n3 source.t6 6.6005
R192 source.n5 source.t12 6.6005
R193 source.n5 source.t16 6.6005
R194 source.n7 source.t15 6.6005
R195 source.n7 source.t38 6.6005
R196 source.n11 source.t31 6.6005
R197 source.n11 source.t29 6.6005
R198 source.n13 source.t20 6.6005
R199 source.n13 source.t22 6.6005
R200 source.n15 source.t27 6.6005
R201 source.n15 source.t25 6.6005
R202 source.n17 source.t21 6.6005
R203 source.n17 source.t19 6.6005
R204 source.n40 source.n39 5.7505
R205 source.n19 source.n18 0.974638
R206 source.n18 source.n16 0.974638
R207 source.n16 source.n14 0.974638
R208 source.n14 source.n12 0.974638
R209 source.n12 source.n10 0.974638
R210 source.n9 source.n8 0.974638
R211 source.n8 source.n6 0.974638
R212 source.n6 source.n4 0.974638
R213 source.n4 source.n2 0.974638
R214 source.n2 source.n0 0.974638
R215 source.n22 source.n20 0.974638
R216 source.n24 source.n22 0.974638
R217 source.n26 source.n24 0.974638
R218 source.n28 source.n26 0.974638
R219 source.n29 source.n28 0.974638
R220 source.n32 source.n30 0.974638
R221 source.n34 source.n32 0.974638
R222 source.n36 source.n34 0.974638
R223 source.n38 source.n36 0.974638
R224 source.n39 source.n38 0.974638
R225 source.n10 source.n9 0.470328
R226 source.n30 source.n29 0.470328
R227 source source.n40 0.188
R228 plus.n11 plus.n10 161.3
R229 plus.n15 plus.n14 161.3
R230 plus.n16 plus.n5 161.3
R231 plus.n18 plus.n17 161.3
R232 plus.n19 plus.n4 161.3
R233 plus.n20 plus.n3 161.3
R234 plus.n25 plus.n24 161.3
R235 plus.n26 plus.n1 161.3
R236 plus.n27 plus.n0 161.3
R237 plus.n29 plus.n28 161.3
R238 plus.n41 plus.n40 161.3
R239 plus.n45 plus.n44 161.3
R240 plus.n46 plus.n35 161.3
R241 plus.n48 plus.n47 161.3
R242 plus.n49 plus.n34 161.3
R243 plus.n50 plus.n33 161.3
R244 plus.n55 plus.n54 161.3
R245 plus.n56 plus.n31 161.3
R246 plus.n57 plus.n30 161.3
R247 plus.n59 plus.n58 161.3
R248 plus.n9 plus.t19 161.269
R249 plus.n39 plus.t3 161.269
R250 plus.n28 plus.t6 139.48
R251 plus.n26 plus.t7 139.48
R252 plus.n2 plus.t9 139.48
R253 plus.n21 plus.t12 139.48
R254 plus.n19 plus.t13 139.48
R255 plus.n5 plus.t17 139.48
R256 plus.n13 plus.t14 139.48
R257 plus.n12 plus.t15 139.48
R258 plus.n8 plus.t18 139.48
R259 plus.n58 plus.t16 139.48
R260 plus.n56 plus.t2 139.48
R261 plus.n32 plus.t5 139.48
R262 plus.n51 plus.t1 139.48
R263 plus.n49 plus.t11 139.48
R264 plus.n35 plus.t0 139.48
R265 plus.n43 plus.t10 139.48
R266 plus.n42 plus.t4 139.48
R267 plus.n38 plus.t8 139.48
R268 plus.n12 plus.n7 80.6037
R269 plus.n13 plus.n6 80.6037
R270 plus.n22 plus.n21 80.6037
R271 plus.n23 plus.n2 80.6037
R272 plus.n42 plus.n37 80.6037
R273 plus.n43 plus.n36 80.6037
R274 plus.n52 plus.n51 80.6037
R275 plus.n53 plus.n32 80.6037
R276 plus.n21 plus.n2 48.2005
R277 plus.n13 plus.n12 48.2005
R278 plus.n51 plus.n32 48.2005
R279 plus.n43 plus.n42 48.2005
R280 plus.n40 plus.n39 44.8565
R281 plus.n10 plus.n9 44.8565
R282 plus.n21 plus.n20 43.0884
R283 plus.n14 plus.n13 43.0884
R284 plus.n51 plus.n50 43.0884
R285 plus.n44 plus.n43 43.0884
R286 plus.n25 plus.n2 40.1672
R287 plus.n12 plus.n11 40.1672
R288 plus.n55 plus.n32 40.1672
R289 plus.n42 plus.n41 40.1672
R290 plus plus.n59 31.9271
R291 plus.n28 plus.n27 27.0217
R292 plus.n58 plus.n57 27.0217
R293 plus.n18 plus.n5 24.1005
R294 plus.n19 plus.n18 24.1005
R295 plus.n49 plus.n48 24.1005
R296 plus.n48 plus.n35 24.1005
R297 plus.n27 plus.n26 21.1793
R298 plus.n57 plus.n56 21.1793
R299 plus.n39 plus.n38 20.1275
R300 plus.n9 plus.n8 20.1275
R301 plus plus.n29 8.93989
R302 plus.n26 plus.n25 8.03383
R303 plus.n11 plus.n8 8.03383
R304 plus.n56 plus.n55 8.03383
R305 plus.n41 plus.n38 8.03383
R306 plus.n20 plus.n19 5.11262
R307 plus.n14 plus.n5 5.11262
R308 plus.n50 plus.n49 5.11262
R309 plus.n44 plus.n35 5.11262
R310 plus.n7 plus.n6 0.380177
R311 plus.n23 plus.n22 0.380177
R312 plus.n53 plus.n52 0.380177
R313 plus.n37 plus.n36 0.380177
R314 plus.n10 plus.n7 0.285035
R315 plus.n15 plus.n6 0.285035
R316 plus.n22 plus.n3 0.285035
R317 plus.n24 plus.n23 0.285035
R318 plus.n54 plus.n53 0.285035
R319 plus.n52 plus.n33 0.285035
R320 plus.n45 plus.n36 0.285035
R321 plus.n40 plus.n37 0.285035
R322 plus.n16 plus.n15 0.189894
R323 plus.n17 plus.n16 0.189894
R324 plus.n17 plus.n4 0.189894
R325 plus.n4 plus.n3 0.189894
R326 plus.n24 plus.n1 0.189894
R327 plus.n1 plus.n0 0.189894
R328 plus.n29 plus.n0 0.189894
R329 plus.n59 plus.n30 0.189894
R330 plus.n31 plus.n30 0.189894
R331 plus.n54 plus.n31 0.189894
R332 plus.n34 plus.n33 0.189894
R333 plus.n47 plus.n34 0.189894
R334 plus.n47 plus.n46 0.189894
R335 plus.n46 plus.n45 0.189894
R336 drain_left.n10 drain_left.n8 80.7472
R337 drain_left.n6 drain_left.n4 80.7471
R338 drain_left.n2 drain_left.n0 80.7471
R339 drain_left.n16 drain_left.n15 79.7731
R340 drain_left.n14 drain_left.n13 79.7731
R341 drain_left.n12 drain_left.n11 79.7731
R342 drain_left.n10 drain_left.n9 79.7731
R343 drain_left.n7 drain_left.n3 79.773
R344 drain_left.n6 drain_left.n5 79.773
R345 drain_left.n2 drain_left.n1 79.773
R346 drain_left drain_left.n7 28.342
R347 drain_left drain_left.n16 6.62735
R348 drain_left.n3 drain_left.t8 6.6005
R349 drain_left.n3 drain_left.t19 6.6005
R350 drain_left.n4 drain_left.t11 6.6005
R351 drain_left.n4 drain_left.t16 6.6005
R352 drain_left.n5 drain_left.t9 6.6005
R353 drain_left.n5 drain_left.t15 6.6005
R354 drain_left.n1 drain_left.t14 6.6005
R355 drain_left.n1 drain_left.t18 6.6005
R356 drain_left.n0 drain_left.t3 6.6005
R357 drain_left.n0 drain_left.t17 6.6005
R358 drain_left.n15 drain_left.t12 6.6005
R359 drain_left.n15 drain_left.t13 6.6005
R360 drain_left.n13 drain_left.t7 6.6005
R361 drain_left.n13 drain_left.t10 6.6005
R362 drain_left.n11 drain_left.t2 6.6005
R363 drain_left.n11 drain_left.t6 6.6005
R364 drain_left.n9 drain_left.t4 6.6005
R365 drain_left.n9 drain_left.t5 6.6005
R366 drain_left.n8 drain_left.t0 6.6005
R367 drain_left.n8 drain_left.t1 6.6005
R368 drain_left.n12 drain_left.n10 0.974638
R369 drain_left.n14 drain_left.n12 0.974638
R370 drain_left.n16 drain_left.n14 0.974638
R371 drain_left.n7 drain_left.n6 0.919292
R372 drain_left.n7 drain_left.n2 0.919292
C0 drain_right minus 3.91605f
C1 drain_right source 8.869861f
C2 drain_right plus 0.483962f
C3 minus source 4.67712f
C4 minus plus 5.47845f
C5 plus source 4.69112f
C6 drain_right drain_left 1.7292f
C7 minus drain_left 0.179123f
C8 drain_left source 8.866981f
C9 plus drain_left 4.23637f
C10 drain_right a_n3202_n1488# 5.82042f
C11 drain_left a_n3202_n1488# 6.2797f
C12 source a_n3202_n1488# 4.184525f
C13 minus a_n3202_n1488# 12.155634f
C14 plus a_n3202_n1488# 13.560131f
C15 drain_left.t3 a_n3202_n1488# 0.06358f
C16 drain_left.t17 a_n3202_n1488# 0.06358f
C17 drain_left.n0 a_n3202_n1488# 0.463284f
C18 drain_left.t14 a_n3202_n1488# 0.06358f
C19 drain_left.t18 a_n3202_n1488# 0.06358f
C20 drain_left.n1 a_n3202_n1488# 0.458532f
C21 drain_left.n2 a_n3202_n1488# 0.768042f
C22 drain_left.t8 a_n3202_n1488# 0.06358f
C23 drain_left.t19 a_n3202_n1488# 0.06358f
C24 drain_left.n3 a_n3202_n1488# 0.458532f
C25 drain_left.t11 a_n3202_n1488# 0.06358f
C26 drain_left.t16 a_n3202_n1488# 0.06358f
C27 drain_left.n4 a_n3202_n1488# 0.463284f
C28 drain_left.t9 a_n3202_n1488# 0.06358f
C29 drain_left.t15 a_n3202_n1488# 0.06358f
C30 drain_left.n5 a_n3202_n1488# 0.458532f
C31 drain_left.n6 a_n3202_n1488# 0.768042f
C32 drain_left.n7 a_n3202_n1488# 1.50733f
C33 drain_left.t0 a_n3202_n1488# 0.06358f
C34 drain_left.t1 a_n3202_n1488# 0.06358f
C35 drain_left.n8 a_n3202_n1488# 0.463286f
C36 drain_left.t4 a_n3202_n1488# 0.06358f
C37 drain_left.t5 a_n3202_n1488# 0.06358f
C38 drain_left.n9 a_n3202_n1488# 0.458535f
C39 drain_left.n10 a_n3202_n1488# 0.772143f
C40 drain_left.t2 a_n3202_n1488# 0.06358f
C41 drain_left.t6 a_n3202_n1488# 0.06358f
C42 drain_left.n11 a_n3202_n1488# 0.458535f
C43 drain_left.n12 a_n3202_n1488# 0.383046f
C44 drain_left.t7 a_n3202_n1488# 0.06358f
C45 drain_left.t10 a_n3202_n1488# 0.06358f
C46 drain_left.n13 a_n3202_n1488# 0.458535f
C47 drain_left.n14 a_n3202_n1488# 0.383046f
C48 drain_left.t12 a_n3202_n1488# 0.06358f
C49 drain_left.t13 a_n3202_n1488# 0.06358f
C50 drain_left.n15 a_n3202_n1488# 0.458535f
C51 drain_left.n16 a_n3202_n1488# 0.623532f
C52 plus.n0 a_n3202_n1488# 0.041034f
C53 plus.t6 a_n3202_n1488# 0.295307f
C54 plus.t7 a_n3202_n1488# 0.295307f
C55 plus.n1 a_n3202_n1488# 0.041034f
C56 plus.t9 a_n3202_n1488# 0.295307f
C57 plus.n2 a_n3202_n1488# 0.179451f
C58 plus.n3 a_n3202_n1488# 0.054754f
C59 plus.t12 a_n3202_n1488# 0.295307f
C60 plus.t13 a_n3202_n1488# 0.295307f
C61 plus.n4 a_n3202_n1488# 0.041034f
C62 plus.t17 a_n3202_n1488# 0.295307f
C63 plus.n5 a_n3202_n1488# 0.168242f
C64 plus.n6 a_n3202_n1488# 0.068346f
C65 plus.t14 a_n3202_n1488# 0.295307f
C66 plus.t15 a_n3202_n1488# 0.295307f
C67 plus.n7 a_n3202_n1488# 0.068346f
C68 plus.t18 a_n3202_n1488# 0.295307f
C69 plus.n8 a_n3202_n1488# 0.171691f
C70 plus.t19 a_n3202_n1488# 0.318349f
C71 plus.n9 a_n3202_n1488# 0.151552f
C72 plus.n10 a_n3202_n1488# 0.188876f
C73 plus.n11 a_n3202_n1488# 0.009311f
C74 plus.n12 a_n3202_n1488# 0.179451f
C75 plus.n13 a_n3202_n1488# 0.179957f
C76 plus.n14 a_n3202_n1488# 0.009311f
C77 plus.n15 a_n3202_n1488# 0.054754f
C78 plus.n16 a_n3202_n1488# 0.041034f
C79 plus.n17 a_n3202_n1488# 0.041034f
C80 plus.n18 a_n3202_n1488# 0.009311f
C81 plus.n19 a_n3202_n1488# 0.168242f
C82 plus.n20 a_n3202_n1488# 0.009311f
C83 plus.n21 a_n3202_n1488# 0.179957f
C84 plus.n22 a_n3202_n1488# 0.068346f
C85 plus.n23 a_n3202_n1488# 0.068346f
C86 plus.n24 a_n3202_n1488# 0.054754f
C87 plus.n25 a_n3202_n1488# 0.009311f
C88 plus.n26 a_n3202_n1488# 0.168242f
C89 plus.n27 a_n3202_n1488# 0.009311f
C90 plus.n28 a_n3202_n1488# 0.167863f
C91 plus.n29 a_n3202_n1488# 0.327211f
C92 plus.n30 a_n3202_n1488# 0.041034f
C93 plus.t16 a_n3202_n1488# 0.295307f
C94 plus.n31 a_n3202_n1488# 0.041034f
C95 plus.t2 a_n3202_n1488# 0.295307f
C96 plus.t5 a_n3202_n1488# 0.295307f
C97 plus.n32 a_n3202_n1488# 0.179451f
C98 plus.n33 a_n3202_n1488# 0.054754f
C99 plus.t1 a_n3202_n1488# 0.295307f
C100 plus.n34 a_n3202_n1488# 0.041034f
C101 plus.t11 a_n3202_n1488# 0.295307f
C102 plus.t0 a_n3202_n1488# 0.295307f
C103 plus.n35 a_n3202_n1488# 0.168242f
C104 plus.n36 a_n3202_n1488# 0.068346f
C105 plus.t10 a_n3202_n1488# 0.295307f
C106 plus.n37 a_n3202_n1488# 0.068346f
C107 plus.t4 a_n3202_n1488# 0.295307f
C108 plus.t8 a_n3202_n1488# 0.295307f
C109 plus.n38 a_n3202_n1488# 0.171691f
C110 plus.t3 a_n3202_n1488# 0.318349f
C111 plus.n39 a_n3202_n1488# 0.151552f
C112 plus.n40 a_n3202_n1488# 0.188876f
C113 plus.n41 a_n3202_n1488# 0.009311f
C114 plus.n42 a_n3202_n1488# 0.179451f
C115 plus.n43 a_n3202_n1488# 0.179957f
C116 plus.n44 a_n3202_n1488# 0.009311f
C117 plus.n45 a_n3202_n1488# 0.054754f
C118 plus.n46 a_n3202_n1488# 0.041034f
C119 plus.n47 a_n3202_n1488# 0.041034f
C120 plus.n48 a_n3202_n1488# 0.009311f
C121 plus.n49 a_n3202_n1488# 0.168242f
C122 plus.n50 a_n3202_n1488# 0.009311f
C123 plus.n51 a_n3202_n1488# 0.179957f
C124 plus.n52 a_n3202_n1488# 0.068346f
C125 plus.n53 a_n3202_n1488# 0.068346f
C126 plus.n54 a_n3202_n1488# 0.054754f
C127 plus.n55 a_n3202_n1488# 0.009311f
C128 plus.n56 a_n3202_n1488# 0.168242f
C129 plus.n57 a_n3202_n1488# 0.009311f
C130 plus.n58 a_n3202_n1488# 0.167863f
C131 plus.n59 a_n3202_n1488# 1.27691f
C132 source.t9 a_n3202_n1488# 0.571448f
C133 source.n0 a_n3202_n1488# 0.850419f
C134 source.t5 a_n3202_n1488# 0.068817f
C135 source.t17 a_n3202_n1488# 0.068817f
C136 source.n1 a_n3202_n1488# 0.436342f
C137 source.n2 a_n3202_n1488# 0.435109f
C138 source.t4 a_n3202_n1488# 0.068817f
C139 source.t6 a_n3202_n1488# 0.068817f
C140 source.n3 a_n3202_n1488# 0.436342f
C141 source.n4 a_n3202_n1488# 0.435109f
C142 source.t12 a_n3202_n1488# 0.068817f
C143 source.t16 a_n3202_n1488# 0.068817f
C144 source.n5 a_n3202_n1488# 0.436342f
C145 source.n6 a_n3202_n1488# 0.435109f
C146 source.t15 a_n3202_n1488# 0.068817f
C147 source.t38 a_n3202_n1488# 0.068817f
C148 source.n7 a_n3202_n1488# 0.436342f
C149 source.n8 a_n3202_n1488# 0.435109f
C150 source.t39 a_n3202_n1488# 0.571448f
C151 source.n9 a_n3202_n1488# 0.440516f
C152 source.t26 a_n3202_n1488# 0.571448f
C153 source.n10 a_n3202_n1488# 0.440516f
C154 source.t31 a_n3202_n1488# 0.068817f
C155 source.t29 a_n3202_n1488# 0.068817f
C156 source.n11 a_n3202_n1488# 0.436342f
C157 source.n12 a_n3202_n1488# 0.435109f
C158 source.t20 a_n3202_n1488# 0.068817f
C159 source.t22 a_n3202_n1488# 0.068817f
C160 source.n13 a_n3202_n1488# 0.436342f
C161 source.n14 a_n3202_n1488# 0.435109f
C162 source.t27 a_n3202_n1488# 0.068817f
C163 source.t25 a_n3202_n1488# 0.068817f
C164 source.n15 a_n3202_n1488# 0.436342f
C165 source.n16 a_n3202_n1488# 0.435109f
C166 source.t21 a_n3202_n1488# 0.068817f
C167 source.t19 a_n3202_n1488# 0.068817f
C168 source.n17 a_n3202_n1488# 0.436342f
C169 source.n18 a_n3202_n1488# 0.435109f
C170 source.t32 a_n3202_n1488# 0.571448f
C171 source.n19 a_n3202_n1488# 1.16286f
C172 source.t10 a_n3202_n1488# 0.571445f
C173 source.n20 a_n3202_n1488# 1.16287f
C174 source.t14 a_n3202_n1488# 0.068817f
C175 source.t3 a_n3202_n1488# 0.068817f
C176 source.n21 a_n3202_n1488# 0.436339f
C177 source.n22 a_n3202_n1488# 0.435112f
C178 source.t7 a_n3202_n1488# 0.068817f
C179 source.t11 a_n3202_n1488# 0.068817f
C180 source.n23 a_n3202_n1488# 0.436339f
C181 source.n24 a_n3202_n1488# 0.435112f
C182 source.t2 a_n3202_n1488# 0.068817f
C183 source.t0 a_n3202_n1488# 0.068817f
C184 source.n25 a_n3202_n1488# 0.436339f
C185 source.n26 a_n3202_n1488# 0.435112f
C186 source.t8 a_n3202_n1488# 0.068817f
C187 source.t13 a_n3202_n1488# 0.068817f
C188 source.n27 a_n3202_n1488# 0.436339f
C189 source.n28 a_n3202_n1488# 0.435112f
C190 source.t1 a_n3202_n1488# 0.571445f
C191 source.n29 a_n3202_n1488# 0.440519f
C192 source.t34 a_n3202_n1488# 0.571445f
C193 source.n30 a_n3202_n1488# 0.440519f
C194 source.t30 a_n3202_n1488# 0.068817f
C195 source.t33 a_n3202_n1488# 0.068817f
C196 source.n31 a_n3202_n1488# 0.436339f
C197 source.n32 a_n3202_n1488# 0.435112f
C198 source.t28 a_n3202_n1488# 0.068817f
C199 source.t37 a_n3202_n1488# 0.068817f
C200 source.n33 a_n3202_n1488# 0.436339f
C201 source.n34 a_n3202_n1488# 0.435112f
C202 source.t23 a_n3202_n1488# 0.068817f
C203 source.t36 a_n3202_n1488# 0.068817f
C204 source.n35 a_n3202_n1488# 0.436339f
C205 source.n36 a_n3202_n1488# 0.435112f
C206 source.t24 a_n3202_n1488# 0.068817f
C207 source.t35 a_n3202_n1488# 0.068817f
C208 source.n37 a_n3202_n1488# 0.436339f
C209 source.n38 a_n3202_n1488# 0.435112f
C210 source.t18 a_n3202_n1488# 0.571445f
C211 source.n39 a_n3202_n1488# 0.636157f
C212 source.n40 a_n3202_n1488# 0.859801f
C213 drain_right.t3 a_n3202_n1488# 0.062625f
C214 drain_right.t7 a_n3202_n1488# 0.062625f
C215 drain_right.n0 a_n3202_n1488# 0.456329f
C216 drain_right.t9 a_n3202_n1488# 0.062625f
C217 drain_right.t8 a_n3202_n1488# 0.062625f
C218 drain_right.n1 a_n3202_n1488# 0.451649f
C219 drain_right.n2 a_n3202_n1488# 0.756511f
C220 drain_right.t19 a_n3202_n1488# 0.062625f
C221 drain_right.t11 a_n3202_n1488# 0.062625f
C222 drain_right.n3 a_n3202_n1488# 0.451649f
C223 drain_right.t2 a_n3202_n1488# 0.062625f
C224 drain_right.t18 a_n3202_n1488# 0.062625f
C225 drain_right.n4 a_n3202_n1488# 0.456329f
C226 drain_right.t13 a_n3202_n1488# 0.062625f
C227 drain_right.t12 a_n3202_n1488# 0.062625f
C228 drain_right.n5 a_n3202_n1488# 0.451649f
C229 drain_right.n6 a_n3202_n1488# 0.756512f
C230 drain_right.n7 a_n3202_n1488# 1.43315f
C231 drain_right.t4 a_n3202_n1488# 0.062625f
C232 drain_right.t5 a_n3202_n1488# 0.062625f
C233 drain_right.n8 a_n3202_n1488# 0.456331f
C234 drain_right.t14 a_n3202_n1488# 0.062625f
C235 drain_right.t0 a_n3202_n1488# 0.062625f
C236 drain_right.n9 a_n3202_n1488# 0.451651f
C237 drain_right.n10 a_n3202_n1488# 0.760552f
C238 drain_right.t1 a_n3202_n1488# 0.062625f
C239 drain_right.t16 a_n3202_n1488# 0.062625f
C240 drain_right.n11 a_n3202_n1488# 0.451651f
C241 drain_right.n12 a_n3202_n1488# 0.377296f
C242 drain_right.t17 a_n3202_n1488# 0.062625f
C243 drain_right.t10 a_n3202_n1488# 0.062625f
C244 drain_right.n13 a_n3202_n1488# 0.451651f
C245 drain_right.n14 a_n3202_n1488# 0.377296f
C246 drain_right.t6 a_n3202_n1488# 0.062625f
C247 drain_right.t15 a_n3202_n1488# 0.062625f
C248 drain_right.n15 a_n3202_n1488# 0.451651f
C249 drain_right.n16 a_n3202_n1488# 0.614172f
C250 minus.n0 a_n3202_n1488# 0.039948f
C251 minus.n1 a_n3202_n1488# 0.009065f
C252 minus.t16 a_n3202_n1488# 0.287498f
C253 minus.n2 a_n3202_n1488# 0.066539f
C254 minus.t12 a_n3202_n1488# 0.287498f
C255 minus.n3 a_n3202_n1488# 0.163793f
C256 minus.n4 a_n3202_n1488# 0.039948f
C257 minus.t15 a_n3202_n1488# 0.287498f
C258 minus.n5 a_n3202_n1488# 0.175198f
C259 minus.n6 a_n3202_n1488# 0.183881f
C260 minus.t11 a_n3202_n1488# 0.309931f
C261 minus.n7 a_n3202_n1488# 0.147544f
C262 minus.t8 a_n3202_n1488# 0.287498f
C263 minus.n8 a_n3202_n1488# 0.167151f
C264 minus.n9 a_n3202_n1488# 0.009065f
C265 minus.t6 a_n3202_n1488# 0.287498f
C266 minus.n10 a_n3202_n1488# 0.174706f
C267 minus.n11 a_n3202_n1488# 0.066539f
C268 minus.n12 a_n3202_n1488# 0.066539f
C269 minus.n13 a_n3202_n1488# 0.053306f
C270 minus.n14 a_n3202_n1488# 0.009065f
C271 minus.t17 a_n3202_n1488# 0.287498f
C272 minus.n15 a_n3202_n1488# 0.163793f
C273 minus.n16 a_n3202_n1488# 0.009065f
C274 minus.n17 a_n3202_n1488# 0.039948f
C275 minus.n18 a_n3202_n1488# 0.039948f
C276 minus.n19 a_n3202_n1488# 0.053306f
C277 minus.n20 a_n3202_n1488# 0.009065f
C278 minus.t10 a_n3202_n1488# 0.287498f
C279 minus.n21 a_n3202_n1488# 0.175198f
C280 minus.t18 a_n3202_n1488# 0.287498f
C281 minus.n22 a_n3202_n1488# 0.174706f
C282 minus.n23 a_n3202_n1488# 0.066539f
C283 minus.n24 a_n3202_n1488# 0.053306f
C284 minus.n25 a_n3202_n1488# 0.039948f
C285 minus.n26 a_n3202_n1488# 0.163793f
C286 minus.n27 a_n3202_n1488# 0.009065f
C287 minus.t5 a_n3202_n1488# 0.287498f
C288 minus.n28 a_n3202_n1488# 0.163424f
C289 minus.n29 a_n3202_n1488# 1.32375f
C290 minus.n30 a_n3202_n1488# 0.039948f
C291 minus.n31 a_n3202_n1488# 0.009065f
C292 minus.n32 a_n3202_n1488# 0.066539f
C293 minus.t14 a_n3202_n1488# 0.287498f
C294 minus.n33 a_n3202_n1488# 0.163793f
C295 minus.n34 a_n3202_n1488# 0.039948f
C296 minus.t9 a_n3202_n1488# 0.287498f
C297 minus.n35 a_n3202_n1488# 0.175198f
C298 minus.n36 a_n3202_n1488# 0.183881f
C299 minus.t3 a_n3202_n1488# 0.309931f
C300 minus.n37 a_n3202_n1488# 0.147544f
C301 minus.t7 a_n3202_n1488# 0.287498f
C302 minus.n38 a_n3202_n1488# 0.167151f
C303 minus.n39 a_n3202_n1488# 0.009065f
C304 minus.t4 a_n3202_n1488# 0.287498f
C305 minus.n40 a_n3202_n1488# 0.174706f
C306 minus.n41 a_n3202_n1488# 0.066539f
C307 minus.n42 a_n3202_n1488# 0.066539f
C308 minus.n43 a_n3202_n1488# 0.053306f
C309 minus.n44 a_n3202_n1488# 0.009065f
C310 minus.t0 a_n3202_n1488# 0.287498f
C311 minus.n45 a_n3202_n1488# 0.163793f
C312 minus.n46 a_n3202_n1488# 0.009065f
C313 minus.n47 a_n3202_n1488# 0.039948f
C314 minus.n48 a_n3202_n1488# 0.039948f
C315 minus.n49 a_n3202_n1488# 0.053306f
C316 minus.n50 a_n3202_n1488# 0.009065f
C317 minus.t1 a_n3202_n1488# 0.287498f
C318 minus.n51 a_n3202_n1488# 0.175198f
C319 minus.t13 a_n3202_n1488# 0.287498f
C320 minus.n52 a_n3202_n1488# 0.174706f
C321 minus.n53 a_n3202_n1488# 0.066539f
C322 minus.n54 a_n3202_n1488# 0.053306f
C323 minus.n55 a_n3202_n1488# 0.039948f
C324 minus.t2 a_n3202_n1488# 0.287498f
C325 minus.n56 a_n3202_n1488# 0.163793f
C326 minus.n57 a_n3202_n1488# 0.009065f
C327 minus.t19 a_n3202_n1488# 0.287498f
C328 minus.n58 a_n3202_n1488# 0.163424f
C329 minus.n59 a_n3202_n1488# 0.280288f
C330 minus.n60 a_n3202_n1488# 1.60811f
.ends

