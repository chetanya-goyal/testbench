* NGSPICE file created from diffpair367.ext - technology: sky130A

.subckt diffpair367 minus drain_right drain_left source plus
X0 drain_right.t15 minus.t0 source.t28 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X1 source.t25 minus.t1 drain_right.t14 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X2 drain_left.t15 plus.t0 source.t3 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 drain_left.t14 plus.t1 source.t11 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 source.t20 minus.t2 drain_right.t13 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X5 drain_right.t12 minus.t3 source.t18 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X6 source.t5 plus.t2 drain_left.t13 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X7 drain_right.t11 minus.t4 source.t21 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X8 a_n2210_n2688# a_n2210_n2688# a_n2210_n2688# a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.5
X9 source.t14 plus.t3 drain_left.t12 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X10 drain_right.t10 minus.t5 source.t22 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X11 drain_right.t9 minus.t6 source.t29 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X12 source.t27 minus.t7 drain_right.t8 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X13 drain_left.t11 plus.t4 source.t15 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X14 a_n2210_n2688# a_n2210_n2688# a_n2210_n2688# a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X15 source.t24 minus.t8 drain_right.t7 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X16 drain_right.t6 minus.t9 source.t19 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X17 source.t4 plus.t5 drain_left.t10 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X18 source.t16 minus.t10 drain_right.t5 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X19 source.t17 minus.t11 drain_right.t4 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X20 drain_right.t3 minus.t12 source.t31 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X21 a_n2210_n2688# a_n2210_n2688# a_n2210_n2688# a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X22 drain_left.t9 plus.t6 source.t8 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X23 drain_left.t8 plus.t7 source.t12 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X24 source.t2 plus.t8 drain_left.t7 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X25 source.t26 minus.t13 drain_right.t2 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X26 a_n2210_n2688# a_n2210_n2688# a_n2210_n2688# a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X27 source.t9 plus.t9 drain_left.t6 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X28 source.t0 plus.t10 drain_left.t5 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X29 source.t13 plus.t11 drain_left.t4 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X30 drain_left.t3 plus.t12 source.t1 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X31 drain_left.t2 plus.t13 source.t7 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X32 source.t10 plus.t14 drain_left.t1 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X33 drain_right.t1 minus.t14 source.t23 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X34 source.t30 minus.t15 drain_right.t0 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X35 drain_left.t0 plus.t15 source.t6 a_n2210_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 minus.n5 minus.t12 533.348
R1 minus.n27 minus.t15 533.348
R2 minus.n6 minus.t2 512.366
R3 minus.n8 minus.t6 512.366
R4 minus.n12 minus.t13 512.366
R5 minus.n13 minus.t4 512.366
R6 minus.n1 minus.t10 512.366
R7 minus.n19 minus.t0 512.366
R8 minus.n20 minus.t11 512.366
R9 minus.n28 minus.t14 512.366
R10 minus.n30 minus.t7 512.366
R11 minus.n34 minus.t5 512.366
R12 minus.n35 minus.t1 512.366
R13 minus.n23 minus.t9 512.366
R14 minus.n41 minus.t8 512.366
R15 minus.n42 minus.t3 512.366
R16 minus.n21 minus.n20 161.3
R17 minus.n19 minus.n0 161.3
R18 minus.n18 minus.n17 161.3
R19 minus.n16 minus.n1 161.3
R20 minus.n15 minus.n14 161.3
R21 minus.n13 minus.n2 161.3
R22 minus.n12 minus.n11 161.3
R23 minus.n10 minus.n3 161.3
R24 minus.n9 minus.n8 161.3
R25 minus.n7 minus.n4 161.3
R26 minus.n43 minus.n42 161.3
R27 minus.n41 minus.n22 161.3
R28 minus.n40 minus.n39 161.3
R29 minus.n38 minus.n23 161.3
R30 minus.n37 minus.n36 161.3
R31 minus.n35 minus.n24 161.3
R32 minus.n34 minus.n33 161.3
R33 minus.n32 minus.n25 161.3
R34 minus.n31 minus.n30 161.3
R35 minus.n29 minus.n26 161.3
R36 minus.n5 minus.n4 70.4033
R37 minus.n27 minus.n26 70.4033
R38 minus.n13 minus.n12 48.2005
R39 minus.n20 minus.n19 48.2005
R40 minus.n35 minus.n34 48.2005
R41 minus.n42 minus.n41 48.2005
R42 minus.n8 minus.n7 37.246
R43 minus.n18 minus.n1 37.246
R44 minus.n30 minus.n29 37.246
R45 minus.n40 minus.n23 37.246
R46 minus.n8 minus.n3 35.7853
R47 minus.n14 minus.n1 35.7853
R48 minus.n30 minus.n25 35.7853
R49 minus.n36 minus.n23 35.7853
R50 minus.n44 minus.n21 35.2808
R51 minus.n6 minus.n5 20.9576
R52 minus.n28 minus.n27 20.9576
R53 minus.n12 minus.n3 12.4157
R54 minus.n14 minus.n13 12.4157
R55 minus.n34 minus.n25 12.4157
R56 minus.n36 minus.n35 12.4157
R57 minus.n7 minus.n6 10.955
R58 minus.n19 minus.n18 10.955
R59 minus.n29 minus.n28 10.955
R60 minus.n41 minus.n40 10.955
R61 minus.n44 minus.n43 6.56111
R62 minus.n21 minus.n0 0.189894
R63 minus.n17 minus.n0 0.189894
R64 minus.n17 minus.n16 0.189894
R65 minus.n16 minus.n15 0.189894
R66 minus.n15 minus.n2 0.189894
R67 minus.n11 minus.n2 0.189894
R68 minus.n11 minus.n10 0.189894
R69 minus.n10 minus.n9 0.189894
R70 minus.n9 minus.n4 0.189894
R71 minus.n31 minus.n26 0.189894
R72 minus.n32 minus.n31 0.189894
R73 minus.n33 minus.n32 0.189894
R74 minus.n33 minus.n24 0.189894
R75 minus.n37 minus.n24 0.189894
R76 minus.n38 minus.n37 0.189894
R77 minus.n39 minus.n38 0.189894
R78 minus.n39 minus.n22 0.189894
R79 minus.n43 minus.n22 0.189894
R80 minus minus.n44 0.188
R81 source.n7 source.t5 51.0588
R82 source.n8 source.t31 51.0588
R83 source.n15 source.t17 51.0588
R84 source.n31 source.t18 51.0586
R85 source.n24 source.t30 51.0586
R86 source.n23 source.t12 51.0586
R87 source.n16 source.t9 51.0586
R88 source.n0 source.t7 51.0586
R89 source.n2 source.n1 48.8588
R90 source.n4 source.n3 48.8588
R91 source.n6 source.n5 48.8588
R92 source.n10 source.n9 48.8588
R93 source.n12 source.n11 48.8588
R94 source.n14 source.n13 48.8588
R95 source.n30 source.n29 48.8586
R96 source.n28 source.n27 48.8586
R97 source.n26 source.n25 48.8586
R98 source.n22 source.n21 48.8586
R99 source.n20 source.n19 48.8586
R100 source.n18 source.n17 48.8586
R101 source.n16 source.n15 19.7305
R102 source.n32 source.n0 14.1098
R103 source.n32 source.n31 5.62119
R104 source.n29 source.t19 2.2005
R105 source.n29 source.t24 2.2005
R106 source.n27 source.t22 2.2005
R107 source.n27 source.t25 2.2005
R108 source.n25 source.t23 2.2005
R109 source.n25 source.t27 2.2005
R110 source.n21 source.t11 2.2005
R111 source.n21 source.t2 2.2005
R112 source.n19 source.t1 2.2005
R113 source.n19 source.t13 2.2005
R114 source.n17 source.t3 2.2005
R115 source.n17 source.t14 2.2005
R116 source.n1 source.t6 2.2005
R117 source.n1 source.t4 2.2005
R118 source.n3 source.t15 2.2005
R119 source.n3 source.t0 2.2005
R120 source.n5 source.t8 2.2005
R121 source.n5 source.t10 2.2005
R122 source.n9 source.t29 2.2005
R123 source.n9 source.t20 2.2005
R124 source.n11 source.t21 2.2005
R125 source.n11 source.t26 2.2005
R126 source.n13 source.t28 2.2005
R127 source.n13 source.t16 2.2005
R128 source.n15 source.n14 0.716017
R129 source.n14 source.n12 0.716017
R130 source.n12 source.n10 0.716017
R131 source.n10 source.n8 0.716017
R132 source.n7 source.n6 0.716017
R133 source.n6 source.n4 0.716017
R134 source.n4 source.n2 0.716017
R135 source.n2 source.n0 0.716017
R136 source.n18 source.n16 0.716017
R137 source.n20 source.n18 0.716017
R138 source.n22 source.n20 0.716017
R139 source.n23 source.n22 0.716017
R140 source.n26 source.n24 0.716017
R141 source.n28 source.n26 0.716017
R142 source.n30 source.n28 0.716017
R143 source.n31 source.n30 0.716017
R144 source.n8 source.n7 0.470328
R145 source.n24 source.n23 0.470328
R146 source source.n32 0.188
R147 drain_right.n9 drain_right.n7 66.2529
R148 drain_right.n5 drain_right.n3 66.2529
R149 drain_right.n2 drain_right.n0 66.2529
R150 drain_right.n9 drain_right.n8 65.5376
R151 drain_right.n11 drain_right.n10 65.5376
R152 drain_right.n13 drain_right.n12 65.5376
R153 drain_right.n5 drain_right.n4 65.5373
R154 drain_right.n2 drain_right.n1 65.5373
R155 drain_right drain_right.n6 29.192
R156 drain_right drain_right.n13 6.36873
R157 drain_right.n3 drain_right.t7 2.2005
R158 drain_right.n3 drain_right.t12 2.2005
R159 drain_right.n4 drain_right.t14 2.2005
R160 drain_right.n4 drain_right.t6 2.2005
R161 drain_right.n1 drain_right.t8 2.2005
R162 drain_right.n1 drain_right.t10 2.2005
R163 drain_right.n0 drain_right.t0 2.2005
R164 drain_right.n0 drain_right.t1 2.2005
R165 drain_right.n7 drain_right.t13 2.2005
R166 drain_right.n7 drain_right.t3 2.2005
R167 drain_right.n8 drain_right.t2 2.2005
R168 drain_right.n8 drain_right.t9 2.2005
R169 drain_right.n10 drain_right.t5 2.2005
R170 drain_right.n10 drain_right.t11 2.2005
R171 drain_right.n12 drain_right.t4 2.2005
R172 drain_right.n12 drain_right.t15 2.2005
R173 drain_right.n13 drain_right.n11 0.716017
R174 drain_right.n11 drain_right.n9 0.716017
R175 drain_right.n6 drain_right.n5 0.302913
R176 drain_right.n6 drain_right.n2 0.302913
R177 plus.n5 plus.t2 533.348
R178 plus.n27 plus.t7 533.348
R179 plus.n20 plus.t13 512.366
R180 plus.n19 plus.t5 512.366
R181 plus.n1 plus.t15 512.366
R182 plus.n13 plus.t10 512.366
R183 plus.n12 plus.t4 512.366
R184 plus.n4 plus.t14 512.366
R185 plus.n6 plus.t6 512.366
R186 plus.n42 plus.t9 512.366
R187 plus.n41 plus.t0 512.366
R188 plus.n23 plus.t3 512.366
R189 plus.n35 plus.t12 512.366
R190 plus.n34 plus.t11 512.366
R191 plus.n26 plus.t1 512.366
R192 plus.n28 plus.t8 512.366
R193 plus.n8 plus.n7 161.3
R194 plus.n9 plus.n4 161.3
R195 plus.n11 plus.n10 161.3
R196 plus.n12 plus.n3 161.3
R197 plus.n13 plus.n2 161.3
R198 plus.n15 plus.n14 161.3
R199 plus.n16 plus.n1 161.3
R200 plus.n18 plus.n17 161.3
R201 plus.n19 plus.n0 161.3
R202 plus.n21 plus.n20 161.3
R203 plus.n30 plus.n29 161.3
R204 plus.n31 plus.n26 161.3
R205 plus.n33 plus.n32 161.3
R206 plus.n34 plus.n25 161.3
R207 plus.n35 plus.n24 161.3
R208 plus.n37 plus.n36 161.3
R209 plus.n38 plus.n23 161.3
R210 plus.n40 plus.n39 161.3
R211 plus.n41 plus.n22 161.3
R212 plus.n43 plus.n42 161.3
R213 plus.n8 plus.n5 70.4033
R214 plus.n30 plus.n27 70.4033
R215 plus.n20 plus.n19 48.2005
R216 plus.n13 plus.n12 48.2005
R217 plus.n42 plus.n41 48.2005
R218 plus.n35 plus.n34 48.2005
R219 plus.n18 plus.n1 37.246
R220 plus.n7 plus.n4 37.246
R221 plus.n40 plus.n23 37.246
R222 plus.n29 plus.n26 37.246
R223 plus.n14 plus.n1 35.7853
R224 plus.n11 plus.n4 35.7853
R225 plus.n36 plus.n23 35.7853
R226 plus.n33 plus.n26 35.7853
R227 plus plus.n43 30.2983
R228 plus.n6 plus.n5 20.9576
R229 plus.n28 plus.n27 20.9576
R230 plus.n14 plus.n13 12.4157
R231 plus.n12 plus.n11 12.4157
R232 plus.n36 plus.n35 12.4157
R233 plus.n34 plus.n33 12.4157
R234 plus plus.n21 11.0687
R235 plus.n19 plus.n18 10.955
R236 plus.n7 plus.n6 10.955
R237 plus.n41 plus.n40 10.955
R238 plus.n29 plus.n28 10.955
R239 plus.n9 plus.n8 0.189894
R240 plus.n10 plus.n9 0.189894
R241 plus.n10 plus.n3 0.189894
R242 plus.n3 plus.n2 0.189894
R243 plus.n15 plus.n2 0.189894
R244 plus.n16 plus.n15 0.189894
R245 plus.n17 plus.n16 0.189894
R246 plus.n17 plus.n0 0.189894
R247 plus.n21 plus.n0 0.189894
R248 plus.n43 plus.n22 0.189894
R249 plus.n39 plus.n22 0.189894
R250 plus.n39 plus.n38 0.189894
R251 plus.n38 plus.n37 0.189894
R252 plus.n37 plus.n24 0.189894
R253 plus.n25 plus.n24 0.189894
R254 plus.n32 plus.n25 0.189894
R255 plus.n32 plus.n31 0.189894
R256 plus.n31 plus.n30 0.189894
R257 drain_left.n9 drain_left.n7 66.2531
R258 drain_left.n5 drain_left.n3 66.2529
R259 drain_left.n2 drain_left.n0 66.2529
R260 drain_left.n11 drain_left.n10 65.5376
R261 drain_left.n9 drain_left.n8 65.5376
R262 drain_left.n13 drain_left.n12 65.5374
R263 drain_left.n5 drain_left.n4 65.5373
R264 drain_left.n2 drain_left.n1 65.5373
R265 drain_left drain_left.n6 29.7452
R266 drain_left drain_left.n13 6.36873
R267 drain_left.n3 drain_left.t7 2.2005
R268 drain_left.n3 drain_left.t8 2.2005
R269 drain_left.n4 drain_left.t4 2.2005
R270 drain_left.n4 drain_left.t14 2.2005
R271 drain_left.n1 drain_left.t12 2.2005
R272 drain_left.n1 drain_left.t3 2.2005
R273 drain_left.n0 drain_left.t6 2.2005
R274 drain_left.n0 drain_left.t15 2.2005
R275 drain_left.n12 drain_left.t10 2.2005
R276 drain_left.n12 drain_left.t2 2.2005
R277 drain_left.n10 drain_left.t5 2.2005
R278 drain_left.n10 drain_left.t0 2.2005
R279 drain_left.n8 drain_left.t1 2.2005
R280 drain_left.n8 drain_left.t11 2.2005
R281 drain_left.n7 drain_left.t13 2.2005
R282 drain_left.n7 drain_left.t9 2.2005
R283 drain_left.n11 drain_left.n9 0.716017
R284 drain_left.n13 drain_left.n11 0.716017
R285 drain_left.n6 drain_left.n5 0.302913
R286 drain_left.n6 drain_left.n2 0.302913
C0 plus drain_left 6.62409f
C1 plus source 6.41499f
C2 drain_right drain_left 1.15071f
C3 drain_right source 18.4298f
C4 minus drain_left 0.172419f
C5 minus source 6.40095f
C6 source drain_left 18.4286f
C7 drain_right plus 0.372806f
C8 minus plus 5.35108f
C9 drain_right minus 6.40692f
C10 drain_right a_n2210_n2688# 5.96854f
C11 drain_left a_n2210_n2688# 6.29199f
C12 source a_n2210_n2688# 7.344686f
C13 minus a_n2210_n2688# 8.538036f
C14 plus a_n2210_n2688# 10.230089f
C15 drain_left.t6 a_n2210_n2688# 0.207589f
C16 drain_left.t15 a_n2210_n2688# 0.207589f
C17 drain_left.n0 a_n2210_n2688# 1.81981f
C18 drain_left.t12 a_n2210_n2688# 0.207589f
C19 drain_left.t3 a_n2210_n2688# 0.207589f
C20 drain_left.n1 a_n2210_n2688# 1.81571f
C21 drain_left.n2 a_n2210_n2688# 0.707818f
C22 drain_left.t7 a_n2210_n2688# 0.207589f
C23 drain_left.t8 a_n2210_n2688# 0.207589f
C24 drain_left.n3 a_n2210_n2688# 1.81981f
C25 drain_left.t4 a_n2210_n2688# 0.207589f
C26 drain_left.t14 a_n2210_n2688# 0.207589f
C27 drain_left.n4 a_n2210_n2688# 1.81571f
C28 drain_left.n5 a_n2210_n2688# 0.707818f
C29 drain_left.n6 a_n2210_n2688# 1.35604f
C30 drain_left.t13 a_n2210_n2688# 0.207589f
C31 drain_left.t9 a_n2210_n2688# 0.207589f
C32 drain_left.n7 a_n2210_n2688# 1.81982f
C33 drain_left.t1 a_n2210_n2688# 0.207589f
C34 drain_left.t11 a_n2210_n2688# 0.207589f
C35 drain_left.n8 a_n2210_n2688# 1.81571f
C36 drain_left.n9 a_n2210_n2688# 0.744426f
C37 drain_left.t5 a_n2210_n2688# 0.207589f
C38 drain_left.t0 a_n2210_n2688# 0.207589f
C39 drain_left.n10 a_n2210_n2688# 1.81571f
C40 drain_left.n11 a_n2210_n2688# 0.368387f
C41 drain_left.t10 a_n2210_n2688# 0.207589f
C42 drain_left.t2 a_n2210_n2688# 0.207589f
C43 drain_left.n12 a_n2210_n2688# 1.8157f
C44 drain_left.n13 a_n2210_n2688# 0.619163f
C45 plus.n0 a_n2210_n2688# 0.04598f
C46 plus.t13 a_n2210_n2688# 0.593394f
C47 plus.t5 a_n2210_n2688# 0.593394f
C48 plus.t15 a_n2210_n2688# 0.593394f
C49 plus.n1 a_n2210_n2688# 0.257722f
C50 plus.n2 a_n2210_n2688# 0.04598f
C51 plus.t10 a_n2210_n2688# 0.593394f
C52 plus.t4 a_n2210_n2688# 0.593394f
C53 plus.n3 a_n2210_n2688# 0.04598f
C54 plus.t14 a_n2210_n2688# 0.593394f
C55 plus.n4 a_n2210_n2688# 0.257722f
C56 plus.t2 a_n2210_n2688# 0.603346f
C57 plus.n5 a_n2210_n2688# 0.243286f
C58 plus.t6 a_n2210_n2688# 0.593394f
C59 plus.n6 a_n2210_n2688# 0.255029f
C60 plus.n7 a_n2210_n2688# 0.010434f
C61 plus.n8 a_n2210_n2688# 0.146394f
C62 plus.n9 a_n2210_n2688# 0.04598f
C63 plus.n10 a_n2210_n2688# 0.04598f
C64 plus.n11 a_n2210_n2688# 0.010434f
C65 plus.n12 a_n2210_n2688# 0.255313f
C66 plus.n13 a_n2210_n2688# 0.255313f
C67 plus.n14 a_n2210_n2688# 0.010434f
C68 plus.n15 a_n2210_n2688# 0.04598f
C69 plus.n16 a_n2210_n2688# 0.04598f
C70 plus.n17 a_n2210_n2688# 0.04598f
C71 plus.n18 a_n2210_n2688# 0.010434f
C72 plus.n19 a_n2210_n2688# 0.255029f
C73 plus.n20 a_n2210_n2688# 0.252903f
C74 plus.n21 a_n2210_n2688# 0.458468f
C75 plus.n22 a_n2210_n2688# 0.04598f
C76 plus.t9 a_n2210_n2688# 0.593394f
C77 plus.t0 a_n2210_n2688# 0.593394f
C78 plus.t3 a_n2210_n2688# 0.593394f
C79 plus.n23 a_n2210_n2688# 0.257722f
C80 plus.n24 a_n2210_n2688# 0.04598f
C81 plus.t12 a_n2210_n2688# 0.593394f
C82 plus.n25 a_n2210_n2688# 0.04598f
C83 plus.t11 a_n2210_n2688# 0.593394f
C84 plus.t1 a_n2210_n2688# 0.593394f
C85 plus.n26 a_n2210_n2688# 0.257722f
C86 plus.t7 a_n2210_n2688# 0.603346f
C87 plus.n27 a_n2210_n2688# 0.243286f
C88 plus.t8 a_n2210_n2688# 0.593394f
C89 plus.n28 a_n2210_n2688# 0.255029f
C90 plus.n29 a_n2210_n2688# 0.010434f
C91 plus.n30 a_n2210_n2688# 0.146394f
C92 plus.n31 a_n2210_n2688# 0.04598f
C93 plus.n32 a_n2210_n2688# 0.04598f
C94 plus.n33 a_n2210_n2688# 0.010434f
C95 plus.n34 a_n2210_n2688# 0.255313f
C96 plus.n35 a_n2210_n2688# 0.255313f
C97 plus.n36 a_n2210_n2688# 0.010434f
C98 plus.n37 a_n2210_n2688# 0.04598f
C99 plus.n38 a_n2210_n2688# 0.04598f
C100 plus.n39 a_n2210_n2688# 0.04598f
C101 plus.n40 a_n2210_n2688# 0.010434f
C102 plus.n41 a_n2210_n2688# 0.255029f
C103 plus.n42 a_n2210_n2688# 0.252903f
C104 plus.n43 a_n2210_n2688# 1.36677f
C105 drain_right.t0 a_n2210_n2688# 0.206873f
C106 drain_right.t1 a_n2210_n2688# 0.206873f
C107 drain_right.n0 a_n2210_n2688# 1.81354f
C108 drain_right.t8 a_n2210_n2688# 0.206873f
C109 drain_right.t10 a_n2210_n2688# 0.206873f
C110 drain_right.n1 a_n2210_n2688# 1.80945f
C111 drain_right.n2 a_n2210_n2688# 0.705377f
C112 drain_right.t7 a_n2210_n2688# 0.206873f
C113 drain_right.t12 a_n2210_n2688# 0.206873f
C114 drain_right.n3 a_n2210_n2688# 1.81354f
C115 drain_right.t14 a_n2210_n2688# 0.206873f
C116 drain_right.t6 a_n2210_n2688# 0.206873f
C117 drain_right.n4 a_n2210_n2688# 1.80945f
C118 drain_right.n5 a_n2210_n2688# 0.705377f
C119 drain_right.n6 a_n2210_n2688# 1.29186f
C120 drain_right.t13 a_n2210_n2688# 0.206873f
C121 drain_right.t3 a_n2210_n2688# 0.206873f
C122 drain_right.n7 a_n2210_n2688# 1.81353f
C123 drain_right.t2 a_n2210_n2688# 0.206873f
C124 drain_right.t9 a_n2210_n2688# 0.206873f
C125 drain_right.n8 a_n2210_n2688# 1.80945f
C126 drain_right.n9 a_n2210_n2688# 0.741866f
C127 drain_right.t5 a_n2210_n2688# 0.206873f
C128 drain_right.t11 a_n2210_n2688# 0.206873f
C129 drain_right.n10 a_n2210_n2688# 1.80945f
C130 drain_right.n11 a_n2210_n2688# 0.367117f
C131 drain_right.t4 a_n2210_n2688# 0.206873f
C132 drain_right.t15 a_n2210_n2688# 0.206873f
C133 drain_right.n12 a_n2210_n2688# 1.80945f
C134 drain_right.n13 a_n2210_n2688# 0.61702f
C135 source.t7 a_n2210_n2688# 1.91591f
C136 source.n0 a_n2210_n2688# 1.12518f
C137 source.t6 a_n2210_n2688# 0.17967f
C138 source.t4 a_n2210_n2688# 0.17967f
C139 source.n1 a_n2210_n2688# 1.50408f
C140 source.n2 a_n2210_n2688# 0.351942f
C141 source.t15 a_n2210_n2688# 0.17967f
C142 source.t0 a_n2210_n2688# 0.17967f
C143 source.n3 a_n2210_n2688# 1.50408f
C144 source.n4 a_n2210_n2688# 0.351942f
C145 source.t8 a_n2210_n2688# 0.17967f
C146 source.t10 a_n2210_n2688# 0.17967f
C147 source.n5 a_n2210_n2688# 1.50408f
C148 source.n6 a_n2210_n2688# 0.351942f
C149 source.t5 a_n2210_n2688# 1.91591f
C150 source.n7 a_n2210_n2688# 0.410122f
C151 source.t31 a_n2210_n2688# 1.91591f
C152 source.n8 a_n2210_n2688# 0.410122f
C153 source.t29 a_n2210_n2688# 0.17967f
C154 source.t20 a_n2210_n2688# 0.17967f
C155 source.n9 a_n2210_n2688# 1.50408f
C156 source.n10 a_n2210_n2688# 0.351942f
C157 source.t21 a_n2210_n2688# 0.17967f
C158 source.t26 a_n2210_n2688# 0.17967f
C159 source.n11 a_n2210_n2688# 1.50408f
C160 source.n12 a_n2210_n2688# 0.351942f
C161 source.t28 a_n2210_n2688# 0.17967f
C162 source.t16 a_n2210_n2688# 0.17967f
C163 source.n13 a_n2210_n2688# 1.50408f
C164 source.n14 a_n2210_n2688# 0.351942f
C165 source.t17 a_n2210_n2688# 1.91591f
C166 source.n15 a_n2210_n2688# 1.49683f
C167 source.t9 a_n2210_n2688# 1.91591f
C168 source.n16 a_n2210_n2688# 1.49684f
C169 source.t3 a_n2210_n2688# 0.17967f
C170 source.t14 a_n2210_n2688# 0.17967f
C171 source.n17 a_n2210_n2688# 1.50408f
C172 source.n18 a_n2210_n2688# 0.351947f
C173 source.t1 a_n2210_n2688# 0.17967f
C174 source.t13 a_n2210_n2688# 0.17967f
C175 source.n19 a_n2210_n2688# 1.50408f
C176 source.n20 a_n2210_n2688# 0.351947f
C177 source.t11 a_n2210_n2688# 0.17967f
C178 source.t2 a_n2210_n2688# 0.17967f
C179 source.n21 a_n2210_n2688# 1.50408f
C180 source.n22 a_n2210_n2688# 0.351947f
C181 source.t12 a_n2210_n2688# 1.91591f
C182 source.n23 a_n2210_n2688# 0.410127f
C183 source.t30 a_n2210_n2688# 1.91591f
C184 source.n24 a_n2210_n2688# 0.410127f
C185 source.t23 a_n2210_n2688# 0.17967f
C186 source.t27 a_n2210_n2688# 0.17967f
C187 source.n25 a_n2210_n2688# 1.50408f
C188 source.n26 a_n2210_n2688# 0.351947f
C189 source.t22 a_n2210_n2688# 0.17967f
C190 source.t25 a_n2210_n2688# 0.17967f
C191 source.n27 a_n2210_n2688# 1.50408f
C192 source.n28 a_n2210_n2688# 0.351947f
C193 source.t19 a_n2210_n2688# 0.17967f
C194 source.t24 a_n2210_n2688# 0.17967f
C195 source.n29 a_n2210_n2688# 1.50408f
C196 source.n30 a_n2210_n2688# 0.351947f
C197 source.t18 a_n2210_n2688# 1.91591f
C198 source.n31 a_n2210_n2688# 0.563888f
C199 source.n32 a_n2210_n2688# 1.32257f
C200 minus.n0 a_n2210_n2688# 0.045252f
C201 minus.t10 a_n2210_n2688# 0.583993f
C202 minus.n1 a_n2210_n2688# 0.253639f
C203 minus.n2 a_n2210_n2688# 0.045252f
C204 minus.n3 a_n2210_n2688# 0.010269f
C205 minus.t13 a_n2210_n2688# 0.583993f
C206 minus.n4 a_n2210_n2688# 0.144075f
C207 minus.t2 a_n2210_n2688# 0.583993f
C208 minus.t12 a_n2210_n2688# 0.593787f
C209 minus.n5 a_n2210_n2688# 0.239432f
C210 minus.n6 a_n2210_n2688# 0.250989f
C211 minus.n7 a_n2210_n2688# 0.010269f
C212 minus.t6 a_n2210_n2688# 0.583993f
C213 minus.n8 a_n2210_n2688# 0.253639f
C214 minus.n9 a_n2210_n2688# 0.045252f
C215 minus.n10 a_n2210_n2688# 0.045252f
C216 minus.n11 a_n2210_n2688# 0.045252f
C217 minus.n12 a_n2210_n2688# 0.251268f
C218 minus.t4 a_n2210_n2688# 0.583993f
C219 minus.n13 a_n2210_n2688# 0.251268f
C220 minus.n14 a_n2210_n2688# 0.010269f
C221 minus.n15 a_n2210_n2688# 0.045252f
C222 minus.n16 a_n2210_n2688# 0.045252f
C223 minus.n17 a_n2210_n2688# 0.045252f
C224 minus.n18 a_n2210_n2688# 0.010269f
C225 minus.t0 a_n2210_n2688# 0.583993f
C226 minus.n19 a_n2210_n2688# 0.250989f
C227 minus.t11 a_n2210_n2688# 0.583993f
C228 minus.n20 a_n2210_n2688# 0.248896f
C229 minus.n21 a_n2210_n2688# 1.53847f
C230 minus.n22 a_n2210_n2688# 0.045252f
C231 minus.t9 a_n2210_n2688# 0.583993f
C232 minus.n23 a_n2210_n2688# 0.253639f
C233 minus.n24 a_n2210_n2688# 0.045252f
C234 minus.n25 a_n2210_n2688# 0.010269f
C235 minus.n26 a_n2210_n2688# 0.144075f
C236 minus.t15 a_n2210_n2688# 0.593787f
C237 minus.n27 a_n2210_n2688# 0.239432f
C238 minus.t14 a_n2210_n2688# 0.583993f
C239 minus.n28 a_n2210_n2688# 0.250989f
C240 minus.n29 a_n2210_n2688# 0.010269f
C241 minus.t7 a_n2210_n2688# 0.583993f
C242 minus.n30 a_n2210_n2688# 0.253639f
C243 minus.n31 a_n2210_n2688# 0.045252f
C244 minus.n32 a_n2210_n2688# 0.045252f
C245 minus.n33 a_n2210_n2688# 0.045252f
C246 minus.t5 a_n2210_n2688# 0.583993f
C247 minus.n34 a_n2210_n2688# 0.251268f
C248 minus.t1 a_n2210_n2688# 0.583993f
C249 minus.n35 a_n2210_n2688# 0.251268f
C250 minus.n36 a_n2210_n2688# 0.010269f
C251 minus.n37 a_n2210_n2688# 0.045252f
C252 minus.n38 a_n2210_n2688# 0.045252f
C253 minus.n39 a_n2210_n2688# 0.045252f
C254 minus.n40 a_n2210_n2688# 0.010269f
C255 minus.t8 a_n2210_n2688# 0.583993f
C256 minus.n41 a_n2210_n2688# 0.250989f
C257 minus.t3 a_n2210_n2688# 0.583993f
C258 minus.n42 a_n2210_n2688# 0.248896f
C259 minus.n43 a_n2210_n2688# 0.302341f
C260 minus.n44 a_n2210_n2688# 1.87143f
.ends

