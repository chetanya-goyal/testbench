* NGSPICE file created from diffpair564.ext - technology: sky130A

.subckt diffpair564 minus drain_right drain_left source plus
X0 a_n1496_n4888# a_n1496_n4888# a_n1496_n4888# a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=76 ps=327.6 w=20 l=0.15
X1 source.t15 minus.t0 drain_right.t9 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X2 drain_right.t1 minus.t1 source.t14 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X3 a_n1496_n4888# a_n1496_n4888# a_n1496_n4888# a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X4 drain_left.t9 plus.t0 source.t2 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X5 a_n1496_n4888# a_n1496_n4888# a_n1496_n4888# a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X6 source.t13 minus.t2 drain_right.t3 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X7 source.t16 plus.t1 drain_left.t8 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X8 drain_right.t0 minus.t3 source.t12 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X9 drain_right.t7 minus.t4 source.t11 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X10 drain_right.t6 minus.t5 source.t10 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X11 source.t9 minus.t6 drain_right.t5 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X12 drain_left.t7 plus.t2 source.t1 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X13 drain_left.t6 plus.t3 source.t4 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X14 drain_right.t4 minus.t7 source.t8 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X15 a_n1496_n4888# a_n1496_n4888# a_n1496_n4888# a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X16 source.t7 minus.t8 drain_right.t8 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X17 drain_left.t5 plus.t4 source.t5 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X18 source.t18 plus.t5 drain_left.t4 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X19 drain_left.t3 plus.t6 source.t17 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X20 source.t0 plus.t7 drain_left.t2 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X21 source.t19 plus.t8 drain_left.t1 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X22 drain_right.t2 minus.t9 source.t6 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X23 drain_left.t0 plus.t9 source.t3 a_n1496_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
R0 minus.n9 minus.t4 3466.02
R1 minus.n3 minus.t3 3466.02
R2 minus.n20 minus.t5 3466.02
R3 minus.n14 minus.t1 3466.02
R4 minus.n6 minus.t7 3422.2
R5 minus.n8 minus.t6 3422.2
R6 minus.n2 minus.t2 3422.2
R7 minus.n17 minus.t9 3422.2
R8 minus.n19 minus.t0 3422.2
R9 minus.n13 minus.t8 3422.2
R10 minus.n4 minus.n3 161.489
R11 minus.n15 minus.n14 161.489
R12 minus.n10 minus.n9 161.3
R13 minus.n7 minus.n0 161.3
R14 minus.n6 minus.n5 161.3
R15 minus.n4 minus.n1 161.3
R16 minus.n21 minus.n20 161.3
R17 minus.n18 minus.n11 161.3
R18 minus.n17 minus.n16 161.3
R19 minus.n15 minus.n12 161.3
R20 minus.n7 minus.n6 73.0308
R21 minus.n6 minus.n1 73.0308
R22 minus.n17 minus.n12 73.0308
R23 minus.n18 minus.n17 73.0308
R24 minus.n9 minus.n8 51.1217
R25 minus.n3 minus.n2 51.1217
R26 minus.n14 minus.n13 51.1217
R27 minus.n20 minus.n19 51.1217
R28 minus.n22 minus.n10 40.8622
R29 minus.n8 minus.n7 21.9096
R30 minus.n2 minus.n1 21.9096
R31 minus.n13 minus.n12 21.9096
R32 minus.n19 minus.n18 21.9096
R33 minus.n22 minus.n21 6.51376
R34 minus.n10 minus.n0 0.189894
R35 minus.n5 minus.n0 0.189894
R36 minus.n5 minus.n4 0.189894
R37 minus.n16 minus.n15 0.189894
R38 minus.n16 minus.n11 0.189894
R39 minus.n21 minus.n11 0.189894
R40 minus minus.n22 0.188
R41 drain_right.n1 drain_right.t1 61.8786
R42 drain_right.n7 drain_right.t7 61.3184
R43 drain_right.n6 drain_right.n4 60.3788
R44 drain_right.n3 drain_right.n2 60.1833
R45 drain_right.n6 drain_right.n5 59.8185
R46 drain_right.n1 drain_right.n0 59.8184
R47 drain_right drain_right.n3 35.2559
R48 drain_right drain_right.n7 5.93339
R49 drain_right.n2 drain_right.t9 1.5005
R50 drain_right.n2 drain_right.t6 1.5005
R51 drain_right.n0 drain_right.t8 1.5005
R52 drain_right.n0 drain_right.t2 1.5005
R53 drain_right.n4 drain_right.t3 1.5005
R54 drain_right.n4 drain_right.t0 1.5005
R55 drain_right.n5 drain_right.t5 1.5005
R56 drain_right.n5 drain_right.t4 1.5005
R57 drain_right.n7 drain_right.n6 0.560845
R58 drain_right.n3 drain_right.n1 0.0852402
R59 source.n0 source.t3 44.6397
R60 source.n5 source.t12 44.6396
R61 source.n19 source.t10 44.6395
R62 source.n14 source.t1 44.6395
R63 source.n2 source.n1 43.1397
R64 source.n4 source.n3 43.1397
R65 source.n7 source.n6 43.1397
R66 source.n9 source.n8 43.1397
R67 source.n18 source.n17 43.1396
R68 source.n16 source.n15 43.1396
R69 source.n13 source.n12 43.1396
R70 source.n11 source.n10 43.1396
R71 source.n11 source.n9 28.469
R72 source.n20 source.n0 22.3656
R73 source.n20 source.n19 5.5436
R74 source.n17 source.t6 1.5005
R75 source.n17 source.t15 1.5005
R76 source.n15 source.t14 1.5005
R77 source.n15 source.t7 1.5005
R78 source.n12 source.t2 1.5005
R79 source.n12 source.t0 1.5005
R80 source.n10 source.t5 1.5005
R81 source.n10 source.t16 1.5005
R82 source.n1 source.t17 1.5005
R83 source.n1 source.t18 1.5005
R84 source.n3 source.t4 1.5005
R85 source.n3 source.t19 1.5005
R86 source.n6 source.t8 1.5005
R87 source.n6 source.t13 1.5005
R88 source.n8 source.t11 1.5005
R89 source.n8 source.t9 1.5005
R90 source.n5 source.n4 0.7505
R91 source.n16 source.n14 0.7505
R92 source.n9 source.n7 0.560845
R93 source.n7 source.n5 0.560845
R94 source.n4 source.n2 0.560845
R95 source.n2 source.n0 0.560845
R96 source.n13 source.n11 0.560845
R97 source.n14 source.n13 0.560845
R98 source.n18 source.n16 0.560845
R99 source.n19 source.n18 0.560845
R100 source source.n20 0.188
R101 plus.n3 plus.t3 3466.02
R102 plus.n9 plus.t9 3466.02
R103 plus.n14 plus.t2 3466.02
R104 plus.n20 plus.t4 3466.02
R105 plus.n6 plus.t6 3422.2
R106 plus.n2 plus.t8 3422.2
R107 plus.n8 plus.t5 3422.2
R108 plus.n17 plus.t0 3422.2
R109 plus.n13 plus.t7 3422.2
R110 plus.n19 plus.t1 3422.2
R111 plus.n4 plus.n3 161.489
R112 plus.n15 plus.n14 161.489
R113 plus.n4 plus.n1 161.3
R114 plus.n6 plus.n5 161.3
R115 plus.n7 plus.n0 161.3
R116 plus.n10 plus.n9 161.3
R117 plus.n15 plus.n12 161.3
R118 plus.n17 plus.n16 161.3
R119 plus.n18 plus.n11 161.3
R120 plus.n21 plus.n20 161.3
R121 plus.n6 plus.n1 73.0308
R122 plus.n7 plus.n6 73.0308
R123 plus.n18 plus.n17 73.0308
R124 plus.n17 plus.n12 73.0308
R125 plus.n3 plus.n2 51.1217
R126 plus.n9 plus.n8 51.1217
R127 plus.n20 plus.n19 51.1217
R128 plus.n14 plus.n13 51.1217
R129 plus plus.n21 31.713
R130 plus.n2 plus.n1 21.9096
R131 plus.n8 plus.n7 21.9096
R132 plus.n19 plus.n18 21.9096
R133 plus.n13 plus.n12 21.9096
R134 plus plus.n10 15.188
R135 plus.n5 plus.n4 0.189894
R136 plus.n5 plus.n0 0.189894
R137 plus.n10 plus.n0 0.189894
R138 plus.n21 plus.n11 0.189894
R139 plus.n16 plus.n11 0.189894
R140 plus.n16 plus.n15 0.189894
R141 drain_left.n5 drain_left.t6 61.8788
R142 drain_left.n1 drain_left.t5 61.8786
R143 drain_left.n3 drain_left.n2 60.1833
R144 drain_left.n7 drain_left.n6 59.8185
R145 drain_left.n5 drain_left.n4 59.8185
R146 drain_left.n1 drain_left.n0 59.8184
R147 drain_left drain_left.n3 35.8091
R148 drain_left drain_left.n7 6.21356
R149 drain_left.n2 drain_left.t2 1.5005
R150 drain_left.n2 drain_left.t7 1.5005
R151 drain_left.n0 drain_left.t8 1.5005
R152 drain_left.n0 drain_left.t9 1.5005
R153 drain_left.n6 drain_left.t4 1.5005
R154 drain_left.n6 drain_left.t0 1.5005
R155 drain_left.n4 drain_left.t1 1.5005
R156 drain_left.n4 drain_left.t3 1.5005
R157 drain_left.n7 drain_left.n5 0.560845
R158 drain_left.n3 drain_left.n1 0.0852402
C0 plus drain_left 4.07437f
C1 drain_right minus 3.93606f
C2 source plus 3.03486f
C3 plus minus 6.48496f
C4 drain_right plus 0.300059f
C5 source drain_left 34.3126f
C6 minus drain_left 0.170828f
C7 drain_right drain_left 0.739657f
C8 source minus 3.01975f
C9 drain_right source 34.2954f
C10 drain_right a_n1496_n4888# 8.763481f
C11 drain_left a_n1496_n4888# 9.00537f
C12 source a_n1496_n4888# 8.945076f
C13 minus a_n1496_n4888# 6.040097f
C14 plus a_n1496_n4888# 8.83965f
C15 drain_left.t5 a_n1496_n4888# 5.0775f
C16 drain_left.t8 a_n1496_n4888# 0.609125f
C17 drain_left.t9 a_n1496_n4888# 0.609125f
C18 drain_left.n0 a_n1496_n4888# 4.08958f
C19 drain_left.n1 a_n1496_n4888# 0.653823f
C20 drain_left.t2 a_n1496_n4888# 0.609125f
C21 drain_left.t7 a_n1496_n4888# 0.609125f
C22 drain_left.n2 a_n1496_n4888# 4.09142f
C23 drain_left.n3 a_n1496_n4888# 1.95166f
C24 drain_left.t6 a_n1496_n4888# 5.07752f
C25 drain_left.t1 a_n1496_n4888# 0.609125f
C26 drain_left.t3 a_n1496_n4888# 0.609125f
C27 drain_left.n4 a_n1496_n4888# 4.08958f
C28 drain_left.n5 a_n1496_n4888# 0.685834f
C29 drain_left.t4 a_n1496_n4888# 0.609125f
C30 drain_left.t0 a_n1496_n4888# 0.609125f
C31 drain_left.n6 a_n1496_n4888# 4.08958f
C32 drain_left.n7 a_n1496_n4888# 0.51894f
C33 plus.n0 a_n1496_n4888# 0.059558f
C34 plus.t5 a_n1496_n4888# 0.503228f
C35 plus.t6 a_n1496_n4888# 0.503228f
C36 plus.n1 a_n1496_n4888# 0.025265f
C37 plus.t3 a_n1496_n4888# 0.505685f
C38 plus.t8 a_n1496_n4888# 0.503228f
C39 plus.n2 a_n1496_n4888# 0.196117f
C40 plus.n3 a_n1496_n4888# 0.217171f
C41 plus.n4 a_n1496_n4888# 0.128215f
C42 plus.n5 a_n1496_n4888# 0.059558f
C43 plus.n6 a_n1496_n4888# 0.215874f
C44 plus.n7 a_n1496_n4888# 0.025265f
C45 plus.n8 a_n1496_n4888# 0.196117f
C46 plus.t9 a_n1496_n4888# 0.505685f
C47 plus.n9 a_n1496_n4888# 0.21709f
C48 plus.n10 a_n1496_n4888# 0.906226f
C49 plus.n11 a_n1496_n4888# 0.059558f
C50 plus.t4 a_n1496_n4888# 0.505685f
C51 plus.t1 a_n1496_n4888# 0.503228f
C52 plus.t0 a_n1496_n4888# 0.503228f
C53 plus.n12 a_n1496_n4888# 0.025265f
C54 plus.t7 a_n1496_n4888# 0.503228f
C55 plus.n13 a_n1496_n4888# 0.196117f
C56 plus.t2 a_n1496_n4888# 0.505685f
C57 plus.n14 a_n1496_n4888# 0.217171f
C58 plus.n15 a_n1496_n4888# 0.128215f
C59 plus.n16 a_n1496_n4888# 0.059558f
C60 plus.n17 a_n1496_n4888# 0.215874f
C61 plus.n18 a_n1496_n4888# 0.025265f
C62 plus.n19 a_n1496_n4888# 0.196117f
C63 plus.n20 a_n1496_n4888# 0.21709f
C64 plus.n21 a_n1496_n4888# 1.99395f
C65 source.t3 a_n1496_n4888# 4.9592f
C66 source.n0 a_n1496_n4888# 2.01345f
C67 source.t17 a_n1496_n4888# 0.609788f
C68 source.t18 a_n1496_n4888# 0.609788f
C69 source.n1 a_n1496_n4888# 4.01282f
C70 source.n2 a_n1496_n4888# 0.353444f
C71 source.t4 a_n1496_n4888# 0.609788f
C72 source.t19 a_n1496_n4888# 0.609788f
C73 source.n3 a_n1496_n4888# 4.01282f
C74 source.n4 a_n1496_n4888# 0.369005f
C75 source.t12 a_n1496_n4888# 4.95921f
C76 source.n5 a_n1496_n4888# 0.52023f
C77 source.t8 a_n1496_n4888# 0.609788f
C78 source.t13 a_n1496_n4888# 0.609788f
C79 source.n6 a_n1496_n4888# 4.01282f
C80 source.n7 a_n1496_n4888# 0.353444f
C81 source.t11 a_n1496_n4888# 0.609788f
C82 source.t9 a_n1496_n4888# 0.609788f
C83 source.n8 a_n1496_n4888# 4.01282f
C84 source.n9 a_n1496_n4888# 2.36007f
C85 source.t5 a_n1496_n4888# 0.609788f
C86 source.t16 a_n1496_n4888# 0.609788f
C87 source.n10 a_n1496_n4888# 4.01283f
C88 source.n11 a_n1496_n4888# 2.36006f
C89 source.t2 a_n1496_n4888# 0.609788f
C90 source.t0 a_n1496_n4888# 0.609788f
C91 source.n12 a_n1496_n4888# 4.01283f
C92 source.n13 a_n1496_n4888# 0.353436f
C93 source.t1 a_n1496_n4888# 4.95919f
C94 source.n14 a_n1496_n4888# 0.520255f
C95 source.t14 a_n1496_n4888# 0.609788f
C96 source.t7 a_n1496_n4888# 0.609788f
C97 source.n15 a_n1496_n4888# 4.01283f
C98 source.n16 a_n1496_n4888# 0.368998f
C99 source.t6 a_n1496_n4888# 0.609788f
C100 source.t15 a_n1496_n4888# 0.609788f
C101 source.n17 a_n1496_n4888# 4.01283f
C102 source.n18 a_n1496_n4888# 0.353436f
C103 source.t10 a_n1496_n4888# 4.95919f
C104 source.n19 a_n1496_n4888# 0.642144f
C105 source.n20 a_n1496_n4888# 2.29319f
C106 drain_right.t1 a_n1496_n4888# 5.06418f
C107 drain_right.t8 a_n1496_n4888# 0.607527f
C108 drain_right.t2 a_n1496_n4888# 0.607527f
C109 drain_right.n0 a_n1496_n4888# 4.07885f
C110 drain_right.n1 a_n1496_n4888# 0.652108f
C111 drain_right.t9 a_n1496_n4888# 0.607527f
C112 drain_right.t6 a_n1496_n4888# 0.607527f
C113 drain_right.n2 a_n1496_n4888# 4.08068f
C114 drain_right.n3 a_n1496_n4888# 1.89345f
C115 drain_right.t3 a_n1496_n4888# 0.607527f
C116 drain_right.t0 a_n1496_n4888# 0.607527f
C117 drain_right.n4 a_n1496_n4888# 4.08178f
C118 drain_right.t5 a_n1496_n4888# 0.607527f
C119 drain_right.t4 a_n1496_n4888# 0.607527f
C120 drain_right.n5 a_n1496_n4888# 4.07885f
C121 drain_right.n6 a_n1496_n4888# 0.618705f
C122 drain_right.t7 a_n1496_n4888# 5.06074f
C123 drain_right.n7 a_n1496_n4888# 0.594519f
C124 minus.n0 a_n1496_n4888# 0.058167f
C125 minus.t4 a_n1496_n4888# 0.493874f
C126 minus.t6 a_n1496_n4888# 0.491476f
C127 minus.t7 a_n1496_n4888# 0.491476f
C128 minus.n1 a_n1496_n4888# 0.024675f
C129 minus.t2 a_n1496_n4888# 0.491476f
C130 minus.n2 a_n1496_n4888# 0.191537f
C131 minus.t3 a_n1496_n4888# 0.493874f
C132 minus.n3 a_n1496_n4888# 0.212099f
C133 minus.n4 a_n1496_n4888# 0.12522f
C134 minus.n5 a_n1496_n4888# 0.058167f
C135 minus.n6 a_n1496_n4888# 0.210833f
C136 minus.n7 a_n1496_n4888# 0.024675f
C137 minus.n8 a_n1496_n4888# 0.191537f
C138 minus.n9 a_n1496_n4888# 0.21202f
C139 minus.n10 a_n1496_n4888# 2.47392f
C140 minus.n11 a_n1496_n4888# 0.058167f
C141 minus.t0 a_n1496_n4888# 0.491476f
C142 minus.t9 a_n1496_n4888# 0.491476f
C143 minus.n12 a_n1496_n4888# 0.024675f
C144 minus.t1 a_n1496_n4888# 0.493874f
C145 minus.t8 a_n1496_n4888# 0.491476f
C146 minus.n13 a_n1496_n4888# 0.191537f
C147 minus.n14 a_n1496_n4888# 0.212099f
C148 minus.n15 a_n1496_n4888# 0.12522f
C149 minus.n16 a_n1496_n4888# 0.058167f
C150 minus.n17 a_n1496_n4888# 0.210833f
C151 minus.n18 a_n1496_n4888# 0.024675f
C152 minus.n19 a_n1496_n4888# 0.191537f
C153 minus.t5 a_n1496_n4888# 0.493874f
C154 minus.n20 a_n1496_n4888# 0.21202f
C155 minus.n21 a_n1496_n4888# 0.382163f
C156 minus.n22 a_n1496_n4888# 2.96351f
.ends

