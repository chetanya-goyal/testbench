* NGSPICE file created from diffpair73.ext - technology: sky130A

.subckt diffpair73 minus drain_right drain_left source plus
X0 a_n1846_n1088# a_n1846_n1088# a_n1846_n1088# a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.8
X1 a_n1846_n1088# a_n1846_n1088# a_n1846_n1088# a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X2 source.t15 minus.t0 drain_right.t7 a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X3 source.t14 minus.t1 drain_right.t5 a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X4 drain_right.t0 minus.t2 source.t13 a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X5 drain_left.t7 plus.t0 source.t2 a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X6 drain_left.t6 plus.t1 source.t6 a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X7 source.t12 minus.t3 drain_right.t3 a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X8 drain_right.t1 minus.t4 source.t11 a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X9 a_n1846_n1088# a_n1846_n1088# a_n1846_n1088# a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X10 source.t10 minus.t5 drain_right.t6 a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X11 a_n1846_n1088# a_n1846_n1088# a_n1846_n1088# a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X12 drain_left.t5 plus.t2 source.t7 a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X13 drain_right.t4 minus.t6 source.t9 a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X14 drain_right.t2 minus.t7 source.t8 a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X15 source.t1 plus.t3 drain_left.t4 a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X16 drain_left.t3 plus.t4 source.t3 a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X17 source.t5 plus.t5 drain_left.t2 a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X18 source.t0 plus.t6 drain_left.t1 a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X19 source.t4 plus.t7 drain_left.t0 a_n1846_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
R0 minus.n7 minus.n6 161.3
R1 minus.n5 minus.n0 161.3
R2 minus.n15 minus.n14 161.3
R3 minus.n13 minus.n8 161.3
R4 minus.n2 minus.t4 99.8318
R5 minus.n10 minus.t1 99.8318
R6 minus.n4 minus.n3 80.6037
R7 minus.n12 minus.n11 80.6037
R8 minus.n1 minus.t3 79.2293
R9 minus.n4 minus.t2 79.2293
R10 minus.n6 minus.t5 79.2293
R11 minus.n9 minus.t7 79.2293
R12 minus.n12 minus.t0 79.2293
R13 minus.n14 minus.t6 79.2293
R14 minus.n4 minus.n1 48.2005
R15 minus.n12 minus.n9 48.2005
R16 minus.n5 minus.n4 41.6278
R17 minus.n13 minus.n12 41.6278
R18 minus.n3 minus.n2 31.6158
R19 minus.n11 minus.n10 31.6158
R20 minus.n16 minus.n7 27.9323
R21 minus.n2 minus.n1 17.6494
R22 minus.n10 minus.n9 17.6494
R23 minus.n16 minus.n15 6.65202
R24 minus.n6 minus.n5 6.57323
R25 minus.n14 minus.n13 6.57323
R26 minus.n3 minus.n0 0.285035
R27 minus.n11 minus.n8 0.285035
R28 minus.n7 minus.n0 0.189894
R29 minus.n15 minus.n8 0.189894
R30 minus minus.n16 0.188
R31 drain_right.n5 drain_right.n3 241.107
R32 drain_right.n2 drain_right.n1 240.564
R33 drain_right.n2 drain_right.n0 240.564
R34 drain_right.n5 drain_right.n4 240.132
R35 drain_right drain_right.n2 21.89
R36 drain_right.n1 drain_right.t7 19.8005
R37 drain_right.n1 drain_right.t4 19.8005
R38 drain_right.n0 drain_right.t5 19.8005
R39 drain_right.n0 drain_right.t2 19.8005
R40 drain_right.n3 drain_right.t3 19.8005
R41 drain_right.n3 drain_right.t1 19.8005
R42 drain_right.n4 drain_right.t6 19.8005
R43 drain_right.n4 drain_right.t0 19.8005
R44 drain_right drain_right.n5 6.62735
R45 source.n0 source.t7 243.255
R46 source.n3 source.t0 243.255
R47 source.n4 source.t11 243.255
R48 source.n7 source.t10 243.255
R49 source.n15 source.t9 243.254
R50 source.n12 source.t14 243.254
R51 source.n11 source.t2 243.254
R52 source.n8 source.t4 243.254
R53 source.n2 source.n1 223.454
R54 source.n6 source.n5 223.454
R55 source.n14 source.n13 223.453
R56 source.n10 source.n9 223.453
R57 source.n13 source.t8 19.8005
R58 source.n13 source.t15 19.8005
R59 source.n9 source.t6 19.8005
R60 source.n9 source.t5 19.8005
R61 source.n1 source.t3 19.8005
R62 source.n1 source.t1 19.8005
R63 source.n5 source.t13 19.8005
R64 source.n5 source.t12 19.8005
R65 source.n8 source.n7 13.9285
R66 source.n16 source.n0 8.17853
R67 source.n16 source.n15 5.7505
R68 source.n7 source.n6 0.974638
R69 source.n6 source.n4 0.974638
R70 source.n3 source.n2 0.974638
R71 source.n2 source.n0 0.974638
R72 source.n10 source.n8 0.974638
R73 source.n11 source.n10 0.974638
R74 source.n14 source.n12 0.974638
R75 source.n15 source.n14 0.974638
R76 source.n4 source.n3 0.470328
R77 source.n12 source.n11 0.470328
R78 source source.n16 0.188
R79 plus.n5 plus.n0 161.3
R80 plus.n7 plus.n6 161.3
R81 plus.n13 plus.n8 161.3
R82 plus.n15 plus.n14 161.3
R83 plus.n2 plus.t6 99.8318
R84 plus.n10 plus.t0 99.8318
R85 plus.n4 plus.n1 80.6037
R86 plus.n12 plus.n9 80.6037
R87 plus.n6 plus.t2 79.2293
R88 plus.n4 plus.t3 79.2293
R89 plus.n3 plus.t4 79.2293
R90 plus.n14 plus.t7 79.2293
R91 plus.n12 plus.t1 79.2293
R92 plus.n11 plus.t5 79.2293
R93 plus.n4 plus.n3 48.2005
R94 plus.n12 plus.n11 48.2005
R95 plus.n5 plus.n4 41.6278
R96 plus.n13 plus.n12 41.6278
R97 plus.n2 plus.n1 31.6158
R98 plus.n10 plus.n9 31.6158
R99 plus plus.n15 25.9801
R100 plus.n3 plus.n2 17.6494
R101 plus.n11 plus.n10 17.6494
R102 plus plus.n7 8.12929
R103 plus.n6 plus.n5 6.57323
R104 plus.n14 plus.n13 6.57323
R105 plus.n1 plus.n0 0.285035
R106 plus.n9 plus.n8 0.285035
R107 plus.n7 plus.n0 0.189894
R108 plus.n15 plus.n8 0.189894
R109 drain_left.n5 drain_left.n3 241.107
R110 drain_left.n2 drain_left.n1 240.564
R111 drain_left.n2 drain_left.n0 240.564
R112 drain_left.n5 drain_left.n4 240.132
R113 drain_left drain_left.n2 22.4432
R114 drain_left.n1 drain_left.t2 19.8005
R115 drain_left.n1 drain_left.t7 19.8005
R116 drain_left.n0 drain_left.t0 19.8005
R117 drain_left.n0 drain_left.t6 19.8005
R118 drain_left.n4 drain_left.t4 19.8005
R119 drain_left.n4 drain_left.t5 19.8005
R120 drain_left.n3 drain_left.t1 19.8005
R121 drain_left.n3 drain_left.t3 19.8005
R122 drain_left drain_left.n5 6.62735
C0 drain_right drain_left 0.873777f
C1 drain_left plus 1.0362f
C2 source drain_left 2.96049f
C3 minus drain_right 0.857095f
C4 minus plus 3.4154f
C5 source minus 1.26458f
C6 drain_right plus 0.342228f
C7 source drain_right 2.96287f
C8 source plus 1.27845f
C9 minus drain_left 0.178628f
C10 drain_right a_n1846_n1088# 3.246674f
C11 drain_left a_n1846_n1088# 3.469461f
C12 source a_n1846_n1088# 2.484419f
C13 minus a_n1846_n1088# 6.243483f
C14 plus a_n1846_n1088# 6.859413f
C15 drain_left.t0 a_n1846_n1088# 0.015001f
C16 drain_left.t6 a_n1846_n1088# 0.015001f
C17 drain_left.n0 a_n1846_n1088# 0.058696f
C18 drain_left.t2 a_n1846_n1088# 0.015001f
C19 drain_left.t7 a_n1846_n1088# 0.015001f
C20 drain_left.n1 a_n1846_n1088# 0.058696f
C21 drain_left.n2 a_n1846_n1088# 0.986895f
C22 drain_left.t1 a_n1846_n1088# 0.015001f
C23 drain_left.t3 a_n1846_n1088# 0.015001f
C24 drain_left.n3 a_n1846_n1088# 0.059337f
C25 drain_left.t4 a_n1846_n1088# 0.015001f
C26 drain_left.t5 a_n1846_n1088# 0.015001f
C27 drain_left.n4 a_n1846_n1088# 0.058288f
C28 drain_left.n5 a_n1846_n1088# 0.680649f
C29 plus.n0 a_n1846_n1088# 0.039292f
C30 plus.t2 a_n1846_n1088# 0.07988f
C31 plus.t3 a_n1846_n1088# 0.07988f
C32 plus.n1 a_n1846_n1088# 0.168528f
C33 plus.t4 a_n1846_n1088# 0.07988f
C34 plus.t6 a_n1846_n1088# 0.096265f
C35 plus.n2 a_n1846_n1088# 0.065473f
C36 plus.n3 a_n1846_n1088# 0.085425f
C37 plus.n4 a_n1846_n1088# 0.084945f
C38 plus.n5 a_n1846_n1088# 0.006682f
C39 plus.n6 a_n1846_n1088# 0.073906f
C40 plus.n7 a_n1846_n1088# 0.212921f
C41 plus.n8 a_n1846_n1088# 0.039292f
C42 plus.t7 a_n1846_n1088# 0.07988f
C43 plus.n9 a_n1846_n1088# 0.168528f
C44 plus.t1 a_n1846_n1088# 0.07988f
C45 plus.t0 a_n1846_n1088# 0.096265f
C46 plus.n10 a_n1846_n1088# 0.065473f
C47 plus.t5 a_n1846_n1088# 0.07988f
C48 plus.n11 a_n1846_n1088# 0.085425f
C49 plus.n12 a_n1846_n1088# 0.084945f
C50 plus.n13 a_n1846_n1088# 0.006682f
C51 plus.n14 a_n1846_n1088# 0.073906f
C52 plus.n15 a_n1846_n1088# 0.660615f
C53 source.t7 a_n1846_n1088# 0.09884f
C54 source.n0 a_n1846_n1088# 0.480096f
C55 source.t3 a_n1846_n1088# 0.017758f
C56 source.t1 a_n1846_n1088# 0.017758f
C57 source.n1 a_n1846_n1088# 0.057593f
C58 source.n2 a_n1846_n1088# 0.279094f
C59 source.t0 a_n1846_n1088# 0.09884f
C60 source.n3 a_n1846_n1088# 0.249761f
C61 source.t11 a_n1846_n1088# 0.09884f
C62 source.n4 a_n1846_n1088# 0.249761f
C63 source.t13 a_n1846_n1088# 0.017758f
C64 source.t12 a_n1846_n1088# 0.017758f
C65 source.n5 a_n1846_n1088# 0.057593f
C66 source.n6 a_n1846_n1088# 0.279094f
C67 source.t10 a_n1846_n1088# 0.09884f
C68 source.n7 a_n1846_n1088# 0.6669f
C69 source.t4 a_n1846_n1088# 0.09884f
C70 source.n8 a_n1846_n1088# 0.6669f
C71 source.t6 a_n1846_n1088# 0.017758f
C72 source.t5 a_n1846_n1088# 0.017758f
C73 source.n9 a_n1846_n1088# 0.057593f
C74 source.n10 a_n1846_n1088# 0.279095f
C75 source.t2 a_n1846_n1088# 0.09884f
C76 source.n11 a_n1846_n1088# 0.249762f
C77 source.t14 a_n1846_n1088# 0.09884f
C78 source.n12 a_n1846_n1088# 0.249762f
C79 source.t8 a_n1846_n1088# 0.017758f
C80 source.t15 a_n1846_n1088# 0.017758f
C81 source.n13 a_n1846_n1088# 0.057593f
C82 source.n14 a_n1846_n1088# 0.279095f
C83 source.t9 a_n1846_n1088# 0.09884f
C84 source.n15 a_n1846_n1088# 0.401215f
C85 source.n16 a_n1846_n1088# 0.468474f
C86 drain_right.t5 a_n1846_n1088# 0.015381f
C87 drain_right.t2 a_n1846_n1088# 0.015381f
C88 drain_right.n0 a_n1846_n1088# 0.060186f
C89 drain_right.t7 a_n1846_n1088# 0.015381f
C90 drain_right.t4 a_n1846_n1088# 0.015381f
C91 drain_right.n1 a_n1846_n1088# 0.060186f
C92 drain_right.n2 a_n1846_n1088# 0.974316f
C93 drain_right.t3 a_n1846_n1088# 0.015381f
C94 drain_right.t1 a_n1846_n1088# 0.015381f
C95 drain_right.n3 a_n1846_n1088# 0.060843f
C96 drain_right.t6 a_n1846_n1088# 0.015381f
C97 drain_right.t0 a_n1846_n1088# 0.015381f
C98 drain_right.n4 a_n1846_n1088# 0.059768f
C99 drain_right.n5 a_n1846_n1088# 0.697925f
C100 minus.n0 a_n1846_n1088# 0.038615f
C101 minus.t3 a_n1846_n1088# 0.078505f
C102 minus.n1 a_n1846_n1088# 0.083954f
C103 minus.t2 a_n1846_n1088# 0.078505f
C104 minus.t4 a_n1846_n1088# 0.094608f
C105 minus.n2 a_n1846_n1088# 0.064346f
C106 minus.n3 a_n1846_n1088# 0.165628f
C107 minus.n4 a_n1846_n1088# 0.083483f
C108 minus.n5 a_n1846_n1088# 0.006567f
C109 minus.t5 a_n1846_n1088# 0.078505f
C110 minus.n6 a_n1846_n1088# 0.072634f
C111 minus.n7 a_n1846_n1088# 0.669272f
C112 minus.n8 a_n1846_n1088# 0.038615f
C113 minus.t7 a_n1846_n1088# 0.078505f
C114 minus.n9 a_n1846_n1088# 0.083954f
C115 minus.t1 a_n1846_n1088# 0.094608f
C116 minus.n10 a_n1846_n1088# 0.064346f
C117 minus.n11 a_n1846_n1088# 0.165628f
C118 minus.t0 a_n1846_n1088# 0.078505f
C119 minus.n12 a_n1846_n1088# 0.083483f
C120 minus.n13 a_n1846_n1088# 0.006567f
C121 minus.t6 a_n1846_n1088# 0.078505f
C122 minus.n14 a_n1846_n1088# 0.072634f
C123 minus.n15 a_n1846_n1088# 0.199486f
C124 minus.n16 a_n1846_n1088# 0.821537f
.ends

