* NGSPICE file created from diffpair354.ext - technology: sky130A

.subckt diffpair354 minus drain_right drain_left source plus
X0 drain_left.t9 plus.t0 source.t17 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X1 drain_right.t9 minus.t0 source.t1 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X2 a_n1472_n2688# a_n1472_n2688# a_n1472_n2688# a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.3
X3 drain_left.t8 plus.t1 source.t18 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X4 drain_right.t8 minus.t1 source.t3 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X5 source.t10 plus.t2 drain_left.t7 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X6 a_n1472_n2688# a_n1472_n2688# a_n1472_n2688# a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X7 drain_left.t6 plus.t3 source.t12 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X8 source.t14 plus.t4 drain_left.t5 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X9 source.t19 plus.t5 drain_left.t4 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X10 source.t4 minus.t2 drain_right.t7 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X11 source.t0 minus.t3 drain_right.t6 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X12 source.t7 minus.t4 drain_right.t5 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X13 a_n1472_n2688# a_n1472_n2688# a_n1472_n2688# a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X14 drain_right.t4 minus.t5 source.t5 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X15 drain_left.t3 plus.t6 source.t11 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X16 drain_left.t2 plus.t7 source.t13 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X17 drain_left.t1 plus.t8 source.t16 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X18 a_n1472_n2688# a_n1472_n2688# a_n1472_n2688# a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X19 drain_right.t3 minus.t6 source.t9 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X20 source.t2 minus.t7 drain_right.t2 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X21 drain_right.t1 minus.t8 source.t6 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X22 drain_right.t0 minus.t9 source.t8 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X23 source.t15 plus.t9 drain_left.t0 a_n1472_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
R0 plus.n3 plus.t1 865.409
R1 plus.n9 plus.t3 865.409
R2 plus.n14 plus.t6 865.409
R3 plus.n20 plus.t0 865.409
R4 plus.n6 plus.t7 827.433
R5 plus.n2 plus.t5 827.433
R6 plus.n8 plus.t9 827.433
R7 plus.n17 plus.t8 827.433
R8 plus.n13 plus.t2 827.433
R9 plus.n19 plus.t4 827.433
R10 plus.n4 plus.n3 161.489
R11 plus.n15 plus.n14 161.489
R12 plus.n4 plus.n1 161.3
R13 plus.n6 plus.n5 161.3
R14 plus.n7 plus.n0 161.3
R15 plus.n10 plus.n9 161.3
R16 plus.n15 plus.n12 161.3
R17 plus.n17 plus.n16 161.3
R18 plus.n18 plus.n11 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n6 plus.n1 73.0308
R21 plus.n7 plus.n6 73.0308
R22 plus.n18 plus.n17 73.0308
R23 plus.n17 plus.n12 73.0308
R24 plus.n3 plus.n2 54.0429
R25 plus.n9 plus.n8 54.0429
R26 plus.n20 plus.n19 54.0429
R27 plus.n14 plus.n13 54.0429
R28 plus plus.n21 27.4289
R29 plus.n2 plus.n1 18.9884
R30 plus.n8 plus.n7 18.9884
R31 plus.n19 plus.n18 18.9884
R32 plus.n13 plus.n12 18.9884
R33 plus plus.n10 10.9948
R34 plus.n5 plus.n4 0.189894
R35 plus.n5 plus.n0 0.189894
R36 plus.n10 plus.n0 0.189894
R37 plus.n21 plus.n11 0.189894
R38 plus.n16 plus.n11 0.189894
R39 plus.n16 plus.n15 0.189894
R40 source.n5 source.t5 51.0588
R41 source.n19 source.t3 51.0586
R42 source.n14 source.t11 51.0586
R43 source.n0 source.t12 51.0586
R44 source.n2 source.n1 48.8588
R45 source.n4 source.n3 48.8588
R46 source.n7 source.n6 48.8588
R47 source.n9 source.n8 48.8588
R48 source.n18 source.n17 48.8586
R49 source.n16 source.n15 48.8586
R50 source.n13 source.n12 48.8586
R51 source.n11 source.n10 48.8586
R52 source.n11 source.n9 20.1012
R53 source.n20 source.n0 14.0236
R54 source.n20 source.n19 5.53498
R55 source.n17 source.t6 2.2005
R56 source.n17 source.t4 2.2005
R57 source.n15 source.t8 2.2005
R58 source.n15 source.t0 2.2005
R59 source.n12 source.t16 2.2005
R60 source.n12 source.t10 2.2005
R61 source.n10 source.t17 2.2005
R62 source.n10 source.t14 2.2005
R63 source.n1 source.t13 2.2005
R64 source.n1 source.t15 2.2005
R65 source.n3 source.t18 2.2005
R66 source.n3 source.t19 2.2005
R67 source.n6 source.t1 2.2005
R68 source.n6 source.t2 2.2005
R69 source.n8 source.t9 2.2005
R70 source.n8 source.t7 2.2005
R71 source.n5 source.n4 0.741879
R72 source.n16 source.n14 0.741879
R73 source.n9 source.n7 0.543603
R74 source.n7 source.n5 0.543603
R75 source.n4 source.n2 0.543603
R76 source.n2 source.n0 0.543603
R77 source.n13 source.n11 0.543603
R78 source.n14 source.n13 0.543603
R79 source.n18 source.n16 0.543603
R80 source.n19 source.n18 0.543603
R81 source source.n20 0.188
R82 drain_left.n5 drain_left.t8 68.2807
R83 drain_left.n1 drain_left.t9 68.2804
R84 drain_left.n3 drain_left.n2 65.8893
R85 drain_left.n5 drain_left.n4 65.5376
R86 drain_left.n7 drain_left.n6 65.5374
R87 drain_left.n1 drain_left.n0 65.5373
R88 drain_left drain_left.n3 27.4025
R89 drain_left drain_left.n7 6.19632
R90 drain_left.n2 drain_left.t7 2.2005
R91 drain_left.n2 drain_left.t3 2.2005
R92 drain_left.n0 drain_left.t5 2.2005
R93 drain_left.n0 drain_left.t1 2.2005
R94 drain_left.n6 drain_left.t0 2.2005
R95 drain_left.n6 drain_left.t6 2.2005
R96 drain_left.n4 drain_left.t4 2.2005
R97 drain_left.n4 drain_left.t2 2.2005
R98 drain_left.n7 drain_left.n5 0.543603
R99 drain_left.n3 drain_left.n1 0.0809298
R100 minus.n9 minus.t6 865.409
R101 minus.n3 minus.t5 865.409
R102 minus.n20 minus.t1 865.409
R103 minus.n14 minus.t9 865.409
R104 minus.n6 minus.t0 827.433
R105 minus.n8 minus.t4 827.433
R106 minus.n2 minus.t7 827.433
R107 minus.n17 minus.t8 827.433
R108 minus.n19 minus.t2 827.433
R109 minus.n13 minus.t3 827.433
R110 minus.n4 minus.n3 161.489
R111 minus.n15 minus.n14 161.489
R112 minus.n10 minus.n9 161.3
R113 minus.n7 minus.n0 161.3
R114 minus.n6 minus.n5 161.3
R115 minus.n4 minus.n1 161.3
R116 minus.n21 minus.n20 161.3
R117 minus.n18 minus.n11 161.3
R118 minus.n17 minus.n16 161.3
R119 minus.n15 minus.n12 161.3
R120 minus.n7 minus.n6 73.0308
R121 minus.n6 minus.n1 73.0308
R122 minus.n17 minus.n12 73.0308
R123 minus.n18 minus.n17 73.0308
R124 minus.n9 minus.n8 54.0429
R125 minus.n3 minus.n2 54.0429
R126 minus.n14 minus.n13 54.0429
R127 minus.n20 minus.n19 54.0429
R128 minus.n22 minus.n10 32.4115
R129 minus.n8 minus.n7 18.9884
R130 minus.n2 minus.n1 18.9884
R131 minus.n13 minus.n12 18.9884
R132 minus.n19 minus.n18 18.9884
R133 minus.n22 minus.n21 6.48724
R134 minus.n10 minus.n0 0.189894
R135 minus.n5 minus.n0 0.189894
R136 minus.n5 minus.n4 0.189894
R137 minus.n16 minus.n15 0.189894
R138 minus.n16 minus.n11 0.189894
R139 minus.n21 minus.n11 0.189894
R140 minus minus.n22 0.188
R141 drain_right.n1 drain_right.t0 68.2804
R142 drain_right.n7 drain_right.t3 67.7376
R143 drain_right.n6 drain_right.n4 66.0805
R144 drain_right.n3 drain_right.n2 65.8893
R145 drain_right.n6 drain_right.n5 65.5376
R146 drain_right.n1 drain_right.n0 65.5373
R147 drain_right drain_right.n3 26.8493
R148 drain_right drain_right.n7 5.92477
R149 drain_right.n2 drain_right.t7 2.2005
R150 drain_right.n2 drain_right.t8 2.2005
R151 drain_right.n0 drain_right.t6 2.2005
R152 drain_right.n0 drain_right.t1 2.2005
R153 drain_right.n4 drain_right.t2 2.2005
R154 drain_right.n4 drain_right.t4 2.2005
R155 drain_right.n5 drain_right.t5 2.2005
R156 drain_right.n5 drain_right.t9 2.2005
R157 drain_right.n7 drain_right.n6 0.543603
R158 drain_right.n3 drain_right.n1 0.0809298
C0 plus minus 4.4323f
C1 drain_right plus 0.296114f
C2 source drain_left 16.3248f
C3 minus drain_left 0.171269f
C4 drain_right drain_left 0.723546f
C5 source minus 2.82482f
C6 drain_right source 16.3162f
C7 plus drain_left 3.23346f
C8 drain_right minus 3.09517f
C9 source plus 2.83935f
C10 drain_right a_n1472_n2688# 5.981639f
C11 drain_left a_n1472_n2688# 6.22002f
C12 source a_n1472_n2688# 5.055253f
C13 minus a_n1472_n2688# 5.490043f
C14 plus a_n1472_n2688# 7.239951f
C15 drain_right.t0 a_n1472_n2688# 2.33394f
C16 drain_right.t6 a_n1472_n2688# 0.209363f
C17 drain_right.t1 a_n1472_n2688# 0.209363f
C18 drain_right.n0 a_n1472_n2688# 1.83123f
C19 drain_right.n1 a_n1472_n2688# 0.670876f
C20 drain_right.t7 a_n1472_n2688# 0.209363f
C21 drain_right.t8 a_n1472_n2688# 0.209363f
C22 drain_right.n2 a_n1472_n2688# 1.83301f
C23 drain_right.n3 a_n1472_n2688# 1.39686f
C24 drain_right.t2 a_n1472_n2688# 0.209363f
C25 drain_right.t4 a_n1472_n2688# 0.209363f
C26 drain_right.n4 a_n1472_n2688# 1.83411f
C27 drain_right.t5 a_n1472_n2688# 0.209363f
C28 drain_right.t9 a_n1472_n2688# 0.209363f
C29 drain_right.n5 a_n1472_n2688# 1.83123f
C30 drain_right.n6 a_n1472_n2688# 0.686637f
C31 drain_right.t3 a_n1472_n2688# 2.331f
C32 drain_right.n7 a_n1472_n2688# 0.615972f
C33 minus.n0 a_n1472_n2688# 0.053074f
C34 minus.t6 a_n1472_n2688# 0.413585f
C35 minus.t4 a_n1472_n2688# 0.406058f
C36 minus.t0 a_n1472_n2688# 0.406058f
C37 minus.n1 a_n1472_n2688# 0.021861f
C38 minus.t7 a_n1472_n2688# 0.406058f
C39 minus.n2 a_n1472_n2688# 0.169563f
C40 minus.t5 a_n1472_n2688# 0.413585f
C41 minus.n3 a_n1472_n2688# 0.185934f
C42 minus.n4 a_n1472_n2688# 0.116546f
C43 minus.n5 a_n1472_n2688# 0.053074f
C44 minus.n6 a_n1472_n2688# 0.187169f
C45 minus.n7 a_n1472_n2688# 0.021861f
C46 minus.n8 a_n1472_n2688# 0.169563f
C47 minus.n9 a_n1472_n2688# 0.18586f
C48 minus.n10 a_n1472_n2688# 1.57102f
C49 minus.n11 a_n1472_n2688# 0.053074f
C50 minus.t2 a_n1472_n2688# 0.406058f
C51 minus.t8 a_n1472_n2688# 0.406058f
C52 minus.n12 a_n1472_n2688# 0.021861f
C53 minus.t9 a_n1472_n2688# 0.413585f
C54 minus.t3 a_n1472_n2688# 0.406058f
C55 minus.n13 a_n1472_n2688# 0.169563f
C56 minus.n14 a_n1472_n2688# 0.185934f
C57 minus.n15 a_n1472_n2688# 0.116546f
C58 minus.n16 a_n1472_n2688# 0.053074f
C59 minus.n17 a_n1472_n2688# 0.187169f
C60 minus.n18 a_n1472_n2688# 0.021861f
C61 minus.n19 a_n1472_n2688# 0.169563f
C62 minus.t1 a_n1472_n2688# 0.413585f
C63 minus.n20 a_n1472_n2688# 0.18586f
C64 minus.n21 a_n1472_n2688# 0.345391f
C65 minus.n22 a_n1472_n2688# 1.92904f
C66 drain_left.t9 a_n1472_n2688# 2.33213f
C67 drain_left.t5 a_n1472_n2688# 0.2092f
C68 drain_left.t1 a_n1472_n2688# 0.2092f
C69 drain_left.n0 a_n1472_n2688# 1.8298f
C70 drain_left.n1 a_n1472_n2688# 0.670355f
C71 drain_left.t7 a_n1472_n2688# 0.2092f
C72 drain_left.t3 a_n1472_n2688# 0.2092f
C73 drain_left.n2 a_n1472_n2688# 1.83159f
C74 drain_left.n3 a_n1472_n2688# 1.45674f
C75 drain_left.t8 a_n1472_n2688# 2.33213f
C76 drain_left.t4 a_n1472_n2688# 0.2092f
C77 drain_left.t2 a_n1472_n2688# 0.2092f
C78 drain_left.n4 a_n1472_n2688# 1.82981f
C79 drain_left.n5 a_n1472_n2688# 0.705722f
C80 drain_left.t0 a_n1472_n2688# 0.2092f
C81 drain_left.t6 a_n1472_n2688# 0.2092f
C82 drain_left.n6 a_n1472_n2688# 1.8298f
C83 drain_left.n7 a_n1472_n2688# 0.58341f
C84 source.t12 a_n1472_n2688# 2.34197f
C85 source.n0 a_n1472_n2688# 1.34669f
C86 source.t13 a_n1472_n2688# 0.219625f
C87 source.t15 a_n1472_n2688# 0.219625f
C88 source.n1 a_n1472_n2688# 1.83856f
C89 source.n2 a_n1472_n2688# 0.395895f
C90 source.t18 a_n1472_n2688# 0.219625f
C91 source.t19 a_n1472_n2688# 0.219625f
C92 source.n3 a_n1472_n2688# 1.83856f
C93 source.n4 a_n1472_n2688# 0.415624f
C94 source.t5 a_n1472_n2688# 2.34197f
C95 source.n5 a_n1472_n2688# 0.51119f
C96 source.t1 a_n1472_n2688# 0.219625f
C97 source.t2 a_n1472_n2688# 0.219625f
C98 source.n6 a_n1472_n2688# 1.83856f
C99 source.n7 a_n1472_n2688# 0.395895f
C100 source.t9 a_n1472_n2688# 0.219625f
C101 source.t7 a_n1472_n2688# 0.219625f
C102 source.n8 a_n1472_n2688# 1.83856f
C103 source.n9 a_n1472_n2688# 1.75386f
C104 source.t17 a_n1472_n2688# 0.219625f
C105 source.t14 a_n1472_n2688# 0.219625f
C106 source.n10 a_n1472_n2688# 1.83855f
C107 source.n11 a_n1472_n2688# 1.75386f
C108 source.t16 a_n1472_n2688# 0.219625f
C109 source.t10 a_n1472_n2688# 0.219625f
C110 source.n12 a_n1472_n2688# 1.83855f
C111 source.n13 a_n1472_n2688# 0.3959f
C112 source.t11 a_n1472_n2688# 2.34197f
C113 source.n14 a_n1472_n2688# 0.511195f
C114 source.t8 a_n1472_n2688# 0.219625f
C115 source.t0 a_n1472_n2688# 0.219625f
C116 source.n15 a_n1472_n2688# 1.83855f
C117 source.n16 a_n1472_n2688# 0.41563f
C118 source.t6 a_n1472_n2688# 0.219625f
C119 source.t4 a_n1472_n2688# 0.219625f
C120 source.n17 a_n1472_n2688# 1.83855f
C121 source.n18 a_n1472_n2688# 0.3959f
C122 source.t3 a_n1472_n2688# 2.34197f
C123 source.n19 a_n1472_n2688# 0.658496f
C124 source.n20 a_n1472_n2688# 1.60755f
C125 plus.n0 a_n1472_n2688# 0.054154f
C126 plus.t9 a_n1472_n2688# 0.414318f
C127 plus.t7 a_n1472_n2688# 0.414318f
C128 plus.n1 a_n1472_n2688# 0.022305f
C129 plus.t1 a_n1472_n2688# 0.421998f
C130 plus.t5 a_n1472_n2688# 0.414318f
C131 plus.n2 a_n1472_n2688# 0.173012f
C132 plus.n3 a_n1472_n2688# 0.189716f
C133 plus.n4 a_n1472_n2688# 0.118916f
C134 plus.n5 a_n1472_n2688# 0.054154f
C135 plus.n6 a_n1472_n2688# 0.190977f
C136 plus.n7 a_n1472_n2688# 0.022305f
C137 plus.n8 a_n1472_n2688# 0.173012f
C138 plus.t3 a_n1472_n2688# 0.421998f
C139 plus.n9 a_n1472_n2688# 0.18964f
C140 plus.n10 a_n1472_n2688# 0.530277f
C141 plus.n11 a_n1472_n2688# 0.054154f
C142 plus.t0 a_n1472_n2688# 0.421998f
C143 plus.t4 a_n1472_n2688# 0.414318f
C144 plus.t8 a_n1472_n2688# 0.414318f
C145 plus.n12 a_n1472_n2688# 0.022305f
C146 plus.t2 a_n1472_n2688# 0.414318f
C147 plus.n13 a_n1472_n2688# 0.173012f
C148 plus.t6 a_n1472_n2688# 0.421998f
C149 plus.n14 a_n1472_n2688# 0.189716f
C150 plus.n15 a_n1472_n2688# 0.118916f
C151 plus.n16 a_n1472_n2688# 0.054154f
C152 plus.n17 a_n1472_n2688# 0.190977f
C153 plus.n18 a_n1472_n2688# 0.022305f
C154 plus.n19 a_n1472_n2688# 0.173012f
C155 plus.n20 a_n1472_n2688# 0.18964f
C156 plus.n21 a_n1472_n2688# 1.39599f
.ends

