* NGSPICE file created from diffpair554.ext - technology: sky130A

.subckt diffpair554 minus drain_right drain_left source plus
X0 drain_left.t9 plus.t0 source.t11 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X1 a_n2072_n3888# a_n2072_n3888# a_n2072_n3888# a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.8
X2 drain_right.t9 minus.t0 source.t3 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X3 drain_right.t8 minus.t1 source.t4 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X4 a_n2072_n3888# a_n2072_n3888# a_n2072_n3888# a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X5 a_n2072_n3888# a_n2072_n3888# a_n2072_n3888# a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X6 drain_right.t7 minus.t2 source.t5 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X7 source.t6 minus.t3 drain_right.t6 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X8 source.t10 plus.t1 drain_left.t8 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X9 source.t7 minus.t4 drain_right.t5 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X10 a_n2072_n3888# a_n2072_n3888# a_n2072_n3888# a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X11 source.t17 plus.t2 drain_left.t7 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X12 drain_right.t4 minus.t5 source.t19 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X13 source.t1 minus.t6 drain_right.t3 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X14 source.t18 minus.t7 drain_right.t2 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X15 drain_right.t1 minus.t8 source.t0 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X16 source.t14 plus.t3 drain_left.t6 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X17 drain_left.t5 plus.t4 source.t9 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X18 drain_left.t4 plus.t5 source.t15 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X19 drain_left.t3 plus.t6 source.t8 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X20 source.t12 plus.t7 drain_left.t2 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X21 drain_left.t1 plus.t8 source.t16 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X22 drain_left.t0 plus.t9 source.t13 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X23 drain_right.t0 minus.t9 source.t2 a_n2072_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
R0 plus.n3 plus.t9 524.176
R1 plus.n13 plus.t0 524.176
R2 plus.n8 plus.t6 500.979
R3 plus.n6 plus.t3 500.979
R4 plus.n5 plus.t4 500.979
R5 plus.n4 plus.t7 500.979
R6 plus.n18 plus.t5 500.979
R7 plus.n16 plus.t1 500.979
R8 plus.n15 plus.t8 500.979
R9 plus.n14 plus.t2 500.979
R10 plus.n7 plus.n0 161.3
R11 plus.n9 plus.n8 161.3
R12 plus.n17 plus.n10 161.3
R13 plus.n19 plus.n18 161.3
R14 plus.n5 plus.n2 80.6037
R15 plus.n6 plus.n1 80.6037
R16 plus.n15 plus.n12 80.6037
R17 plus.n16 plus.n11 80.6037
R18 plus.n6 plus.n5 48.2005
R19 plus.n5 plus.n4 48.2005
R20 plus.n16 plus.n15 48.2005
R21 plus.n15 plus.n14 48.2005
R22 plus plus.n19 32.1638
R23 plus.n7 plus.n6 32.1338
R24 plus.n17 plus.n16 32.1338
R25 plus.n3 plus.n2 31.8629
R26 plus.n13 plus.n12 31.8629
R27 plus.n4 plus.n3 16.2333
R28 plus.n14 plus.n13 16.2333
R29 plus.n8 plus.n7 16.0672
R30 plus.n18 plus.n17 16.0672
R31 plus plus.n9 13.4569
R32 plus.n2 plus.n1 0.380177
R33 plus.n12 plus.n11 0.380177
R34 plus.n1 plus.n0 0.285035
R35 plus.n11 plus.n10 0.285035
R36 plus.n9 plus.n0 0.189894
R37 plus.n19 plus.n10 0.189894
R38 source.n5 source.t19 45.521
R39 source.n19 source.t3 45.5208
R40 source.n14 source.t11 45.5208
R41 source.n0 source.t8 45.5208
R42 source.n2 source.n1 44.201
R43 source.n4 source.n3 44.201
R44 source.n7 source.n6 44.201
R45 source.n9 source.n8 44.201
R46 source.n18 source.n17 44.2008
R47 source.n16 source.n15 44.2008
R48 source.n13 source.n12 44.2008
R49 source.n11 source.n10 44.2008
R50 source.n11 source.n9 25.5087
R51 source.n20 source.n0 18.7846
R52 source.n20 source.n19 5.7505
R53 source.n17 source.t2 1.3205
R54 source.n17 source.t6 1.3205
R55 source.n15 source.t4 1.3205
R56 source.n15 source.t1 1.3205
R57 source.n12 source.t16 1.3205
R58 source.n12 source.t17 1.3205
R59 source.n10 source.t15 1.3205
R60 source.n10 source.t10 1.3205
R61 source.n1 source.t9 1.3205
R62 source.n1 source.t14 1.3205
R63 source.n3 source.t13 1.3205
R64 source.n3 source.t12 1.3205
R65 source.n6 source.t5 1.3205
R66 source.n6 source.t7 1.3205
R67 source.n8 source.t0 1.3205
R68 source.n8 source.t18 1.3205
R69 source.n9 source.n7 0.974638
R70 source.n7 source.n5 0.974638
R71 source.n4 source.n2 0.974638
R72 source.n2 source.n0 0.974638
R73 source.n13 source.n11 0.974638
R74 source.n14 source.n13 0.974638
R75 source.n18 source.n16 0.974638
R76 source.n19 source.n18 0.974638
R77 source.n5 source.n4 0.957397
R78 source.n16 source.n14 0.957397
R79 source source.n20 0.188
R80 drain_left.n5 drain_left.t0 63.1739
R81 drain_left.n1 drain_left.t4 63.1737
R82 drain_left.n3 drain_left.n2 61.5548
R83 drain_left.n5 drain_left.n4 60.8798
R84 drain_left.n7 drain_left.n6 60.8796
R85 drain_left.n1 drain_left.n0 60.8796
R86 drain_left drain_left.n3 33.7799
R87 drain_left drain_left.n7 6.62735
R88 drain_left.n2 drain_left.t7 1.3205
R89 drain_left.n2 drain_left.t9 1.3205
R90 drain_left.n0 drain_left.t8 1.3205
R91 drain_left.n0 drain_left.t1 1.3205
R92 drain_left.n6 drain_left.t6 1.3205
R93 drain_left.n6 drain_left.t3 1.3205
R94 drain_left.n4 drain_left.t2 1.3205
R95 drain_left.n4 drain_left.t5 1.3205
R96 drain_left.n7 drain_left.n5 0.974638
R97 drain_left.n3 drain_left.n1 0.188688
R98 minus.n3 minus.t5 524.176
R99 minus.n13 minus.t1 524.176
R100 minus.n2 minus.t4 500.979
R101 minus.n1 minus.t2 500.979
R102 minus.n6 minus.t7 500.979
R103 minus.n8 minus.t8 500.979
R104 minus.n12 minus.t6 500.979
R105 minus.n11 minus.t9 500.979
R106 minus.n16 minus.t3 500.979
R107 minus.n18 minus.t0 500.979
R108 minus.n9 minus.n8 161.3
R109 minus.n7 minus.n0 161.3
R110 minus.n19 minus.n18 161.3
R111 minus.n17 minus.n10 161.3
R112 minus.n6 minus.n5 80.6037
R113 minus.n4 minus.n1 80.6037
R114 minus.n16 minus.n15 80.6037
R115 minus.n14 minus.n11 80.6037
R116 minus.n2 minus.n1 48.2005
R117 minus.n6 minus.n1 48.2005
R118 minus.n12 minus.n11 48.2005
R119 minus.n16 minus.n11 48.2005
R120 minus.n20 minus.n9 39.4191
R121 minus.n7 minus.n6 32.1338
R122 minus.n17 minus.n16 32.1338
R123 minus.n4 minus.n3 31.8629
R124 minus.n14 minus.n13 31.8629
R125 minus.n3 minus.n2 16.2333
R126 minus.n13 minus.n12 16.2333
R127 minus.n8 minus.n7 16.0672
R128 minus.n18 minus.n17 16.0672
R129 minus.n20 minus.n19 6.67664
R130 minus.n5 minus.n4 0.380177
R131 minus.n15 minus.n14 0.380177
R132 minus.n5 minus.n0 0.285035
R133 minus.n15 minus.n10 0.285035
R134 minus.n9 minus.n0 0.189894
R135 minus.n19 minus.n10 0.189894
R136 minus minus.n20 0.188
R137 drain_right.n1 drain_right.t8 63.1737
R138 drain_right.n7 drain_right.t1 62.1998
R139 drain_right.n6 drain_right.n4 61.8538
R140 drain_right.n3 drain_right.n2 61.5548
R141 drain_right.n6 drain_right.n5 60.8798
R142 drain_right.n1 drain_right.n0 60.8796
R143 drain_right drain_right.n3 33.2267
R144 drain_right drain_right.n7 6.14028
R145 drain_right.n2 drain_right.t6 1.3205
R146 drain_right.n2 drain_right.t9 1.3205
R147 drain_right.n0 drain_right.t3 1.3205
R148 drain_right.n0 drain_right.t0 1.3205
R149 drain_right.n4 drain_right.t5 1.3205
R150 drain_right.n4 drain_right.t4 1.3205
R151 drain_right.n5 drain_right.t2 1.3205
R152 drain_right.n5 drain_right.t7 1.3205
R153 drain_right.n7 drain_right.n6 0.974638
R154 drain_right.n3 drain_right.n1 0.188688
C0 plus minus 6.27997f
C1 plus source 8.64156f
C2 drain_left minus 0.172418f
C3 drain_right minus 8.86352f
C4 drain_left source 16.3041f
C5 drain_right source 16.2967f
C6 drain_left plus 9.063499f
C7 drain_right plus 0.360609f
C8 drain_left drain_right 1.03481f
C9 minus source 8.626941f
C10 drain_right a_n2072_n3888# 7.86728f
C11 drain_left a_n2072_n3888# 8.17925f
C12 source a_n2072_n3888# 7.742919f
C13 minus a_n2072_n3888# 8.318291f
C14 plus a_n2072_n3888# 10.09949f
C15 drain_right.t8 a_n2072_n3888# 3.26115f
C16 drain_right.t3 a_n2072_n3888# 0.282194f
C17 drain_right.t0 a_n2072_n3888# 0.282194f
C18 drain_right.n0 a_n2072_n3888# 2.5507f
C19 drain_right.n1 a_n2072_n3888# 0.625573f
C20 drain_right.t6 a_n2072_n3888# 0.282194f
C21 drain_right.t9 a_n2072_n3888# 0.282194f
C22 drain_right.n2 a_n2072_n3888# 2.55434f
C23 drain_right.n3 a_n2072_n3888# 1.69669f
C24 drain_right.t5 a_n2072_n3888# 0.282194f
C25 drain_right.t4 a_n2072_n3888# 0.282194f
C26 drain_right.n4 a_n2072_n3888# 2.55627f
C27 drain_right.t2 a_n2072_n3888# 0.282194f
C28 drain_right.t7 a_n2072_n3888# 0.282194f
C29 drain_right.n5 a_n2072_n3888# 2.55071f
C30 drain_right.n6 a_n2072_n3888# 0.692913f
C31 drain_right.t1 a_n2072_n3888# 3.25585f
C32 drain_right.n7 a_n2072_n3888# 0.567568f
C33 minus.n0 a_n2072_n3888# 0.05393f
C34 minus.t2 a_n2072_n3888# 1.3782f
C35 minus.n1 a_n2072_n3888# 0.540568f
C36 minus.t7 a_n2072_n3888# 1.3782f
C37 minus.t5 a_n2072_n3888# 1.40171f
C38 minus.t4 a_n2072_n3888# 1.3782f
C39 minus.n2 a_n2072_n3888# 0.53959f
C40 minus.n3 a_n2072_n3888# 0.512267f
C41 minus.n4 a_n2072_n3888# 0.24802f
C42 minus.n5 a_n2072_n3888# 0.067318f
C43 minus.n6 a_n2072_n3888# 0.537827f
C44 minus.n7 a_n2072_n3888# 0.009171f
C45 minus.t8 a_n2072_n3888# 1.3782f
C46 minus.n8 a_n2072_n3888# 0.525915f
C47 minus.n9 a_n2072_n3888# 1.63349f
C48 minus.n10 a_n2072_n3888# 0.05393f
C49 minus.t9 a_n2072_n3888# 1.3782f
C50 minus.n11 a_n2072_n3888# 0.540568f
C51 minus.t1 a_n2072_n3888# 1.40171f
C52 minus.t6 a_n2072_n3888# 1.3782f
C53 minus.n12 a_n2072_n3888# 0.53959f
C54 minus.n13 a_n2072_n3888# 0.512267f
C55 minus.n14 a_n2072_n3888# 0.24802f
C56 minus.n15 a_n2072_n3888# 0.067318f
C57 minus.t3 a_n2072_n3888# 1.3782f
C58 minus.n16 a_n2072_n3888# 0.537827f
C59 minus.n17 a_n2072_n3888# 0.009171f
C60 minus.t0 a_n2072_n3888# 1.3782f
C61 minus.n18 a_n2072_n3888# 0.525915f
C62 minus.n19 a_n2072_n3888# 0.280911f
C63 minus.n20 a_n2072_n3888# 1.96079f
C64 drain_left.t4 a_n2072_n3888# 3.27493f
C65 drain_left.t8 a_n2072_n3888# 0.283386f
C66 drain_left.t1 a_n2072_n3888# 0.283386f
C67 drain_left.n0 a_n2072_n3888# 2.56148f
C68 drain_left.n1 a_n2072_n3888# 0.628216f
C69 drain_left.t7 a_n2072_n3888# 0.283386f
C70 drain_left.t9 a_n2072_n3888# 0.283386f
C71 drain_left.n2 a_n2072_n3888# 2.56514f
C72 drain_left.n3 a_n2072_n3888# 1.75345f
C73 drain_left.t0 a_n2072_n3888# 3.27493f
C74 drain_left.t2 a_n2072_n3888# 0.283386f
C75 drain_left.t5 a_n2072_n3888# 0.283386f
C76 drain_left.n4 a_n2072_n3888# 2.56148f
C77 drain_left.n5 a_n2072_n3888# 0.685813f
C78 drain_left.t6 a_n2072_n3888# 0.283386f
C79 drain_left.t3 a_n2072_n3888# 0.283386f
C80 drain_left.n6 a_n2072_n3888# 2.56148f
C81 drain_left.n7 a_n2072_n3888# 0.560287f
C82 source.t8 a_n2072_n3888# 3.28272f
C83 source.n0 a_n2072_n3888# 1.57581f
C84 source.t9 a_n2072_n3888# 0.292927f
C85 source.t14 a_n2072_n3888# 0.292927f
C86 source.n1 a_n2072_n3888# 2.57312f
C87 source.n2 a_n2072_n3888# 0.398559f
C88 source.t13 a_n2072_n3888# 0.292927f
C89 source.t12 a_n2072_n3888# 0.292927f
C90 source.n3 a_n2072_n3888# 2.57312f
C91 source.n4 a_n2072_n3888# 0.397186f
C92 source.t19 a_n2072_n3888# 3.28272f
C93 source.n5 a_n2072_n3888# 0.486473f
C94 source.t5 a_n2072_n3888# 0.292927f
C95 source.t7 a_n2072_n3888# 0.292927f
C96 source.n6 a_n2072_n3888# 2.57312f
C97 source.n7 a_n2072_n3888# 0.398559f
C98 source.t0 a_n2072_n3888# 0.292927f
C99 source.t18 a_n2072_n3888# 0.292927f
C100 source.n8 a_n2072_n3888# 2.57312f
C101 source.n9 a_n2072_n3888# 1.98828f
C102 source.t15 a_n2072_n3888# 0.292927f
C103 source.t10 a_n2072_n3888# 0.292927f
C104 source.n10 a_n2072_n3888# 2.57312f
C105 source.n11 a_n2072_n3888# 1.98829f
C106 source.t16 a_n2072_n3888# 0.292927f
C107 source.t17 a_n2072_n3888# 0.292927f
C108 source.n12 a_n2072_n3888# 2.57312f
C109 source.n13 a_n2072_n3888# 0.398562f
C110 source.t11 a_n2072_n3888# 3.28272f
C111 source.n14 a_n2072_n3888# 0.486477f
C112 source.t4 a_n2072_n3888# 0.292927f
C113 source.t1 a_n2072_n3888# 0.292927f
C114 source.n15 a_n2072_n3888# 2.57312f
C115 source.n16 a_n2072_n3888# 0.397189f
C116 source.t2 a_n2072_n3888# 0.292927f
C117 source.t6 a_n2072_n3888# 0.292927f
C118 source.n17 a_n2072_n3888# 2.57312f
C119 source.n18 a_n2072_n3888# 0.398562f
C120 source.t3 a_n2072_n3888# 3.28272f
C121 source.n19 a_n2072_n3888# 0.614242f
C122 source.n20 a_n2072_n3888# 1.82754f
C123 plus.n0 a_n2072_n3888# 0.054571f
C124 plus.t6 a_n2072_n3888# 1.39457f
C125 plus.t3 a_n2072_n3888# 1.39457f
C126 plus.n1 a_n2072_n3888# 0.068118f
C127 plus.t4 a_n2072_n3888# 1.39457f
C128 plus.n2 a_n2072_n3888# 0.250966f
C129 plus.t7 a_n2072_n3888# 1.39457f
C130 plus.t9 a_n2072_n3888# 1.41836f
C131 plus.n3 a_n2072_n3888# 0.518351f
C132 plus.n4 a_n2072_n3888# 0.546f
C133 plus.n5 a_n2072_n3888# 0.546989f
C134 plus.n6 a_n2072_n3888# 0.544215f
C135 plus.n7 a_n2072_n3888# 0.00928f
C136 plus.n8 a_n2072_n3888# 0.532162f
C137 plus.n9 a_n2072_n3888# 0.533746f
C138 plus.n10 a_n2072_n3888# 0.054571f
C139 plus.t5 a_n2072_n3888# 1.39457f
C140 plus.n11 a_n2072_n3888# 0.068118f
C141 plus.t1 a_n2072_n3888# 1.39457f
C142 plus.n12 a_n2072_n3888# 0.250966f
C143 plus.t8 a_n2072_n3888# 1.39457f
C144 plus.t0 a_n2072_n3888# 1.41836f
C145 plus.n13 a_n2072_n3888# 0.518351f
C146 plus.t2 a_n2072_n3888# 1.39457f
C147 plus.n14 a_n2072_n3888# 0.546f
C148 plus.n15 a_n2072_n3888# 0.546989f
C149 plus.n16 a_n2072_n3888# 0.544215f
C150 plus.n17 a_n2072_n3888# 0.00928f
C151 plus.n18 a_n2072_n3888# 0.532162f
C152 plus.n19 a_n2072_n3888# 1.36614f
.ends

