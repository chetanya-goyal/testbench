* NGSPICE file created from diffpair625.ext - technology: sky130A

.subckt diffpair625 minus drain_right drain_left source plus
X0 drain_left.t11 plus.t0 source.t14 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X1 source.t2 minus.t0 drain_right.t11 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X2 source.t15 plus.t1 drain_left.t10 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X3 drain_right.t10 minus.t1 source.t7 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X4 source.t16 plus.t2 drain_left.t9 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X5 source.t1 minus.t2 drain_right.t9 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X6 a_n2158_n4888# a_n2158_n4888# a_n2158_n4888# a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.7
X7 source.t5 minus.t3 drain_right.t8 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X8 source.t20 plus.t3 drain_left.t8 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X9 source.t11 plus.t4 drain_left.t7 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X10 source.t13 plus.t5 drain_left.t6 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X11 drain_right.t7 minus.t4 source.t6 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X12 source.t22 minus.t5 drain_right.t6 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X13 drain_right.t5 minus.t6 source.t8 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X14 drain_right.t4 minus.t7 source.t0 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X15 drain_left.t5 plus.t6 source.t10 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X16 drain_left.t4 plus.t7 source.t12 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X17 source.t9 plus.t8 drain_left.t3 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X18 drain_left.t2 plus.t9 source.t19 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X19 a_n2158_n4888# a_n2158_n4888# a_n2158_n4888# a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X20 drain_right.t3 minus.t8 source.t23 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X21 drain_left.t1 plus.t10 source.t18 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X22 drain_left.t0 plus.t11 source.t17 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X23 a_n2158_n4888# a_n2158_n4888# a_n2158_n4888# a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X24 drain_right.t2 minus.t9 source.t4 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X25 source.t3 minus.t10 drain_right.t1 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X26 source.t21 minus.t11 drain_right.t0 a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X27 a_n2158_n4888# a_n2158_n4888# a_n2158_n4888# a_n2158_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
R0 plus.n5 plus.t4 767.995
R1 plus.n23 plus.t0 767.995
R2 plus.n16 plus.t7 744.691
R3 plus.n14 plus.t3 744.691
R4 plus.n2 plus.t6 744.691
R5 plus.n8 plus.t2 744.691
R6 plus.n4 plus.t10 744.691
R7 plus.n34 plus.t5 744.691
R8 plus.n32 plus.t9 744.691
R9 plus.n20 plus.t8 744.691
R10 plus.n26 plus.t11 744.691
R11 plus.n22 plus.t1 744.691
R12 plus.n7 plus.n6 161.3
R13 plus.n8 plus.n3 161.3
R14 plus.n10 plus.n9 161.3
R15 plus.n11 plus.n2 161.3
R16 plus.n13 plus.n12 161.3
R17 plus.n14 plus.n1 161.3
R18 plus.n15 plus.n0 161.3
R19 plus.n17 plus.n16 161.3
R20 plus.n25 plus.n24 161.3
R21 plus.n26 plus.n21 161.3
R22 plus.n28 plus.n27 161.3
R23 plus.n29 plus.n20 161.3
R24 plus.n31 plus.n30 161.3
R25 plus.n32 plus.n19 161.3
R26 plus.n33 plus.n18 161.3
R27 plus.n35 plus.n34 161.3
R28 plus.n6 plus.n5 44.8907
R29 plus.n24 plus.n23 44.8907
R30 plus plus.n35 34.3513
R31 plus.n16 plus.n15 32.8641
R32 plus.n34 plus.n33 32.8641
R33 plus.n14 plus.n13 28.4823
R34 plus.n7 plus.n4 28.4823
R35 plus.n32 plus.n31 28.4823
R36 plus.n25 plus.n22 28.4823
R37 plus.n9 plus.n8 24.1005
R38 plus.n9 plus.n2 24.1005
R39 plus.n27 plus.n20 24.1005
R40 plus.n27 plus.n26 24.1005
R41 plus.n13 plus.n2 19.7187
R42 plus.n8 plus.n7 19.7187
R43 plus.n31 plus.n20 19.7187
R44 plus.n26 plus.n25 19.7187
R45 plus.n5 plus.n4 18.4104
R46 plus.n23 plus.n22 18.4104
R47 plus.n15 plus.n14 15.3369
R48 plus.n33 plus.n32 15.3369
R49 plus plus.n17 15.3187
R50 plus.n6 plus.n3 0.189894
R51 plus.n10 plus.n3 0.189894
R52 plus.n11 plus.n10 0.189894
R53 plus.n12 plus.n11 0.189894
R54 plus.n12 plus.n1 0.189894
R55 plus.n1 plus.n0 0.189894
R56 plus.n17 plus.n0 0.189894
R57 plus.n35 plus.n18 0.189894
R58 plus.n19 plus.n18 0.189894
R59 plus.n30 plus.n19 0.189894
R60 plus.n30 plus.n29 0.189894
R61 plus.n29 plus.n28 0.189894
R62 plus.n28 plus.n21 0.189894
R63 plus.n24 plus.n21 0.189894
R64 source.n0 source.t12 44.1297
R65 source.n5 source.t11 44.1296
R66 source.n6 source.t23 44.1296
R67 source.n11 source.t21 44.1296
R68 source.n23 source.t4 44.1295
R69 source.n18 source.t22 44.1295
R70 source.n17 source.t14 44.1295
R71 source.n12 source.t13 44.1295
R72 source.n2 source.n1 43.1397
R73 source.n4 source.n3 43.1397
R74 source.n8 source.n7 43.1397
R75 source.n10 source.n9 43.1397
R76 source.n22 source.n21 43.1396
R77 source.n20 source.n19 43.1396
R78 source.n16 source.n15 43.1396
R79 source.n14 source.n13 43.1396
R80 source.n12 source.n11 28.2363
R81 source.n24 source.n0 22.5294
R82 source.n24 source.n23 5.7074
R83 source.n21 source.t7 0.9905
R84 source.n21 source.t5 0.9905
R85 source.n19 source.t6 0.9905
R86 source.n19 source.t2 0.9905
R87 source.n15 source.t17 0.9905
R88 source.n15 source.t15 0.9905
R89 source.n13 source.t19 0.9905
R90 source.n13 source.t9 0.9905
R91 source.n1 source.t10 0.9905
R92 source.n1 source.t20 0.9905
R93 source.n3 source.t18 0.9905
R94 source.n3 source.t16 0.9905
R95 source.n7 source.t0 0.9905
R96 source.n7 source.t1 0.9905
R97 source.n9 source.t8 0.9905
R98 source.n9 source.t3 0.9905
R99 source.n11 source.n10 0.888431
R100 source.n10 source.n8 0.888431
R101 source.n8 source.n6 0.888431
R102 source.n5 source.n4 0.888431
R103 source.n4 source.n2 0.888431
R104 source.n2 source.n0 0.888431
R105 source.n14 source.n12 0.888431
R106 source.n16 source.n14 0.888431
R107 source.n17 source.n16 0.888431
R108 source.n20 source.n18 0.888431
R109 source.n22 source.n20 0.888431
R110 source.n23 source.n22 0.888431
R111 source.n6 source.n5 0.470328
R112 source.n18 source.n17 0.470328
R113 source source.n24 0.188
R114 drain_left.n6 drain_left.n4 60.7064
R115 drain_left.n3 drain_left.n2 60.651
R116 drain_left.n3 drain_left.n0 60.651
R117 drain_left.n8 drain_left.n7 59.8185
R118 drain_left.n6 drain_left.n5 59.8185
R119 drain_left.n3 drain_left.n1 59.8184
R120 drain_left drain_left.n3 37.8673
R121 drain_left drain_left.n8 6.54115
R122 drain_left.n1 drain_left.t3 0.9905
R123 drain_left.n1 drain_left.t0 0.9905
R124 drain_left.n2 drain_left.t10 0.9905
R125 drain_left.n2 drain_left.t11 0.9905
R126 drain_left.n0 drain_left.t6 0.9905
R127 drain_left.n0 drain_left.t2 0.9905
R128 drain_left.n7 drain_left.t8 0.9905
R129 drain_left.n7 drain_left.t4 0.9905
R130 drain_left.n5 drain_left.t9 0.9905
R131 drain_left.n5 drain_left.t5 0.9905
R132 drain_left.n4 drain_left.t7 0.9905
R133 drain_left.n4 drain_left.t1 0.9905
R134 drain_left.n8 drain_left.n6 0.888431
R135 minus.n5 minus.t8 767.995
R136 minus.n23 minus.t5 767.995
R137 minus.n4 minus.t2 744.691
R138 minus.n8 minus.t7 744.691
R139 minus.n10 minus.t10 744.691
R140 minus.n14 minus.t6 744.691
R141 minus.n16 minus.t11 744.691
R142 minus.n22 minus.t4 744.691
R143 minus.n26 minus.t0 744.691
R144 minus.n28 minus.t1 744.691
R145 minus.n32 minus.t3 744.691
R146 minus.n34 minus.t9 744.691
R147 minus.n17 minus.n16 161.3
R148 minus.n15 minus.n0 161.3
R149 minus.n14 minus.n13 161.3
R150 minus.n12 minus.n1 161.3
R151 minus.n11 minus.n10 161.3
R152 minus.n9 minus.n2 161.3
R153 minus.n8 minus.n7 161.3
R154 minus.n6 minus.n3 161.3
R155 minus.n35 minus.n34 161.3
R156 minus.n33 minus.n18 161.3
R157 minus.n32 minus.n31 161.3
R158 minus.n30 minus.n19 161.3
R159 minus.n29 minus.n28 161.3
R160 minus.n27 minus.n20 161.3
R161 minus.n26 minus.n25 161.3
R162 minus.n24 minus.n21 161.3
R163 minus.n6 minus.n5 44.8907
R164 minus.n24 minus.n23 44.8907
R165 minus.n36 minus.n17 43.5005
R166 minus.n16 minus.n15 32.8641
R167 minus.n34 minus.n33 32.8641
R168 minus.n4 minus.n3 28.4823
R169 minus.n14 minus.n1 28.4823
R170 minus.n22 minus.n21 28.4823
R171 minus.n32 minus.n19 28.4823
R172 minus.n10 minus.n9 24.1005
R173 minus.n9 minus.n8 24.1005
R174 minus.n27 minus.n26 24.1005
R175 minus.n28 minus.n27 24.1005
R176 minus.n8 minus.n3 19.7187
R177 minus.n10 minus.n1 19.7187
R178 minus.n26 minus.n21 19.7187
R179 minus.n28 minus.n19 19.7187
R180 minus.n5 minus.n4 18.4104
R181 minus.n23 minus.n22 18.4104
R182 minus.n15 minus.n14 15.3369
R183 minus.n33 minus.n32 15.3369
R184 minus.n36 minus.n35 6.64444
R185 minus.n17 minus.n0 0.189894
R186 minus.n13 minus.n0 0.189894
R187 minus.n13 minus.n12 0.189894
R188 minus.n12 minus.n11 0.189894
R189 minus.n11 minus.n2 0.189894
R190 minus.n7 minus.n2 0.189894
R191 minus.n7 minus.n6 0.189894
R192 minus.n25 minus.n24 0.189894
R193 minus.n25 minus.n20 0.189894
R194 minus.n29 minus.n20 0.189894
R195 minus.n30 minus.n29 0.189894
R196 minus.n31 minus.n30 0.189894
R197 minus.n31 minus.n18 0.189894
R198 minus.n35 minus.n18 0.189894
R199 minus minus.n36 0.188
R200 drain_right.n6 drain_right.n4 60.7064
R201 drain_right.n3 drain_right.n2 60.651
R202 drain_right.n3 drain_right.n0 60.651
R203 drain_right.n6 drain_right.n5 59.8185
R204 drain_right.n8 drain_right.n7 59.8185
R205 drain_right.n3 drain_right.n1 59.8184
R206 drain_right drain_right.n3 37.3141
R207 drain_right drain_right.n8 6.54115
R208 drain_right.n1 drain_right.t11 0.9905
R209 drain_right.n1 drain_right.t10 0.9905
R210 drain_right.n2 drain_right.t8 0.9905
R211 drain_right.n2 drain_right.t2 0.9905
R212 drain_right.n0 drain_right.t6 0.9905
R213 drain_right.n0 drain_right.t7 0.9905
R214 drain_right.n4 drain_right.t9 0.9905
R215 drain_right.n4 drain_right.t3 0.9905
R216 drain_right.n5 drain_right.t1 0.9905
R217 drain_right.n5 drain_right.t4 0.9905
R218 drain_right.n7 drain_right.t0 0.9905
R219 drain_right.n7 drain_right.t5 0.9905
R220 drain_right.n8 drain_right.n6 0.888431
C0 drain_right plus 0.366822f
C1 minus drain_right 12.8186f
C2 source drain_left 23.9667f
C3 source drain_right 23.9687f
C4 minus plus 7.31627f
C5 drain_left drain_right 1.08491f
C6 source plus 12.4143f
C7 drain_left plus 13.0303f
C8 minus source 12.4003f
C9 minus drain_left 0.17184f
C10 drain_right a_n2158_n4888# 7.68712f
C11 drain_left a_n2158_n4888# 7.99557f
C12 source a_n2158_n4888# 13.60714f
C13 minus a_n2158_n4888# 9.048603f
C14 plus a_n2158_n4888# 11.156811f
C15 drain_right.t6 a_n2158_n4888# 0.430672f
C16 drain_right.t7 a_n2158_n4888# 0.430672f
C17 drain_right.n0 a_n2158_n4888# 3.94269f
C18 drain_right.t11 a_n2158_n4888# 0.430672f
C19 drain_right.t10 a_n2158_n4888# 0.430672f
C20 drain_right.n1 a_n2158_n4888# 3.9373f
C21 drain_right.t8 a_n2158_n4888# 0.430672f
C22 drain_right.t2 a_n2158_n4888# 0.430672f
C23 drain_right.n2 a_n2158_n4888# 3.94269f
C24 drain_right.n3 a_n2158_n4888# 3.01154f
C25 drain_right.t9 a_n2158_n4888# 0.430672f
C26 drain_right.t3 a_n2158_n4888# 0.430672f
C27 drain_right.n4 a_n2158_n4888# 3.9431f
C28 drain_right.t1 a_n2158_n4888# 0.430672f
C29 drain_right.t4 a_n2158_n4888# 0.430672f
C30 drain_right.n5 a_n2158_n4888# 3.93729f
C31 drain_right.n6 a_n2158_n4888# 0.776939f
C32 drain_right.t0 a_n2158_n4888# 0.430672f
C33 drain_right.t5 a_n2158_n4888# 0.430672f
C34 drain_right.n7 a_n2158_n4888# 3.93729f
C35 drain_right.n8 a_n2158_n4888# 0.62691f
C36 minus.n0 a_n2158_n4888# 0.04138f
C37 minus.n1 a_n2158_n4888# 0.00939f
C38 minus.t6 a_n2158_n4888# 1.64057f
C39 minus.n2 a_n2158_n4888# 0.04138f
C40 minus.n3 a_n2158_n4888# 0.00939f
C41 minus.t7 a_n2158_n4888# 1.64057f
C42 minus.t8 a_n2158_n4888# 1.65913f
C43 minus.t2 a_n2158_n4888# 1.64057f
C44 minus.n4 a_n2158_n4888# 0.616392f
C45 minus.n5 a_n2158_n4888# 0.596907f
C46 minus.n6 a_n2158_n4888# 0.173594f
C47 minus.n7 a_n2158_n4888# 0.04138f
C48 minus.n8 a_n2158_n4888# 0.611764f
C49 minus.n9 a_n2158_n4888# 0.00939f
C50 minus.t10 a_n2158_n4888# 1.64057f
C51 minus.n10 a_n2158_n4888# 0.611764f
C52 minus.n11 a_n2158_n4888# 0.04138f
C53 minus.n12 a_n2158_n4888# 0.04138f
C54 minus.n13 a_n2158_n4888# 0.04138f
C55 minus.n14 a_n2158_n4888# 0.611764f
C56 minus.n15 a_n2158_n4888# 0.00939f
C57 minus.t11 a_n2158_n4888# 1.64057f
C58 minus.n16 a_n2158_n4888# 0.609851f
C59 minus.n17 a_n2158_n4888# 1.93298f
C60 minus.n18 a_n2158_n4888# 0.04138f
C61 minus.n19 a_n2158_n4888# 0.00939f
C62 minus.n20 a_n2158_n4888# 0.04138f
C63 minus.n21 a_n2158_n4888# 0.00939f
C64 minus.t5 a_n2158_n4888# 1.65913f
C65 minus.t4 a_n2158_n4888# 1.64057f
C66 minus.n22 a_n2158_n4888# 0.616392f
C67 minus.n23 a_n2158_n4888# 0.596907f
C68 minus.n24 a_n2158_n4888# 0.173594f
C69 minus.n25 a_n2158_n4888# 0.04138f
C70 minus.t0 a_n2158_n4888# 1.64057f
C71 minus.n26 a_n2158_n4888# 0.611764f
C72 minus.n27 a_n2158_n4888# 0.00939f
C73 minus.t1 a_n2158_n4888# 1.64057f
C74 minus.n28 a_n2158_n4888# 0.611764f
C75 minus.n29 a_n2158_n4888# 0.04138f
C76 minus.n30 a_n2158_n4888# 0.04138f
C77 minus.n31 a_n2158_n4888# 0.04138f
C78 minus.t3 a_n2158_n4888# 1.64057f
C79 minus.n32 a_n2158_n4888# 0.611764f
C80 minus.n33 a_n2158_n4888# 0.00939f
C81 minus.t9 a_n2158_n4888# 1.64057f
C82 minus.n34 a_n2158_n4888# 0.609851f
C83 minus.n35 a_n2158_n4888# 0.284518f
C84 minus.n36 a_n2158_n4888# 2.29558f
C85 drain_left.t6 a_n2158_n4888# 0.431762f
C86 drain_left.t2 a_n2158_n4888# 0.431762f
C87 drain_left.n0 a_n2158_n4888# 3.95267f
C88 drain_left.t3 a_n2158_n4888# 0.431762f
C89 drain_left.t0 a_n2158_n4888# 0.431762f
C90 drain_left.n1 a_n2158_n4888# 3.94726f
C91 drain_left.t10 a_n2158_n4888# 0.431762f
C92 drain_left.t11 a_n2158_n4888# 0.431762f
C93 drain_left.n2 a_n2158_n4888# 3.95267f
C94 drain_left.n3 a_n2158_n4888# 3.07578f
C95 drain_left.t7 a_n2158_n4888# 0.431762f
C96 drain_left.t1 a_n2158_n4888# 0.431762f
C97 drain_left.n4 a_n2158_n4888# 3.95308f
C98 drain_left.t9 a_n2158_n4888# 0.431762f
C99 drain_left.t5 a_n2158_n4888# 0.431762f
C100 drain_left.n5 a_n2158_n4888# 3.94726f
C101 drain_left.n6 a_n2158_n4888# 0.778905f
C102 drain_left.t8 a_n2158_n4888# 0.431762f
C103 drain_left.t4 a_n2158_n4888# 0.431762f
C104 drain_left.n7 a_n2158_n4888# 3.94726f
C105 drain_left.n8 a_n2158_n4888# 0.628496f
C106 source.t12 a_n2158_n4888# 3.84554f
C107 source.n0 a_n2158_n4888# 1.67292f
C108 source.t10 a_n2158_n4888# 0.336491f
C109 source.t20 a_n2158_n4888# 0.336491f
C110 source.n1 a_n2158_n4888# 3.00837f
C111 source.n2 a_n2158_n4888# 0.340456f
C112 source.t18 a_n2158_n4888# 0.336491f
C113 source.t16 a_n2158_n4888# 0.336491f
C114 source.n3 a_n2158_n4888# 3.00837f
C115 source.n4 a_n2158_n4888# 0.340456f
C116 source.t11 a_n2158_n4888# 3.84555f
C117 source.n5 a_n2158_n4888# 0.392293f
C118 source.t23 a_n2158_n4888# 3.84555f
C119 source.n6 a_n2158_n4888# 0.392293f
C120 source.t0 a_n2158_n4888# 0.336491f
C121 source.t1 a_n2158_n4888# 0.336491f
C122 source.n7 a_n2158_n4888# 3.00837f
C123 source.n8 a_n2158_n4888# 0.340456f
C124 source.t8 a_n2158_n4888# 0.336491f
C125 source.t3 a_n2158_n4888# 0.336491f
C126 source.n9 a_n2158_n4888# 3.00837f
C127 source.n10 a_n2158_n4888# 0.340456f
C128 source.t21 a_n2158_n4888# 3.84555f
C129 source.n11 a_n2158_n4888# 2.06025f
C130 source.t13 a_n2158_n4888# 3.84553f
C131 source.n12 a_n2158_n4888# 2.06027f
C132 source.t19 a_n2158_n4888# 0.336491f
C133 source.t9 a_n2158_n4888# 0.336491f
C134 source.n13 a_n2158_n4888# 3.00838f
C135 source.n14 a_n2158_n4888# 0.34045f
C136 source.t17 a_n2158_n4888# 0.336491f
C137 source.t15 a_n2158_n4888# 0.336491f
C138 source.n15 a_n2158_n4888# 3.00838f
C139 source.n16 a_n2158_n4888# 0.34045f
C140 source.t14 a_n2158_n4888# 3.84553f
C141 source.n17 a_n2158_n4888# 0.392315f
C142 source.t22 a_n2158_n4888# 3.84553f
C143 source.n18 a_n2158_n4888# 0.392315f
C144 source.t6 a_n2158_n4888# 0.336491f
C145 source.t2 a_n2158_n4888# 0.336491f
C146 source.n19 a_n2158_n4888# 3.00838f
C147 source.n20 a_n2158_n4888# 0.34045f
C148 source.t7 a_n2158_n4888# 0.336491f
C149 source.t5 a_n2158_n4888# 0.336491f
C150 source.n21 a_n2158_n4888# 3.00838f
C151 source.n22 a_n2158_n4888# 0.34045f
C152 source.t4 a_n2158_n4888# 3.84553f
C153 source.n23 a_n2158_n4888# 0.531194f
C154 source.n24 a_n2158_n4888# 1.93155f
C155 plus.n0 a_n2158_n4888# 0.041742f
C156 plus.t7 a_n2158_n4888# 1.65493f
C157 plus.t3 a_n2158_n4888# 1.65493f
C158 plus.n1 a_n2158_n4888# 0.041742f
C159 plus.t6 a_n2158_n4888# 1.65493f
C160 plus.n2 a_n2158_n4888# 0.617118f
C161 plus.n3 a_n2158_n4888# 0.041742f
C162 plus.t2 a_n2158_n4888# 1.65493f
C163 plus.t10 a_n2158_n4888# 1.65493f
C164 plus.n4 a_n2158_n4888# 0.621787f
C165 plus.t4 a_n2158_n4888# 1.67365f
C166 plus.n5 a_n2158_n4888# 0.60213f
C167 plus.n6 a_n2158_n4888# 0.175113f
C168 plus.n7 a_n2158_n4888# 0.009472f
C169 plus.n8 a_n2158_n4888# 0.617118f
C170 plus.n9 a_n2158_n4888# 0.009472f
C171 plus.n10 a_n2158_n4888# 0.041742f
C172 plus.n11 a_n2158_n4888# 0.041742f
C173 plus.n12 a_n2158_n4888# 0.041742f
C174 plus.n13 a_n2158_n4888# 0.009472f
C175 plus.n14 a_n2158_n4888# 0.617118f
C176 plus.n15 a_n2158_n4888# 0.009472f
C177 plus.n16 a_n2158_n4888# 0.615188f
C178 plus.n17 a_n2158_n4888# 0.647656f
C179 plus.n18 a_n2158_n4888# 0.041742f
C180 plus.t5 a_n2158_n4888# 1.65493f
C181 plus.n19 a_n2158_n4888# 0.041742f
C182 plus.t9 a_n2158_n4888# 1.65493f
C183 plus.t8 a_n2158_n4888# 1.65493f
C184 plus.n20 a_n2158_n4888# 0.617118f
C185 plus.n21 a_n2158_n4888# 0.041742f
C186 plus.t11 a_n2158_n4888# 1.65493f
C187 plus.t1 a_n2158_n4888# 1.65493f
C188 plus.n22 a_n2158_n4888# 0.621787f
C189 plus.t0 a_n2158_n4888# 1.67365f
C190 plus.n23 a_n2158_n4888# 0.60213f
C191 plus.n24 a_n2158_n4888# 0.175113f
C192 plus.n25 a_n2158_n4888# 0.009472f
C193 plus.n26 a_n2158_n4888# 0.617118f
C194 plus.n27 a_n2158_n4888# 0.009472f
C195 plus.n28 a_n2158_n4888# 0.041742f
C196 plus.n29 a_n2158_n4888# 0.041742f
C197 plus.n30 a_n2158_n4888# 0.041742f
C198 plus.n31 a_n2158_n4888# 0.009472f
C199 plus.n32 a_n2158_n4888# 0.617118f
C200 plus.n33 a_n2158_n4888# 0.009472f
C201 plus.n34 a_n2158_n4888# 0.615188f
C202 plus.n35 a_n2158_n4888# 1.55206f
.ends

