* NGSPICE file created from diffpair298.ext - technology: sky130A

.subckt diffpair298 minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t36 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X1 source.t32 plus.t1 drain_left.t18 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X2 source.t38 plus.t2 drain_left.t17 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X3 drain_left.t16 plus.t3 source.t21 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X4 source.t0 minus.t0 drain_right.t19 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X5 source.t26 plus.t4 drain_left.t15 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X6 drain_right.t18 minus.t1 source.t1 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X7 drain_left.t14 plus.t5 source.t23 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X8 source.t3 minus.t2 drain_right.t17 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X9 source.t9 minus.t3 drain_right.t16 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X10 drain_right.t15 minus.t4 source.t12 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X11 drain_right.t14 minus.t5 source.t10 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X12 drain_right.t13 minus.t6 source.t19 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X13 source.t5 minus.t7 drain_right.t12 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X14 source.t13 minus.t8 drain_right.t11 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X15 a_n2762_n2088# a_n2762_n2088# a_n2762_n2088# a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.6
X16 drain_left.t13 plus.t6 source.t28 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X17 drain_left.t12 plus.t7 source.t27 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X18 a_n2762_n2088# a_n2762_n2088# a_n2762_n2088# a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.6
X19 source.t22 plus.t8 drain_left.t11 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X20 a_n2762_n2088# a_n2762_n2088# a_n2762_n2088# a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.6
X21 drain_right.t10 minus.t9 source.t16 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X22 source.t35 plus.t9 drain_left.t10 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X23 source.t2 minus.t10 drain_right.t9 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X24 a_n2762_n2088# a_n2762_n2088# a_n2762_n2088# a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.6
X25 drain_right.t8 minus.t11 source.t15 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X26 drain_left.t9 plus.t10 source.t33 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X27 drain_right.t7 minus.t12 source.t4 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X28 source.t39 plus.t11 drain_left.t8 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X29 source.t20 plus.t12 drain_left.t7 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X30 drain_left.t6 plus.t13 source.t30 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X31 source.t17 minus.t13 drain_right.t6 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X32 source.t29 plus.t14 drain_left.t5 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X33 drain_right.t5 minus.t14 source.t8 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X34 drain_right.t4 minus.t15 source.t14 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X35 drain_left.t4 plus.t15 source.t37 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X36 source.t34 plus.t16 drain_left.t3 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X37 drain_left.t2 plus.t17 source.t25 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X38 source.t7 minus.t16 drain_right.t3 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X39 drain_right.t2 minus.t17 source.t11 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X40 source.t31 plus.t18 drain_left.t1 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X41 drain_left.t0 plus.t19 source.t24 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X42 source.t18 minus.t18 drain_right.t1 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X43 source.t6 minus.t19 drain_right.t0 a_n2762_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
R0 plus.n8 plus.t16 333.293
R1 plus.n36 plus.t10 333.293
R2 plus.n26 plus.t0 306.473
R3 plus.n25 plus.t2 306.473
R4 plus.n24 plus.t3 306.473
R5 plus.n2 plus.t4 306.473
R6 plus.n18 plus.t5 306.473
R7 plus.n4 plus.t9 306.473
R8 plus.n12 plus.t13 306.473
R9 plus.n6 plus.t14 306.473
R10 plus.n7 plus.t15 306.473
R11 plus.n54 plus.t8 306.473
R12 plus.n53 plus.t19 306.473
R13 plus.n52 plus.t12 306.473
R14 plus.n30 plus.t7 306.473
R15 plus.n46 plus.t18 306.473
R16 plus.n32 plus.t17 306.473
R17 plus.n40 plus.t11 306.473
R18 plus.n34 plus.t6 306.473
R19 plus.n35 plus.t1 306.473
R20 plus.n9 plus.n6 161.3
R21 plus.n11 plus.n10 161.3
R22 plus.n12 plus.n5 161.3
R23 plus.n14 plus.n13 161.3
R24 plus.n15 plus.n4 161.3
R25 plus.n17 plus.n16 161.3
R26 plus.n18 plus.n3 161.3
R27 plus.n20 plus.n19 161.3
R28 plus.n21 plus.n2 161.3
R29 plus.n23 plus.n22 161.3
R30 plus.n24 plus.n1 161.3
R31 plus.n27 plus.n26 161.3
R32 plus.n37 plus.n34 161.3
R33 plus.n39 plus.n38 161.3
R34 plus.n40 plus.n33 161.3
R35 plus.n42 plus.n41 161.3
R36 plus.n43 plus.n32 161.3
R37 plus.n45 plus.n44 161.3
R38 plus.n46 plus.n31 161.3
R39 plus.n48 plus.n47 161.3
R40 plus.n49 plus.n30 161.3
R41 plus.n51 plus.n50 161.3
R42 plus.n52 plus.n29 161.3
R43 plus.n55 plus.n54 161.3
R44 plus.n25 plus.n0 80.6037
R45 plus.n53 plus.n28 80.6037
R46 plus.n26 plus.n25 48.2005
R47 plus.n25 plus.n24 48.2005
R48 plus.n7 plus.n6 48.2005
R49 plus.n54 plus.n53 48.2005
R50 plus.n53 plus.n52 48.2005
R51 plus.n35 plus.n34 48.2005
R52 plus.n9 plus.n8 45.1367
R53 plus.n37 plus.n36 45.1367
R54 plus.n23 plus.n2 44.549
R55 plus.n12 plus.n11 44.549
R56 plus.n51 plus.n30 44.549
R57 plus.n40 plus.n39 44.549
R58 plus.n19 plus.n18 34.3247
R59 plus.n13 plus.n4 34.3247
R60 plus.n47 plus.n46 34.3247
R61 plus.n41 plus.n32 34.3247
R62 plus plus.n55 31.321
R63 plus.n17 plus.n4 24.1005
R64 plus.n18 plus.n17 24.1005
R65 plus.n46 plus.n45 24.1005
R66 plus.n45 plus.n32 24.1005
R67 plus.n19 plus.n2 13.8763
R68 plus.n13 plus.n12 13.8763
R69 plus.n47 plus.n30 13.8763
R70 plus.n41 plus.n40 13.8763
R71 plus.n8 plus.n7 13.3799
R72 plus.n36 plus.n35 13.3799
R73 plus plus.n27 10.0005
R74 plus.n24 plus.n23 3.65202
R75 plus.n11 plus.n6 3.65202
R76 plus.n52 plus.n51 3.65202
R77 plus.n39 plus.n34 3.65202
R78 plus.n1 plus.n0 0.285035
R79 plus.n27 plus.n0 0.285035
R80 plus.n55 plus.n28 0.285035
R81 plus.n29 plus.n28 0.285035
R82 plus.n10 plus.n9 0.189894
R83 plus.n10 plus.n5 0.189894
R84 plus.n14 plus.n5 0.189894
R85 plus.n15 plus.n14 0.189894
R86 plus.n16 plus.n15 0.189894
R87 plus.n16 plus.n3 0.189894
R88 plus.n20 plus.n3 0.189894
R89 plus.n21 plus.n20 0.189894
R90 plus.n22 plus.n21 0.189894
R91 plus.n22 plus.n1 0.189894
R92 plus.n50 plus.n29 0.189894
R93 plus.n50 plus.n49 0.189894
R94 plus.n49 plus.n48 0.189894
R95 plus.n48 plus.n31 0.189894
R96 plus.n44 plus.n31 0.189894
R97 plus.n44 plus.n43 0.189894
R98 plus.n43 plus.n42 0.189894
R99 plus.n42 plus.n33 0.189894
R100 plus.n38 plus.n33 0.189894
R101 plus.n38 plus.n37 0.189894
R102 source.n282 source.n256 289.615
R103 source.n242 source.n216 289.615
R104 source.n210 source.n184 289.615
R105 source.n170 source.n144 289.615
R106 source.n26 source.n0 289.615
R107 source.n66 source.n40 289.615
R108 source.n98 source.n72 289.615
R109 source.n138 source.n112 289.615
R110 source.n267 source.n266 185
R111 source.n264 source.n263 185
R112 source.n273 source.n272 185
R113 source.n275 source.n274 185
R114 source.n260 source.n259 185
R115 source.n281 source.n280 185
R116 source.n283 source.n282 185
R117 source.n227 source.n226 185
R118 source.n224 source.n223 185
R119 source.n233 source.n232 185
R120 source.n235 source.n234 185
R121 source.n220 source.n219 185
R122 source.n241 source.n240 185
R123 source.n243 source.n242 185
R124 source.n195 source.n194 185
R125 source.n192 source.n191 185
R126 source.n201 source.n200 185
R127 source.n203 source.n202 185
R128 source.n188 source.n187 185
R129 source.n209 source.n208 185
R130 source.n211 source.n210 185
R131 source.n155 source.n154 185
R132 source.n152 source.n151 185
R133 source.n161 source.n160 185
R134 source.n163 source.n162 185
R135 source.n148 source.n147 185
R136 source.n169 source.n168 185
R137 source.n171 source.n170 185
R138 source.n27 source.n26 185
R139 source.n25 source.n24 185
R140 source.n4 source.n3 185
R141 source.n19 source.n18 185
R142 source.n17 source.n16 185
R143 source.n8 source.n7 185
R144 source.n11 source.n10 185
R145 source.n67 source.n66 185
R146 source.n65 source.n64 185
R147 source.n44 source.n43 185
R148 source.n59 source.n58 185
R149 source.n57 source.n56 185
R150 source.n48 source.n47 185
R151 source.n51 source.n50 185
R152 source.n99 source.n98 185
R153 source.n97 source.n96 185
R154 source.n76 source.n75 185
R155 source.n91 source.n90 185
R156 source.n89 source.n88 185
R157 source.n80 source.n79 185
R158 source.n83 source.n82 185
R159 source.n139 source.n138 185
R160 source.n137 source.n136 185
R161 source.n116 source.n115 185
R162 source.n131 source.n130 185
R163 source.n129 source.n128 185
R164 source.n120 source.n119 185
R165 source.n123 source.n122 185
R166 source.t12 source.n265 147.661
R167 source.t5 source.n225 147.661
R168 source.t33 source.n193 147.661
R169 source.t22 source.n153 147.661
R170 source.t36 source.n9 147.661
R171 source.t34 source.n49 147.661
R172 source.t8 source.n81 147.661
R173 source.t0 source.n121 147.661
R174 source.n266 source.n263 104.615
R175 source.n273 source.n263 104.615
R176 source.n274 source.n273 104.615
R177 source.n274 source.n259 104.615
R178 source.n281 source.n259 104.615
R179 source.n282 source.n281 104.615
R180 source.n226 source.n223 104.615
R181 source.n233 source.n223 104.615
R182 source.n234 source.n233 104.615
R183 source.n234 source.n219 104.615
R184 source.n241 source.n219 104.615
R185 source.n242 source.n241 104.615
R186 source.n194 source.n191 104.615
R187 source.n201 source.n191 104.615
R188 source.n202 source.n201 104.615
R189 source.n202 source.n187 104.615
R190 source.n209 source.n187 104.615
R191 source.n210 source.n209 104.615
R192 source.n154 source.n151 104.615
R193 source.n161 source.n151 104.615
R194 source.n162 source.n161 104.615
R195 source.n162 source.n147 104.615
R196 source.n169 source.n147 104.615
R197 source.n170 source.n169 104.615
R198 source.n26 source.n25 104.615
R199 source.n25 source.n3 104.615
R200 source.n18 source.n3 104.615
R201 source.n18 source.n17 104.615
R202 source.n17 source.n7 104.615
R203 source.n10 source.n7 104.615
R204 source.n66 source.n65 104.615
R205 source.n65 source.n43 104.615
R206 source.n58 source.n43 104.615
R207 source.n58 source.n57 104.615
R208 source.n57 source.n47 104.615
R209 source.n50 source.n47 104.615
R210 source.n98 source.n97 104.615
R211 source.n97 source.n75 104.615
R212 source.n90 source.n75 104.615
R213 source.n90 source.n89 104.615
R214 source.n89 source.n79 104.615
R215 source.n82 source.n79 104.615
R216 source.n138 source.n137 104.615
R217 source.n137 source.n115 104.615
R218 source.n130 source.n115 104.615
R219 source.n130 source.n129 104.615
R220 source.n129 source.n119 104.615
R221 source.n122 source.n119 104.615
R222 source.n266 source.t12 52.3082
R223 source.n226 source.t5 52.3082
R224 source.n194 source.t33 52.3082
R225 source.n154 source.t22 52.3082
R226 source.n10 source.t36 52.3082
R227 source.n50 source.t34 52.3082
R228 source.n82 source.t8 52.3082
R229 source.n122 source.t0 52.3082
R230 source.n33 source.n32 50.512
R231 source.n35 source.n34 50.512
R232 source.n37 source.n36 50.512
R233 source.n39 source.n38 50.512
R234 source.n105 source.n104 50.512
R235 source.n107 source.n106 50.512
R236 source.n109 source.n108 50.512
R237 source.n111 source.n110 50.512
R238 source.n255 source.n254 50.5119
R239 source.n253 source.n252 50.5119
R240 source.n251 source.n250 50.5119
R241 source.n249 source.n248 50.5119
R242 source.n183 source.n182 50.5119
R243 source.n181 source.n180 50.5119
R244 source.n179 source.n178 50.5119
R245 source.n177 source.n176 50.5119
R246 source.n287 source.n286 32.1853
R247 source.n247 source.n246 32.1853
R248 source.n215 source.n214 32.1853
R249 source.n175 source.n174 32.1853
R250 source.n31 source.n30 32.1853
R251 source.n71 source.n70 32.1853
R252 source.n103 source.n102 32.1853
R253 source.n143 source.n142 32.1853
R254 source.n175 source.n143 17.544
R255 source.n267 source.n265 15.6674
R256 source.n227 source.n225 15.6674
R257 source.n195 source.n193 15.6674
R258 source.n155 source.n153 15.6674
R259 source.n11 source.n9 15.6674
R260 source.n51 source.n49 15.6674
R261 source.n83 source.n81 15.6674
R262 source.n123 source.n121 15.6674
R263 source.n268 source.n264 12.8005
R264 source.n228 source.n224 12.8005
R265 source.n196 source.n192 12.8005
R266 source.n156 source.n152 12.8005
R267 source.n12 source.n8 12.8005
R268 source.n52 source.n48 12.8005
R269 source.n84 source.n80 12.8005
R270 source.n124 source.n120 12.8005
R271 source.n272 source.n271 12.0247
R272 source.n232 source.n231 12.0247
R273 source.n200 source.n199 12.0247
R274 source.n160 source.n159 12.0247
R275 source.n16 source.n15 12.0247
R276 source.n56 source.n55 12.0247
R277 source.n88 source.n87 12.0247
R278 source.n128 source.n127 12.0247
R279 source.n288 source.n31 11.8802
R280 source.n275 source.n262 11.249
R281 source.n235 source.n222 11.249
R282 source.n203 source.n190 11.249
R283 source.n163 source.n150 11.249
R284 source.n19 source.n6 11.249
R285 source.n59 source.n46 11.249
R286 source.n91 source.n78 11.249
R287 source.n131 source.n118 11.249
R288 source.n276 source.n260 10.4732
R289 source.n236 source.n220 10.4732
R290 source.n204 source.n188 10.4732
R291 source.n164 source.n148 10.4732
R292 source.n20 source.n4 10.4732
R293 source.n60 source.n44 10.4732
R294 source.n92 source.n76 10.4732
R295 source.n132 source.n116 10.4732
R296 source.n280 source.n279 9.69747
R297 source.n240 source.n239 9.69747
R298 source.n208 source.n207 9.69747
R299 source.n168 source.n167 9.69747
R300 source.n24 source.n23 9.69747
R301 source.n64 source.n63 9.69747
R302 source.n96 source.n95 9.69747
R303 source.n136 source.n135 9.69747
R304 source.n286 source.n285 9.45567
R305 source.n246 source.n245 9.45567
R306 source.n214 source.n213 9.45567
R307 source.n174 source.n173 9.45567
R308 source.n30 source.n29 9.45567
R309 source.n70 source.n69 9.45567
R310 source.n102 source.n101 9.45567
R311 source.n142 source.n141 9.45567
R312 source.n285 source.n284 9.3005
R313 source.n258 source.n257 9.3005
R314 source.n279 source.n278 9.3005
R315 source.n277 source.n276 9.3005
R316 source.n262 source.n261 9.3005
R317 source.n271 source.n270 9.3005
R318 source.n269 source.n268 9.3005
R319 source.n245 source.n244 9.3005
R320 source.n218 source.n217 9.3005
R321 source.n239 source.n238 9.3005
R322 source.n237 source.n236 9.3005
R323 source.n222 source.n221 9.3005
R324 source.n231 source.n230 9.3005
R325 source.n229 source.n228 9.3005
R326 source.n213 source.n212 9.3005
R327 source.n186 source.n185 9.3005
R328 source.n207 source.n206 9.3005
R329 source.n205 source.n204 9.3005
R330 source.n190 source.n189 9.3005
R331 source.n199 source.n198 9.3005
R332 source.n197 source.n196 9.3005
R333 source.n173 source.n172 9.3005
R334 source.n146 source.n145 9.3005
R335 source.n167 source.n166 9.3005
R336 source.n165 source.n164 9.3005
R337 source.n150 source.n149 9.3005
R338 source.n159 source.n158 9.3005
R339 source.n157 source.n156 9.3005
R340 source.n29 source.n28 9.3005
R341 source.n2 source.n1 9.3005
R342 source.n23 source.n22 9.3005
R343 source.n21 source.n20 9.3005
R344 source.n6 source.n5 9.3005
R345 source.n15 source.n14 9.3005
R346 source.n13 source.n12 9.3005
R347 source.n69 source.n68 9.3005
R348 source.n42 source.n41 9.3005
R349 source.n63 source.n62 9.3005
R350 source.n61 source.n60 9.3005
R351 source.n46 source.n45 9.3005
R352 source.n55 source.n54 9.3005
R353 source.n53 source.n52 9.3005
R354 source.n101 source.n100 9.3005
R355 source.n74 source.n73 9.3005
R356 source.n95 source.n94 9.3005
R357 source.n93 source.n92 9.3005
R358 source.n78 source.n77 9.3005
R359 source.n87 source.n86 9.3005
R360 source.n85 source.n84 9.3005
R361 source.n141 source.n140 9.3005
R362 source.n114 source.n113 9.3005
R363 source.n135 source.n134 9.3005
R364 source.n133 source.n132 9.3005
R365 source.n118 source.n117 9.3005
R366 source.n127 source.n126 9.3005
R367 source.n125 source.n124 9.3005
R368 source.n283 source.n258 8.92171
R369 source.n243 source.n218 8.92171
R370 source.n211 source.n186 8.92171
R371 source.n171 source.n146 8.92171
R372 source.n27 source.n2 8.92171
R373 source.n67 source.n42 8.92171
R374 source.n99 source.n74 8.92171
R375 source.n139 source.n114 8.92171
R376 source.n284 source.n256 8.14595
R377 source.n244 source.n216 8.14595
R378 source.n212 source.n184 8.14595
R379 source.n172 source.n144 8.14595
R380 source.n28 source.n0 8.14595
R381 source.n68 source.n40 8.14595
R382 source.n100 source.n72 8.14595
R383 source.n140 source.n112 8.14595
R384 source.n286 source.n256 5.81868
R385 source.n246 source.n216 5.81868
R386 source.n214 source.n184 5.81868
R387 source.n174 source.n144 5.81868
R388 source.n30 source.n0 5.81868
R389 source.n70 source.n40 5.81868
R390 source.n102 source.n72 5.81868
R391 source.n142 source.n112 5.81868
R392 source.n288 source.n287 5.66429
R393 source.n284 source.n283 5.04292
R394 source.n244 source.n243 5.04292
R395 source.n212 source.n211 5.04292
R396 source.n172 source.n171 5.04292
R397 source.n28 source.n27 5.04292
R398 source.n68 source.n67 5.04292
R399 source.n100 source.n99 5.04292
R400 source.n140 source.n139 5.04292
R401 source.n269 source.n265 4.38594
R402 source.n229 source.n225 4.38594
R403 source.n197 source.n193 4.38594
R404 source.n157 source.n153 4.38594
R405 source.n13 source.n9 4.38594
R406 source.n53 source.n49 4.38594
R407 source.n85 source.n81 4.38594
R408 source.n125 source.n121 4.38594
R409 source.n280 source.n258 4.26717
R410 source.n240 source.n218 4.26717
R411 source.n208 source.n186 4.26717
R412 source.n168 source.n146 4.26717
R413 source.n24 source.n2 4.26717
R414 source.n64 source.n42 4.26717
R415 source.n96 source.n74 4.26717
R416 source.n136 source.n114 4.26717
R417 source.n279 source.n260 3.49141
R418 source.n239 source.n220 3.49141
R419 source.n207 source.n188 3.49141
R420 source.n167 source.n148 3.49141
R421 source.n23 source.n4 3.49141
R422 source.n63 source.n44 3.49141
R423 source.n95 source.n76 3.49141
R424 source.n135 source.n116 3.49141
R425 source.n254 source.t16 3.3005
R426 source.n254 source.t18 3.3005
R427 source.n252 source.t14 3.3005
R428 source.n252 source.t9 3.3005
R429 source.n250 source.t15 3.3005
R430 source.n250 source.t7 3.3005
R431 source.n248 source.t11 3.3005
R432 source.n248 source.t6 3.3005
R433 source.n182 source.t28 3.3005
R434 source.n182 source.t32 3.3005
R435 source.n180 source.t25 3.3005
R436 source.n180 source.t39 3.3005
R437 source.n178 source.t27 3.3005
R438 source.n178 source.t31 3.3005
R439 source.n176 source.t24 3.3005
R440 source.n176 source.t20 3.3005
R441 source.n32 source.t21 3.3005
R442 source.n32 source.t38 3.3005
R443 source.n34 source.t23 3.3005
R444 source.n34 source.t26 3.3005
R445 source.n36 source.t30 3.3005
R446 source.n36 source.t35 3.3005
R447 source.n38 source.t37 3.3005
R448 source.n38 source.t29 3.3005
R449 source.n104 source.t4 3.3005
R450 source.n104 source.t17 3.3005
R451 source.n106 source.t10 3.3005
R452 source.n106 source.t2 3.3005
R453 source.n108 source.t19 3.3005
R454 source.n108 source.t13 3.3005
R455 source.n110 source.t1 3.3005
R456 source.n110 source.t3 3.3005
R457 source.n276 source.n275 2.71565
R458 source.n236 source.n235 2.71565
R459 source.n204 source.n203 2.71565
R460 source.n164 source.n163 2.71565
R461 source.n20 source.n19 2.71565
R462 source.n60 source.n59 2.71565
R463 source.n92 source.n91 2.71565
R464 source.n132 source.n131 2.71565
R465 source.n272 source.n262 1.93989
R466 source.n232 source.n222 1.93989
R467 source.n200 source.n190 1.93989
R468 source.n160 source.n150 1.93989
R469 source.n16 source.n6 1.93989
R470 source.n56 source.n46 1.93989
R471 source.n88 source.n78 1.93989
R472 source.n128 source.n118 1.93989
R473 source.n271 source.n264 1.16414
R474 source.n231 source.n224 1.16414
R475 source.n199 source.n192 1.16414
R476 source.n159 source.n152 1.16414
R477 source.n15 source.n8 1.16414
R478 source.n55 source.n48 1.16414
R479 source.n87 source.n80 1.16414
R480 source.n127 source.n120 1.16414
R481 source.n143 source.n111 0.802224
R482 source.n111 source.n109 0.802224
R483 source.n109 source.n107 0.802224
R484 source.n107 source.n105 0.802224
R485 source.n105 source.n103 0.802224
R486 source.n71 source.n39 0.802224
R487 source.n39 source.n37 0.802224
R488 source.n37 source.n35 0.802224
R489 source.n35 source.n33 0.802224
R490 source.n33 source.n31 0.802224
R491 source.n177 source.n175 0.802224
R492 source.n179 source.n177 0.802224
R493 source.n181 source.n179 0.802224
R494 source.n183 source.n181 0.802224
R495 source.n215 source.n183 0.802224
R496 source.n249 source.n247 0.802224
R497 source.n251 source.n249 0.802224
R498 source.n253 source.n251 0.802224
R499 source.n255 source.n253 0.802224
R500 source.n287 source.n255 0.802224
R501 source.n103 source.n71 0.470328
R502 source.n247 source.n215 0.470328
R503 source.n268 source.n267 0.388379
R504 source.n228 source.n227 0.388379
R505 source.n196 source.n195 0.388379
R506 source.n156 source.n155 0.388379
R507 source.n12 source.n11 0.388379
R508 source.n52 source.n51 0.388379
R509 source.n84 source.n83 0.388379
R510 source.n124 source.n123 0.388379
R511 source source.n288 0.188
R512 source.n270 source.n269 0.155672
R513 source.n270 source.n261 0.155672
R514 source.n277 source.n261 0.155672
R515 source.n278 source.n277 0.155672
R516 source.n278 source.n257 0.155672
R517 source.n285 source.n257 0.155672
R518 source.n230 source.n229 0.155672
R519 source.n230 source.n221 0.155672
R520 source.n237 source.n221 0.155672
R521 source.n238 source.n237 0.155672
R522 source.n238 source.n217 0.155672
R523 source.n245 source.n217 0.155672
R524 source.n198 source.n197 0.155672
R525 source.n198 source.n189 0.155672
R526 source.n205 source.n189 0.155672
R527 source.n206 source.n205 0.155672
R528 source.n206 source.n185 0.155672
R529 source.n213 source.n185 0.155672
R530 source.n158 source.n157 0.155672
R531 source.n158 source.n149 0.155672
R532 source.n165 source.n149 0.155672
R533 source.n166 source.n165 0.155672
R534 source.n166 source.n145 0.155672
R535 source.n173 source.n145 0.155672
R536 source.n29 source.n1 0.155672
R537 source.n22 source.n1 0.155672
R538 source.n22 source.n21 0.155672
R539 source.n21 source.n5 0.155672
R540 source.n14 source.n5 0.155672
R541 source.n14 source.n13 0.155672
R542 source.n69 source.n41 0.155672
R543 source.n62 source.n41 0.155672
R544 source.n62 source.n61 0.155672
R545 source.n61 source.n45 0.155672
R546 source.n54 source.n45 0.155672
R547 source.n54 source.n53 0.155672
R548 source.n101 source.n73 0.155672
R549 source.n94 source.n73 0.155672
R550 source.n94 source.n93 0.155672
R551 source.n93 source.n77 0.155672
R552 source.n86 source.n77 0.155672
R553 source.n86 source.n85 0.155672
R554 source.n141 source.n113 0.155672
R555 source.n134 source.n113 0.155672
R556 source.n134 source.n133 0.155672
R557 source.n133 source.n117 0.155672
R558 source.n126 source.n117 0.155672
R559 source.n126 source.n125 0.155672
R560 drain_left.n10 drain_left.n8 67.9925
R561 drain_left.n6 drain_left.n4 67.9924
R562 drain_left.n2 drain_left.n0 67.9924
R563 drain_left.n14 drain_left.n13 67.1908
R564 drain_left.n12 drain_left.n11 67.1908
R565 drain_left.n10 drain_left.n9 67.1908
R566 drain_left.n16 drain_left.n15 67.1907
R567 drain_left.n7 drain_left.n3 67.1907
R568 drain_left.n6 drain_left.n5 67.1907
R569 drain_left.n2 drain_left.n1 67.1907
R570 drain_left drain_left.n7 29.2354
R571 drain_left drain_left.n16 6.45494
R572 drain_left.n3 drain_left.t1 3.3005
R573 drain_left.n3 drain_left.t2 3.3005
R574 drain_left.n4 drain_left.t18 3.3005
R575 drain_left.n4 drain_left.t9 3.3005
R576 drain_left.n5 drain_left.t8 3.3005
R577 drain_left.n5 drain_left.t13 3.3005
R578 drain_left.n1 drain_left.t7 3.3005
R579 drain_left.n1 drain_left.t12 3.3005
R580 drain_left.n0 drain_left.t11 3.3005
R581 drain_left.n0 drain_left.t0 3.3005
R582 drain_left.n15 drain_left.t17 3.3005
R583 drain_left.n15 drain_left.t19 3.3005
R584 drain_left.n13 drain_left.t15 3.3005
R585 drain_left.n13 drain_left.t16 3.3005
R586 drain_left.n11 drain_left.t10 3.3005
R587 drain_left.n11 drain_left.t14 3.3005
R588 drain_left.n9 drain_left.t5 3.3005
R589 drain_left.n9 drain_left.t6 3.3005
R590 drain_left.n8 drain_left.t3 3.3005
R591 drain_left.n8 drain_left.t4 3.3005
R592 drain_left.n12 drain_left.n10 0.802224
R593 drain_left.n14 drain_left.n12 0.802224
R594 drain_left.n16 drain_left.n14 0.802224
R595 drain_left.n7 drain_left.n6 0.746878
R596 drain_left.n7 drain_left.n2 0.746878
R597 minus.n6 minus.t14 333.293
R598 minus.n34 minus.t7 333.293
R599 minus.n7 minus.t13 306.473
R600 minus.n8 minus.t12 306.473
R601 minus.n12 minus.t10 306.473
R602 minus.n14 minus.t5 306.473
R603 minus.n18 minus.t8 306.473
R604 minus.n20 minus.t6 306.473
R605 minus.n24 minus.t2 306.473
R606 minus.n25 minus.t1 306.473
R607 minus.n26 minus.t0 306.473
R608 minus.n35 minus.t17 306.473
R609 minus.n36 minus.t19 306.473
R610 minus.n40 minus.t11 306.473
R611 minus.n42 minus.t16 306.473
R612 minus.n46 minus.t15 306.473
R613 minus.n48 minus.t3 306.473
R614 minus.n52 minus.t9 306.473
R615 minus.n53 minus.t18 306.473
R616 minus.n54 minus.t4 306.473
R617 minus.n27 minus.n26 161.3
R618 minus.n24 minus.n23 161.3
R619 minus.n22 minus.n1 161.3
R620 minus.n21 minus.n20 161.3
R621 minus.n19 minus.n2 161.3
R622 minus.n18 minus.n17 161.3
R623 minus.n16 minus.n3 161.3
R624 minus.n15 minus.n14 161.3
R625 minus.n13 minus.n4 161.3
R626 minus.n12 minus.n11 161.3
R627 minus.n10 minus.n5 161.3
R628 minus.n9 minus.n8 161.3
R629 minus.n55 minus.n54 161.3
R630 minus.n52 minus.n51 161.3
R631 minus.n50 minus.n29 161.3
R632 minus.n49 minus.n48 161.3
R633 minus.n47 minus.n30 161.3
R634 minus.n46 minus.n45 161.3
R635 minus.n44 minus.n31 161.3
R636 minus.n43 minus.n42 161.3
R637 minus.n41 minus.n32 161.3
R638 minus.n40 minus.n39 161.3
R639 minus.n38 minus.n33 161.3
R640 minus.n37 minus.n36 161.3
R641 minus.n25 minus.n0 80.6037
R642 minus.n53 minus.n28 80.6037
R643 minus.n8 minus.n7 48.2005
R644 minus.n25 minus.n24 48.2005
R645 minus.n26 minus.n25 48.2005
R646 minus.n36 minus.n35 48.2005
R647 minus.n53 minus.n52 48.2005
R648 minus.n54 minus.n53 48.2005
R649 minus.n9 minus.n6 45.1367
R650 minus.n37 minus.n34 45.1367
R651 minus.n12 minus.n5 44.549
R652 minus.n20 minus.n1 44.549
R653 minus.n40 minus.n33 44.549
R654 minus.n48 minus.n29 44.549
R655 minus.n56 minus.n27 35.1672
R656 minus.n14 minus.n13 34.3247
R657 minus.n19 minus.n18 34.3247
R658 minus.n42 minus.n41 34.3247
R659 minus.n47 minus.n46 34.3247
R660 minus.n18 minus.n3 24.1005
R661 minus.n14 minus.n3 24.1005
R662 minus.n42 minus.n31 24.1005
R663 minus.n46 minus.n31 24.1005
R664 minus.n13 minus.n12 13.8763
R665 minus.n20 minus.n19 13.8763
R666 minus.n41 minus.n40 13.8763
R667 minus.n48 minus.n47 13.8763
R668 minus.n7 minus.n6 13.3799
R669 minus.n35 minus.n34 13.3799
R670 minus.n56 minus.n55 6.62929
R671 minus.n8 minus.n5 3.65202
R672 minus.n24 minus.n1 3.65202
R673 minus.n36 minus.n33 3.65202
R674 minus.n52 minus.n29 3.65202
R675 minus.n27 minus.n0 0.285035
R676 minus.n23 minus.n0 0.285035
R677 minus.n51 minus.n28 0.285035
R678 minus.n55 minus.n28 0.285035
R679 minus.n23 minus.n22 0.189894
R680 minus.n22 minus.n21 0.189894
R681 minus.n21 minus.n2 0.189894
R682 minus.n17 minus.n2 0.189894
R683 minus.n17 minus.n16 0.189894
R684 minus.n16 minus.n15 0.189894
R685 minus.n15 minus.n4 0.189894
R686 minus.n11 minus.n4 0.189894
R687 minus.n11 minus.n10 0.189894
R688 minus.n10 minus.n9 0.189894
R689 minus.n38 minus.n37 0.189894
R690 minus.n39 minus.n38 0.189894
R691 minus.n39 minus.n32 0.189894
R692 minus.n43 minus.n32 0.189894
R693 minus.n44 minus.n43 0.189894
R694 minus.n45 minus.n44 0.189894
R695 minus.n45 minus.n30 0.189894
R696 minus.n49 minus.n30 0.189894
R697 minus.n50 minus.n49 0.189894
R698 minus.n51 minus.n50 0.189894
R699 minus minus.n56 0.188
R700 drain_right.n6 drain_right.n4 67.9924
R701 drain_right.n2 drain_right.n0 67.9924
R702 drain_right.n10 drain_right.n8 67.9924
R703 drain_right.n10 drain_right.n9 67.1908
R704 drain_right.n12 drain_right.n11 67.1908
R705 drain_right.n14 drain_right.n13 67.1908
R706 drain_right.n16 drain_right.n15 67.1908
R707 drain_right.n7 drain_right.n3 67.1907
R708 drain_right.n6 drain_right.n5 67.1907
R709 drain_right.n2 drain_right.n1 67.1907
R710 drain_right drain_right.n7 28.6822
R711 drain_right drain_right.n16 6.45494
R712 drain_right.n3 drain_right.t3 3.3005
R713 drain_right.n3 drain_right.t4 3.3005
R714 drain_right.n4 drain_right.t1 3.3005
R715 drain_right.n4 drain_right.t15 3.3005
R716 drain_right.n5 drain_right.t16 3.3005
R717 drain_right.n5 drain_right.t10 3.3005
R718 drain_right.n1 drain_right.t0 3.3005
R719 drain_right.n1 drain_right.t8 3.3005
R720 drain_right.n0 drain_right.t12 3.3005
R721 drain_right.n0 drain_right.t2 3.3005
R722 drain_right.n8 drain_right.t6 3.3005
R723 drain_right.n8 drain_right.t5 3.3005
R724 drain_right.n9 drain_right.t9 3.3005
R725 drain_right.n9 drain_right.t7 3.3005
R726 drain_right.n11 drain_right.t11 3.3005
R727 drain_right.n11 drain_right.t14 3.3005
R728 drain_right.n13 drain_right.t17 3.3005
R729 drain_right.n13 drain_right.t13 3.3005
R730 drain_right.n15 drain_right.t19 3.3005
R731 drain_right.n15 drain_right.t18 3.3005
R732 drain_right.n16 drain_right.n14 0.802224
R733 drain_right.n14 drain_right.n12 0.802224
R734 drain_right.n12 drain_right.n10 0.802224
R735 drain_right.n7 drain_right.n6 0.746878
R736 drain_right.n7 drain_right.n2 0.746878
C0 drain_right minus 6.08018f
C1 drain_left source 14.9889f
C2 minus plus 5.48165f
C3 drain_left minus 0.173552f
C4 drain_right plus 0.431663f
C5 minus source 6.4822f
C6 drain_left drain_right 1.48676f
C7 drain_left plus 6.35483f
C8 drain_right source 14.990701f
C9 source plus 6.49621f
C10 drain_right a_n2762_n2088# 5.99527f
C11 drain_left a_n2762_n2088# 6.3961f
C12 source a_n2762_n2088# 5.740417f
C13 minus a_n2762_n2088# 10.534765f
C14 plus a_n2762_n2088# 12.10784f
C15 drain_right.t12 a_n2762_n2088# 0.132342f
C16 drain_right.t2 a_n2762_n2088# 0.132342f
C17 drain_right.n0 a_n2762_n2088# 1.10824f
C18 drain_right.t0 a_n2762_n2088# 0.132342f
C19 drain_right.t8 a_n2762_n2088# 0.132342f
C20 drain_right.n1 a_n2762_n2088# 1.10373f
C21 drain_right.n2 a_n2762_n2088# 0.744143f
C22 drain_right.t3 a_n2762_n2088# 0.132342f
C23 drain_right.t4 a_n2762_n2088# 0.132342f
C24 drain_right.n3 a_n2762_n2088# 1.10373f
C25 drain_right.t1 a_n2762_n2088# 0.132342f
C26 drain_right.t15 a_n2762_n2088# 0.132342f
C27 drain_right.n4 a_n2762_n2088# 1.10824f
C28 drain_right.t16 a_n2762_n2088# 0.132342f
C29 drain_right.t10 a_n2762_n2088# 0.132342f
C30 drain_right.n5 a_n2762_n2088# 1.10373f
C31 drain_right.n6 a_n2762_n2088# 0.744143f
C32 drain_right.n7 a_n2762_n2088# 1.52873f
C33 drain_right.t6 a_n2762_n2088# 0.132342f
C34 drain_right.t5 a_n2762_n2088# 0.132342f
C35 drain_right.n8 a_n2762_n2088# 1.10824f
C36 drain_right.t9 a_n2762_n2088# 0.132342f
C37 drain_right.t7 a_n2762_n2088# 0.132342f
C38 drain_right.n9 a_n2762_n2088# 1.10374f
C39 drain_right.n10 a_n2762_n2088# 0.748248f
C40 drain_right.t11 a_n2762_n2088# 0.132342f
C41 drain_right.t14 a_n2762_n2088# 0.132342f
C42 drain_right.n11 a_n2762_n2088# 1.10374f
C43 drain_right.n12 a_n2762_n2088# 0.370753f
C44 drain_right.t17 a_n2762_n2088# 0.132342f
C45 drain_right.t13 a_n2762_n2088# 0.132342f
C46 drain_right.n13 a_n2762_n2088# 1.10374f
C47 drain_right.n14 a_n2762_n2088# 0.370753f
C48 drain_right.t19 a_n2762_n2088# 0.132342f
C49 drain_right.t18 a_n2762_n2088# 0.132342f
C50 drain_right.n15 a_n2762_n2088# 1.10374f
C51 drain_right.n16 a_n2762_n2088# 0.614144f
C52 minus.n0 a_n2762_n2088# 0.056694f
C53 minus.n1 a_n2762_n2088# 0.009664f
C54 minus.t2 a_n2762_n2088# 0.44469f
C55 minus.n2 a_n2762_n2088# 0.042587f
C56 minus.n3 a_n2762_n2088# 0.009664f
C57 minus.t8 a_n2762_n2088# 0.44469f
C58 minus.n4 a_n2762_n2088# 0.042587f
C59 minus.n5 a_n2762_n2088# 0.009664f
C60 minus.t10 a_n2762_n2088# 0.44469f
C61 minus.t14 a_n2762_n2088# 0.461402f
C62 minus.n6 a_n2762_n2088# 0.191746f
C63 minus.t13 a_n2762_n2088# 0.44469f
C64 minus.n7 a_n2762_n2088# 0.217206f
C65 minus.t12 a_n2762_n2088# 0.44469f
C66 minus.n8 a_n2762_n2088# 0.208199f
C67 minus.n9 a_n2762_n2088# 0.181773f
C68 minus.n10 a_n2762_n2088# 0.042587f
C69 minus.n11 a_n2762_n2088# 0.042587f
C70 minus.n12 a_n2762_n2088# 0.209381f
C71 minus.n13 a_n2762_n2088# 0.009664f
C72 minus.t5 a_n2762_n2088# 0.44469f
C73 minus.n14 a_n2762_n2088# 0.209381f
C74 minus.n15 a_n2762_n2088# 0.042587f
C75 minus.n16 a_n2762_n2088# 0.042587f
C76 minus.n17 a_n2762_n2088# 0.042587f
C77 minus.n18 a_n2762_n2088# 0.209381f
C78 minus.n19 a_n2762_n2088# 0.009664f
C79 minus.t6 a_n2762_n2088# 0.44469f
C80 minus.n20 a_n2762_n2088# 0.209381f
C81 minus.n21 a_n2762_n2088# 0.042587f
C82 minus.n22 a_n2762_n2088# 0.042587f
C83 minus.n23 a_n2762_n2088# 0.056827f
C84 minus.n24 a_n2762_n2088# 0.208199f
C85 minus.t1 a_n2762_n2088# 0.44469f
C86 minus.n25 a_n2762_n2088# 0.217206f
C87 minus.t0 a_n2762_n2088# 0.44469f
C88 minus.n26 a_n2762_n2088# 0.207543f
C89 minus.n27 a_n2762_n2088# 1.45705f
C90 minus.n28 a_n2762_n2088# 0.056694f
C91 minus.n29 a_n2762_n2088# 0.009664f
C92 minus.n30 a_n2762_n2088# 0.042587f
C93 minus.n31 a_n2762_n2088# 0.009664f
C94 minus.n32 a_n2762_n2088# 0.042587f
C95 minus.n33 a_n2762_n2088# 0.009664f
C96 minus.t7 a_n2762_n2088# 0.461402f
C97 minus.n34 a_n2762_n2088# 0.191746f
C98 minus.t17 a_n2762_n2088# 0.44469f
C99 minus.n35 a_n2762_n2088# 0.217206f
C100 minus.t19 a_n2762_n2088# 0.44469f
C101 minus.n36 a_n2762_n2088# 0.208199f
C102 minus.n37 a_n2762_n2088# 0.181773f
C103 minus.n38 a_n2762_n2088# 0.042587f
C104 minus.n39 a_n2762_n2088# 0.042587f
C105 minus.t11 a_n2762_n2088# 0.44469f
C106 minus.n40 a_n2762_n2088# 0.209381f
C107 minus.n41 a_n2762_n2088# 0.009664f
C108 minus.t16 a_n2762_n2088# 0.44469f
C109 minus.n42 a_n2762_n2088# 0.209381f
C110 minus.n43 a_n2762_n2088# 0.042587f
C111 minus.n44 a_n2762_n2088# 0.042587f
C112 minus.n45 a_n2762_n2088# 0.042587f
C113 minus.t15 a_n2762_n2088# 0.44469f
C114 minus.n46 a_n2762_n2088# 0.209381f
C115 minus.n47 a_n2762_n2088# 0.009664f
C116 minus.t3 a_n2762_n2088# 0.44469f
C117 minus.n48 a_n2762_n2088# 0.209381f
C118 minus.n49 a_n2762_n2088# 0.042587f
C119 minus.n50 a_n2762_n2088# 0.042587f
C120 minus.n51 a_n2762_n2088# 0.056827f
C121 minus.t9 a_n2762_n2088# 0.44469f
C122 minus.n52 a_n2762_n2088# 0.208199f
C123 minus.t18 a_n2762_n2088# 0.44469f
C124 minus.n53 a_n2762_n2088# 0.217206f
C125 minus.t4 a_n2762_n2088# 0.44469f
C126 minus.n54 a_n2762_n2088# 0.207543f
C127 minus.n55 a_n2762_n2088# 0.305554f
C128 minus.n56 a_n2762_n2088# 1.75317f
C129 drain_left.t11 a_n2762_n2088# 0.133533f
C130 drain_left.t0 a_n2762_n2088# 0.133533f
C131 drain_left.n0 a_n2762_n2088# 1.11821f
C132 drain_left.t7 a_n2762_n2088# 0.133533f
C133 drain_left.t12 a_n2762_n2088# 0.133533f
C134 drain_left.n1 a_n2762_n2088# 1.11366f
C135 drain_left.n2 a_n2762_n2088# 0.750838f
C136 drain_left.t1 a_n2762_n2088# 0.133533f
C137 drain_left.t2 a_n2762_n2088# 0.133533f
C138 drain_left.n3 a_n2762_n2088# 1.11366f
C139 drain_left.t18 a_n2762_n2088# 0.133533f
C140 drain_left.t9 a_n2762_n2088# 0.133533f
C141 drain_left.n4 a_n2762_n2088# 1.11821f
C142 drain_left.t8 a_n2762_n2088# 0.133533f
C143 drain_left.t13 a_n2762_n2088# 0.133533f
C144 drain_left.n5 a_n2762_n2088# 1.11366f
C145 drain_left.n6 a_n2762_n2088# 0.750838f
C146 drain_left.n7 a_n2762_n2088# 1.59886f
C147 drain_left.t3 a_n2762_n2088# 0.133533f
C148 drain_left.t4 a_n2762_n2088# 0.133533f
C149 drain_left.n8 a_n2762_n2088# 1.11821f
C150 drain_left.t5 a_n2762_n2088# 0.133533f
C151 drain_left.t6 a_n2762_n2088# 0.133533f
C152 drain_left.n9 a_n2762_n2088# 1.11367f
C153 drain_left.n10 a_n2762_n2088# 0.754975f
C154 drain_left.t10 a_n2762_n2088# 0.133533f
C155 drain_left.t14 a_n2762_n2088# 0.133533f
C156 drain_left.n11 a_n2762_n2088# 1.11367f
C157 drain_left.n12 a_n2762_n2088# 0.374088f
C158 drain_left.t15 a_n2762_n2088# 0.133533f
C159 drain_left.t16 a_n2762_n2088# 0.133533f
C160 drain_left.n13 a_n2762_n2088# 1.11367f
C161 drain_left.n14 a_n2762_n2088# 0.374088f
C162 drain_left.t17 a_n2762_n2088# 0.133533f
C163 drain_left.t19 a_n2762_n2088# 0.133533f
C164 drain_left.n15 a_n2762_n2088# 1.11366f
C165 drain_left.n16 a_n2762_n2088# 0.619675f
C166 source.n0 a_n2762_n2088# 0.037321f
C167 source.n1 a_n2762_n2088# 0.026552f
C168 source.n2 a_n2762_n2088# 0.014268f
C169 source.n3 a_n2762_n2088# 0.033724f
C170 source.n4 a_n2762_n2088# 0.015107f
C171 source.n5 a_n2762_n2088# 0.026552f
C172 source.n6 a_n2762_n2088# 0.014268f
C173 source.n7 a_n2762_n2088# 0.033724f
C174 source.n8 a_n2762_n2088# 0.015107f
C175 source.n9 a_n2762_n2088# 0.113624f
C176 source.t36 a_n2762_n2088# 0.054966f
C177 source.n10 a_n2762_n2088# 0.025293f
C178 source.n11 a_n2762_n2088# 0.01992f
C179 source.n12 a_n2762_n2088# 0.014268f
C180 source.n13 a_n2762_n2088# 0.631779f
C181 source.n14 a_n2762_n2088# 0.026552f
C182 source.n15 a_n2762_n2088# 0.014268f
C183 source.n16 a_n2762_n2088# 0.015107f
C184 source.n17 a_n2762_n2088# 0.033724f
C185 source.n18 a_n2762_n2088# 0.033724f
C186 source.n19 a_n2762_n2088# 0.015107f
C187 source.n20 a_n2762_n2088# 0.014268f
C188 source.n21 a_n2762_n2088# 0.026552f
C189 source.n22 a_n2762_n2088# 0.026552f
C190 source.n23 a_n2762_n2088# 0.014268f
C191 source.n24 a_n2762_n2088# 0.015107f
C192 source.n25 a_n2762_n2088# 0.033724f
C193 source.n26 a_n2762_n2088# 0.073007f
C194 source.n27 a_n2762_n2088# 0.015107f
C195 source.n28 a_n2762_n2088# 0.014268f
C196 source.n29 a_n2762_n2088# 0.061374f
C197 source.n30 a_n2762_n2088# 0.04085f
C198 source.n31 a_n2762_n2088# 0.681027f
C199 source.t21 a_n2762_n2088# 0.125893f
C200 source.t38 a_n2762_n2088# 0.125893f
C201 source.n32 a_n2762_n2088# 0.980466f
C202 source.n33 a_n2762_n2088# 0.386085f
C203 source.t23 a_n2762_n2088# 0.125893f
C204 source.t26 a_n2762_n2088# 0.125893f
C205 source.n34 a_n2762_n2088# 0.980466f
C206 source.n35 a_n2762_n2088# 0.386085f
C207 source.t30 a_n2762_n2088# 0.125893f
C208 source.t35 a_n2762_n2088# 0.125893f
C209 source.n36 a_n2762_n2088# 0.980466f
C210 source.n37 a_n2762_n2088# 0.386085f
C211 source.t37 a_n2762_n2088# 0.125893f
C212 source.t29 a_n2762_n2088# 0.125893f
C213 source.n38 a_n2762_n2088# 0.980466f
C214 source.n39 a_n2762_n2088# 0.386085f
C215 source.n40 a_n2762_n2088# 0.037321f
C216 source.n41 a_n2762_n2088# 0.026552f
C217 source.n42 a_n2762_n2088# 0.014268f
C218 source.n43 a_n2762_n2088# 0.033724f
C219 source.n44 a_n2762_n2088# 0.015107f
C220 source.n45 a_n2762_n2088# 0.026552f
C221 source.n46 a_n2762_n2088# 0.014268f
C222 source.n47 a_n2762_n2088# 0.033724f
C223 source.n48 a_n2762_n2088# 0.015107f
C224 source.n49 a_n2762_n2088# 0.113624f
C225 source.t34 a_n2762_n2088# 0.054966f
C226 source.n50 a_n2762_n2088# 0.025293f
C227 source.n51 a_n2762_n2088# 0.01992f
C228 source.n52 a_n2762_n2088# 0.014268f
C229 source.n53 a_n2762_n2088# 0.631779f
C230 source.n54 a_n2762_n2088# 0.026552f
C231 source.n55 a_n2762_n2088# 0.014268f
C232 source.n56 a_n2762_n2088# 0.015107f
C233 source.n57 a_n2762_n2088# 0.033724f
C234 source.n58 a_n2762_n2088# 0.033724f
C235 source.n59 a_n2762_n2088# 0.015107f
C236 source.n60 a_n2762_n2088# 0.014268f
C237 source.n61 a_n2762_n2088# 0.026552f
C238 source.n62 a_n2762_n2088# 0.026552f
C239 source.n63 a_n2762_n2088# 0.014268f
C240 source.n64 a_n2762_n2088# 0.015107f
C241 source.n65 a_n2762_n2088# 0.033724f
C242 source.n66 a_n2762_n2088# 0.073007f
C243 source.n67 a_n2762_n2088# 0.015107f
C244 source.n68 a_n2762_n2088# 0.014268f
C245 source.n69 a_n2762_n2088# 0.061374f
C246 source.n70 a_n2762_n2088# 0.04085f
C247 source.n71 a_n2762_n2088# 0.131467f
C248 source.n72 a_n2762_n2088# 0.037321f
C249 source.n73 a_n2762_n2088# 0.026552f
C250 source.n74 a_n2762_n2088# 0.014268f
C251 source.n75 a_n2762_n2088# 0.033724f
C252 source.n76 a_n2762_n2088# 0.015107f
C253 source.n77 a_n2762_n2088# 0.026552f
C254 source.n78 a_n2762_n2088# 0.014268f
C255 source.n79 a_n2762_n2088# 0.033724f
C256 source.n80 a_n2762_n2088# 0.015107f
C257 source.n81 a_n2762_n2088# 0.113624f
C258 source.t8 a_n2762_n2088# 0.054966f
C259 source.n82 a_n2762_n2088# 0.025293f
C260 source.n83 a_n2762_n2088# 0.01992f
C261 source.n84 a_n2762_n2088# 0.014268f
C262 source.n85 a_n2762_n2088# 0.631779f
C263 source.n86 a_n2762_n2088# 0.026552f
C264 source.n87 a_n2762_n2088# 0.014268f
C265 source.n88 a_n2762_n2088# 0.015107f
C266 source.n89 a_n2762_n2088# 0.033724f
C267 source.n90 a_n2762_n2088# 0.033724f
C268 source.n91 a_n2762_n2088# 0.015107f
C269 source.n92 a_n2762_n2088# 0.014268f
C270 source.n93 a_n2762_n2088# 0.026552f
C271 source.n94 a_n2762_n2088# 0.026552f
C272 source.n95 a_n2762_n2088# 0.014268f
C273 source.n96 a_n2762_n2088# 0.015107f
C274 source.n97 a_n2762_n2088# 0.033724f
C275 source.n98 a_n2762_n2088# 0.073007f
C276 source.n99 a_n2762_n2088# 0.015107f
C277 source.n100 a_n2762_n2088# 0.014268f
C278 source.n101 a_n2762_n2088# 0.061374f
C279 source.n102 a_n2762_n2088# 0.04085f
C280 source.n103 a_n2762_n2088# 0.131467f
C281 source.t4 a_n2762_n2088# 0.125893f
C282 source.t17 a_n2762_n2088# 0.125893f
C283 source.n104 a_n2762_n2088# 0.980466f
C284 source.n105 a_n2762_n2088# 0.386085f
C285 source.t10 a_n2762_n2088# 0.125893f
C286 source.t2 a_n2762_n2088# 0.125893f
C287 source.n106 a_n2762_n2088# 0.980466f
C288 source.n107 a_n2762_n2088# 0.386085f
C289 source.t19 a_n2762_n2088# 0.125893f
C290 source.t13 a_n2762_n2088# 0.125893f
C291 source.n108 a_n2762_n2088# 0.980466f
C292 source.n109 a_n2762_n2088# 0.386085f
C293 source.t1 a_n2762_n2088# 0.125893f
C294 source.t3 a_n2762_n2088# 0.125893f
C295 source.n110 a_n2762_n2088# 0.980466f
C296 source.n111 a_n2762_n2088# 0.386085f
C297 source.n112 a_n2762_n2088# 0.037321f
C298 source.n113 a_n2762_n2088# 0.026552f
C299 source.n114 a_n2762_n2088# 0.014268f
C300 source.n115 a_n2762_n2088# 0.033724f
C301 source.n116 a_n2762_n2088# 0.015107f
C302 source.n117 a_n2762_n2088# 0.026552f
C303 source.n118 a_n2762_n2088# 0.014268f
C304 source.n119 a_n2762_n2088# 0.033724f
C305 source.n120 a_n2762_n2088# 0.015107f
C306 source.n121 a_n2762_n2088# 0.113624f
C307 source.t0 a_n2762_n2088# 0.054966f
C308 source.n122 a_n2762_n2088# 0.025293f
C309 source.n123 a_n2762_n2088# 0.01992f
C310 source.n124 a_n2762_n2088# 0.014268f
C311 source.n125 a_n2762_n2088# 0.631779f
C312 source.n126 a_n2762_n2088# 0.026552f
C313 source.n127 a_n2762_n2088# 0.014268f
C314 source.n128 a_n2762_n2088# 0.015107f
C315 source.n129 a_n2762_n2088# 0.033724f
C316 source.n130 a_n2762_n2088# 0.033724f
C317 source.n131 a_n2762_n2088# 0.015107f
C318 source.n132 a_n2762_n2088# 0.014268f
C319 source.n133 a_n2762_n2088# 0.026552f
C320 source.n134 a_n2762_n2088# 0.026552f
C321 source.n135 a_n2762_n2088# 0.014268f
C322 source.n136 a_n2762_n2088# 0.015107f
C323 source.n137 a_n2762_n2088# 0.033724f
C324 source.n138 a_n2762_n2088# 0.073007f
C325 source.n139 a_n2762_n2088# 0.015107f
C326 source.n140 a_n2762_n2088# 0.014268f
C327 source.n141 a_n2762_n2088# 0.061374f
C328 source.n142 a_n2762_n2088# 0.04085f
C329 source.n143 a_n2762_n2088# 1.02922f
C330 source.n144 a_n2762_n2088# 0.037321f
C331 source.n145 a_n2762_n2088# 0.026552f
C332 source.n146 a_n2762_n2088# 0.014268f
C333 source.n147 a_n2762_n2088# 0.033724f
C334 source.n148 a_n2762_n2088# 0.015107f
C335 source.n149 a_n2762_n2088# 0.026552f
C336 source.n150 a_n2762_n2088# 0.014268f
C337 source.n151 a_n2762_n2088# 0.033724f
C338 source.n152 a_n2762_n2088# 0.015107f
C339 source.n153 a_n2762_n2088# 0.113624f
C340 source.t22 a_n2762_n2088# 0.054966f
C341 source.n154 a_n2762_n2088# 0.025293f
C342 source.n155 a_n2762_n2088# 0.01992f
C343 source.n156 a_n2762_n2088# 0.014268f
C344 source.n157 a_n2762_n2088# 0.631779f
C345 source.n158 a_n2762_n2088# 0.026552f
C346 source.n159 a_n2762_n2088# 0.014268f
C347 source.n160 a_n2762_n2088# 0.015107f
C348 source.n161 a_n2762_n2088# 0.033724f
C349 source.n162 a_n2762_n2088# 0.033724f
C350 source.n163 a_n2762_n2088# 0.015107f
C351 source.n164 a_n2762_n2088# 0.014268f
C352 source.n165 a_n2762_n2088# 0.026552f
C353 source.n166 a_n2762_n2088# 0.026552f
C354 source.n167 a_n2762_n2088# 0.014268f
C355 source.n168 a_n2762_n2088# 0.015107f
C356 source.n169 a_n2762_n2088# 0.033724f
C357 source.n170 a_n2762_n2088# 0.073007f
C358 source.n171 a_n2762_n2088# 0.015107f
C359 source.n172 a_n2762_n2088# 0.014268f
C360 source.n173 a_n2762_n2088# 0.061374f
C361 source.n174 a_n2762_n2088# 0.04085f
C362 source.n175 a_n2762_n2088# 1.02922f
C363 source.t24 a_n2762_n2088# 0.125893f
C364 source.t20 a_n2762_n2088# 0.125893f
C365 source.n176 a_n2762_n2088# 0.980459f
C366 source.n177 a_n2762_n2088# 0.386091f
C367 source.t27 a_n2762_n2088# 0.125893f
C368 source.t31 a_n2762_n2088# 0.125893f
C369 source.n178 a_n2762_n2088# 0.980459f
C370 source.n179 a_n2762_n2088# 0.386091f
C371 source.t25 a_n2762_n2088# 0.125893f
C372 source.t39 a_n2762_n2088# 0.125893f
C373 source.n180 a_n2762_n2088# 0.980459f
C374 source.n181 a_n2762_n2088# 0.386091f
C375 source.t28 a_n2762_n2088# 0.125893f
C376 source.t32 a_n2762_n2088# 0.125893f
C377 source.n182 a_n2762_n2088# 0.980459f
C378 source.n183 a_n2762_n2088# 0.386091f
C379 source.n184 a_n2762_n2088# 0.037321f
C380 source.n185 a_n2762_n2088# 0.026552f
C381 source.n186 a_n2762_n2088# 0.014268f
C382 source.n187 a_n2762_n2088# 0.033724f
C383 source.n188 a_n2762_n2088# 0.015107f
C384 source.n189 a_n2762_n2088# 0.026552f
C385 source.n190 a_n2762_n2088# 0.014268f
C386 source.n191 a_n2762_n2088# 0.033724f
C387 source.n192 a_n2762_n2088# 0.015107f
C388 source.n193 a_n2762_n2088# 0.113624f
C389 source.t33 a_n2762_n2088# 0.054966f
C390 source.n194 a_n2762_n2088# 0.025293f
C391 source.n195 a_n2762_n2088# 0.01992f
C392 source.n196 a_n2762_n2088# 0.014268f
C393 source.n197 a_n2762_n2088# 0.631779f
C394 source.n198 a_n2762_n2088# 0.026552f
C395 source.n199 a_n2762_n2088# 0.014268f
C396 source.n200 a_n2762_n2088# 0.015107f
C397 source.n201 a_n2762_n2088# 0.033724f
C398 source.n202 a_n2762_n2088# 0.033724f
C399 source.n203 a_n2762_n2088# 0.015107f
C400 source.n204 a_n2762_n2088# 0.014268f
C401 source.n205 a_n2762_n2088# 0.026552f
C402 source.n206 a_n2762_n2088# 0.026552f
C403 source.n207 a_n2762_n2088# 0.014268f
C404 source.n208 a_n2762_n2088# 0.015107f
C405 source.n209 a_n2762_n2088# 0.033724f
C406 source.n210 a_n2762_n2088# 0.073007f
C407 source.n211 a_n2762_n2088# 0.015107f
C408 source.n212 a_n2762_n2088# 0.014268f
C409 source.n213 a_n2762_n2088# 0.061374f
C410 source.n214 a_n2762_n2088# 0.04085f
C411 source.n215 a_n2762_n2088# 0.131467f
C412 source.n216 a_n2762_n2088# 0.037321f
C413 source.n217 a_n2762_n2088# 0.026552f
C414 source.n218 a_n2762_n2088# 0.014268f
C415 source.n219 a_n2762_n2088# 0.033724f
C416 source.n220 a_n2762_n2088# 0.015107f
C417 source.n221 a_n2762_n2088# 0.026552f
C418 source.n222 a_n2762_n2088# 0.014268f
C419 source.n223 a_n2762_n2088# 0.033724f
C420 source.n224 a_n2762_n2088# 0.015107f
C421 source.n225 a_n2762_n2088# 0.113624f
C422 source.t5 a_n2762_n2088# 0.054966f
C423 source.n226 a_n2762_n2088# 0.025293f
C424 source.n227 a_n2762_n2088# 0.01992f
C425 source.n228 a_n2762_n2088# 0.014268f
C426 source.n229 a_n2762_n2088# 0.631779f
C427 source.n230 a_n2762_n2088# 0.026552f
C428 source.n231 a_n2762_n2088# 0.014268f
C429 source.n232 a_n2762_n2088# 0.015107f
C430 source.n233 a_n2762_n2088# 0.033724f
C431 source.n234 a_n2762_n2088# 0.033724f
C432 source.n235 a_n2762_n2088# 0.015107f
C433 source.n236 a_n2762_n2088# 0.014268f
C434 source.n237 a_n2762_n2088# 0.026552f
C435 source.n238 a_n2762_n2088# 0.026552f
C436 source.n239 a_n2762_n2088# 0.014268f
C437 source.n240 a_n2762_n2088# 0.015107f
C438 source.n241 a_n2762_n2088# 0.033724f
C439 source.n242 a_n2762_n2088# 0.073007f
C440 source.n243 a_n2762_n2088# 0.015107f
C441 source.n244 a_n2762_n2088# 0.014268f
C442 source.n245 a_n2762_n2088# 0.061374f
C443 source.n246 a_n2762_n2088# 0.04085f
C444 source.n247 a_n2762_n2088# 0.131467f
C445 source.t11 a_n2762_n2088# 0.125893f
C446 source.t6 a_n2762_n2088# 0.125893f
C447 source.n248 a_n2762_n2088# 0.980459f
C448 source.n249 a_n2762_n2088# 0.386091f
C449 source.t15 a_n2762_n2088# 0.125893f
C450 source.t7 a_n2762_n2088# 0.125893f
C451 source.n250 a_n2762_n2088# 0.980459f
C452 source.n251 a_n2762_n2088# 0.386091f
C453 source.t14 a_n2762_n2088# 0.125893f
C454 source.t9 a_n2762_n2088# 0.125893f
C455 source.n252 a_n2762_n2088# 0.980459f
C456 source.n253 a_n2762_n2088# 0.386091f
C457 source.t16 a_n2762_n2088# 0.125893f
C458 source.t18 a_n2762_n2088# 0.125893f
C459 source.n254 a_n2762_n2088# 0.980459f
C460 source.n255 a_n2762_n2088# 0.386091f
C461 source.n256 a_n2762_n2088# 0.037321f
C462 source.n257 a_n2762_n2088# 0.026552f
C463 source.n258 a_n2762_n2088# 0.014268f
C464 source.n259 a_n2762_n2088# 0.033724f
C465 source.n260 a_n2762_n2088# 0.015107f
C466 source.n261 a_n2762_n2088# 0.026552f
C467 source.n262 a_n2762_n2088# 0.014268f
C468 source.n263 a_n2762_n2088# 0.033724f
C469 source.n264 a_n2762_n2088# 0.015107f
C470 source.n265 a_n2762_n2088# 0.113624f
C471 source.t12 a_n2762_n2088# 0.054966f
C472 source.n266 a_n2762_n2088# 0.025293f
C473 source.n267 a_n2762_n2088# 0.01992f
C474 source.n268 a_n2762_n2088# 0.014268f
C475 source.n269 a_n2762_n2088# 0.631779f
C476 source.n270 a_n2762_n2088# 0.026552f
C477 source.n271 a_n2762_n2088# 0.014268f
C478 source.n272 a_n2762_n2088# 0.015107f
C479 source.n273 a_n2762_n2088# 0.033724f
C480 source.n274 a_n2762_n2088# 0.033724f
C481 source.n275 a_n2762_n2088# 0.015107f
C482 source.n276 a_n2762_n2088# 0.014268f
C483 source.n277 a_n2762_n2088# 0.026552f
C484 source.n278 a_n2762_n2088# 0.026552f
C485 source.n279 a_n2762_n2088# 0.014268f
C486 source.n280 a_n2762_n2088# 0.015107f
C487 source.n281 a_n2762_n2088# 0.033724f
C488 source.n282 a_n2762_n2088# 0.073007f
C489 source.n283 a_n2762_n2088# 0.015107f
C490 source.n284 a_n2762_n2088# 0.014268f
C491 source.n285 a_n2762_n2088# 0.061374f
C492 source.n286 a_n2762_n2088# 0.04085f
C493 source.n287 a_n2762_n2088# 0.298887f
C494 source.n288 a_n2762_n2088# 1.09742f
C495 plus.n0 a_n2762_n2088# 0.057909f
C496 plus.t0 a_n2762_n2088# 0.454222f
C497 plus.t2 a_n2762_n2088# 0.454222f
C498 plus.t3 a_n2762_n2088# 0.454222f
C499 plus.n1 a_n2762_n2088# 0.058045f
C500 plus.t4 a_n2762_n2088# 0.454222f
C501 plus.n2 a_n2762_n2088# 0.213869f
C502 plus.n3 a_n2762_n2088# 0.043499f
C503 plus.t5 a_n2762_n2088# 0.454222f
C504 plus.t9 a_n2762_n2088# 0.454222f
C505 plus.n4 a_n2762_n2088# 0.213869f
C506 plus.n5 a_n2762_n2088# 0.043499f
C507 plus.t13 a_n2762_n2088# 0.454222f
C508 plus.t14 a_n2762_n2088# 0.454222f
C509 plus.n6 a_n2762_n2088# 0.212662f
C510 plus.t15 a_n2762_n2088# 0.454222f
C511 plus.n7 a_n2762_n2088# 0.221862f
C512 plus.t16 a_n2762_n2088# 0.471292f
C513 plus.n8 a_n2762_n2088# 0.195856f
C514 plus.n9 a_n2762_n2088# 0.185669f
C515 plus.n10 a_n2762_n2088# 0.043499f
C516 plus.n11 a_n2762_n2088# 0.009871f
C517 plus.n12 a_n2762_n2088# 0.213869f
C518 plus.n13 a_n2762_n2088# 0.009871f
C519 plus.n14 a_n2762_n2088# 0.043499f
C520 plus.n15 a_n2762_n2088# 0.043499f
C521 plus.n16 a_n2762_n2088# 0.043499f
C522 plus.n17 a_n2762_n2088# 0.009871f
C523 plus.n18 a_n2762_n2088# 0.213869f
C524 plus.n19 a_n2762_n2088# 0.009871f
C525 plus.n20 a_n2762_n2088# 0.043499f
C526 plus.n21 a_n2762_n2088# 0.043499f
C527 plus.n22 a_n2762_n2088# 0.043499f
C528 plus.n23 a_n2762_n2088# 0.009871f
C529 plus.n24 a_n2762_n2088# 0.212662f
C530 plus.n25 a_n2762_n2088# 0.221862f
C531 plus.n26 a_n2762_n2088# 0.211991f
C532 plus.n27 a_n2762_n2088# 0.40105f
C533 plus.n28 a_n2762_n2088# 0.057909f
C534 plus.t8 a_n2762_n2088# 0.454222f
C535 plus.t19 a_n2762_n2088# 0.454222f
C536 plus.n29 a_n2762_n2088# 0.058045f
C537 plus.t12 a_n2762_n2088# 0.454222f
C538 plus.t7 a_n2762_n2088# 0.454222f
C539 plus.n30 a_n2762_n2088# 0.213869f
C540 plus.n31 a_n2762_n2088# 0.043499f
C541 plus.t18 a_n2762_n2088# 0.454222f
C542 plus.t17 a_n2762_n2088# 0.454222f
C543 plus.n32 a_n2762_n2088# 0.213869f
C544 plus.n33 a_n2762_n2088# 0.043499f
C545 plus.t11 a_n2762_n2088# 0.454222f
C546 plus.t6 a_n2762_n2088# 0.454222f
C547 plus.n34 a_n2762_n2088# 0.212662f
C548 plus.t1 a_n2762_n2088# 0.454222f
C549 plus.n35 a_n2762_n2088# 0.221862f
C550 plus.t10 a_n2762_n2088# 0.471292f
C551 plus.n36 a_n2762_n2088# 0.195856f
C552 plus.n37 a_n2762_n2088# 0.185669f
C553 plus.n38 a_n2762_n2088# 0.043499f
C554 plus.n39 a_n2762_n2088# 0.009871f
C555 plus.n40 a_n2762_n2088# 0.213869f
C556 plus.n41 a_n2762_n2088# 0.009871f
C557 plus.n42 a_n2762_n2088# 0.043499f
C558 plus.n43 a_n2762_n2088# 0.043499f
C559 plus.n44 a_n2762_n2088# 0.043499f
C560 plus.n45 a_n2762_n2088# 0.009871f
C561 plus.n46 a_n2762_n2088# 0.213869f
C562 plus.n47 a_n2762_n2088# 0.009871f
C563 plus.n48 a_n2762_n2088# 0.043499f
C564 plus.n49 a_n2762_n2088# 0.043499f
C565 plus.n50 a_n2762_n2088# 0.043499f
C566 plus.n51 a_n2762_n2088# 0.009871f
C567 plus.n52 a_n2762_n2088# 0.212662f
C568 plus.n53 a_n2762_n2088# 0.221862f
C569 plus.n54 a_n2762_n2088# 0.211991f
C570 plus.n55 a_n2762_n2088# 1.34975f
.ends

