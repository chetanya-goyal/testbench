* NGSPICE file created from diffpair220.ext - technology: sky130A

.subckt diffpair220 minus drain_right drain_left source plus
X0 drain_right minus source a_n1128_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=0.7
X1 drain_right minus source a_n1128_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=0.7
X2 a_n1128_n1492# a_n1128_n1492# a_n1128_n1492# a_n1128_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.7
X3 a_n1128_n1492# a_n1128_n1492# a_n1128_n1492# a_n1128_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X4 drain_left plus source a_n1128_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=0.7
X5 a_n1128_n1492# a_n1128_n1492# a_n1128_n1492# a_n1128_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X6 drain_left plus source a_n1128_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=0.7
X7 a_n1128_n1492# a_n1128_n1492# a_n1128_n1492# a_n1128_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
.ends

