* NGSPICE file created from diffpair335.ext - technology: sky130A

.subckt diffpair335 minus drain_right drain_left source plus
X0 source.t23 minus.t0 drain_right.t4 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X1 source.t22 minus.t1 drain_right.t11 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X2 drain_right.t8 minus.t2 source.t21 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X3 drain_right.t3 minus.t3 source.t20 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X4 drain_right.t9 minus.t4 source.t19 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X5 a_n1458_n2688# a_n1458_n2688# a_n1458_n2688# a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.2
X6 drain_right.t0 minus.t5 source.t18 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X7 drain_left.t11 plus.t0 source.t10 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X8 source.t17 minus.t6 drain_right.t6 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X9 source.t16 minus.t7 drain_right.t10 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X10 source.t15 minus.t8 drain_right.t7 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X11 drain_left.t10 plus.t1 source.t1 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X12 source.t5 plus.t2 drain_left.t9 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X13 source.t8 plus.t3 drain_left.t8 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X14 source.t4 plus.t4 drain_left.t7 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X15 a_n1458_n2688# a_n1458_n2688# a_n1458_n2688# a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X16 drain_right.t5 minus.t9 source.t14 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X17 drain_right.t2 minus.t10 source.t13 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X18 a_n1458_n2688# a_n1458_n2688# a_n1458_n2688# a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X19 drain_left.t6 plus.t5 source.t6 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X20 drain_left.t5 plus.t6 source.t11 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X21 drain_left.t4 plus.t7 source.t3 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X22 a_n1458_n2688# a_n1458_n2688# a_n1458_n2688# a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X23 source.t7 plus.t8 drain_left.t3 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X24 drain_left.t2 plus.t9 source.t9 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X25 source.t0 plus.t10 drain_left.t1 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X26 source.t12 minus.t11 drain_right.t1 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
X27 source.t2 plus.t11 drain_left.t0 a_n1458_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.2
R0 minus.n11 minus.t7 1288.62
R1 minus.n2 minus.t9 1288.62
R2 minus.n24 minus.t5 1288.62
R3 minus.n15 minus.t1 1288.62
R4 minus.n10 minus.t10 1241.15
R5 minus.n8 minus.t11 1241.15
R6 minus.n1 minus.t2 1241.15
R7 minus.n3 minus.t8 1241.15
R8 minus.n23 minus.t6 1241.15
R9 minus.n21 minus.t3 1241.15
R10 minus.n14 minus.t0 1241.15
R11 minus.n16 minus.t4 1241.15
R12 minus.n5 minus.n2 161.489
R13 minus.n18 minus.n15 161.489
R14 minus.n12 minus.n11 161.3
R15 minus.n9 minus.n0 161.3
R16 minus.n7 minus.n6 161.3
R17 minus.n5 minus.n4 161.3
R18 minus.n25 minus.n24 161.3
R19 minus.n22 minus.n13 161.3
R20 minus.n20 minus.n19 161.3
R21 minus.n18 minus.n17 161.3
R22 minus.n10 minus.n9 43.0884
R23 minus.n4 minus.n3 43.0884
R24 minus.n17 minus.n16 43.0884
R25 minus.n23 minus.n22 43.0884
R26 minus.n8 minus.n7 38.7066
R27 minus.n7 minus.n1 38.7066
R28 minus.n20 minus.n14 38.7066
R29 minus.n21 minus.n20 38.7066
R30 minus.n9 minus.n8 34.3247
R31 minus.n4 minus.n1 34.3247
R32 minus.n17 minus.n14 34.3247
R33 minus.n22 minus.n21 34.3247
R34 minus.n26 minus.n12 32.3263
R35 minus.n11 minus.n10 29.9429
R36 minus.n3 minus.n2 29.9429
R37 minus.n16 minus.n15 29.9429
R38 minus.n24 minus.n23 29.9429
R39 minus.n26 minus.n25 6.45505
R40 minus.n12 minus.n0 0.189894
R41 minus.n6 minus.n0 0.189894
R42 minus.n6 minus.n5 0.189894
R43 minus.n19 minus.n18 0.189894
R44 minus.n19 minus.n13 0.189894
R45 minus.n25 minus.n13 0.189894
R46 minus minus.n26 0.188
R47 drain_right.n6 drain_right.n4 65.9943
R48 drain_right.n3 drain_right.n2 65.9389
R49 drain_right.n3 drain_right.n0 65.9389
R50 drain_right.n6 drain_right.n5 65.5376
R51 drain_right.n8 drain_right.n7 65.5376
R52 drain_right.n3 drain_right.n1 65.5373
R53 drain_right drain_right.n3 26.8256
R54 drain_right drain_right.n8 6.11011
R55 drain_right.n1 drain_right.t4 2.2005
R56 drain_right.n1 drain_right.t3 2.2005
R57 drain_right.n2 drain_right.t6 2.2005
R58 drain_right.n2 drain_right.t0 2.2005
R59 drain_right.n0 drain_right.t11 2.2005
R60 drain_right.n0 drain_right.t9 2.2005
R61 drain_right.n4 drain_right.t7 2.2005
R62 drain_right.n4 drain_right.t5 2.2005
R63 drain_right.n5 drain_right.t1 2.2005
R64 drain_right.n5 drain_right.t8 2.2005
R65 drain_right.n7 drain_right.t10 2.2005
R66 drain_right.n7 drain_right.t2 2.2005
R67 drain_right.n8 drain_right.n6 0.457397
R68 source.n5 source.t5 51.0588
R69 source.n6 source.t14 51.0588
R70 source.n11 source.t16 51.0588
R71 source.n23 source.t18 51.0586
R72 source.n18 source.t22 51.0586
R73 source.n17 source.t11 51.0586
R74 source.n12 source.t4 51.0586
R75 source.n0 source.t1 51.0586
R76 source.n2 source.n1 48.8588
R77 source.n4 source.n3 48.8588
R78 source.n8 source.n7 48.8588
R79 source.n10 source.n9 48.8588
R80 source.n22 source.n21 48.8586
R81 source.n20 source.n19 48.8586
R82 source.n16 source.n15 48.8586
R83 source.n14 source.n13 48.8586
R84 source.n12 source.n11 19.4719
R85 source.n24 source.n0 13.9805
R86 source.n24 source.n23 5.49188
R87 source.n21 source.t20 2.2005
R88 source.n21 source.t17 2.2005
R89 source.n19 source.t19 2.2005
R90 source.n19 source.t23 2.2005
R91 source.n15 source.t3 2.2005
R92 source.n15 source.t0 2.2005
R93 source.n13 source.t6 2.2005
R94 source.n13 source.t8 2.2005
R95 source.n1 source.t9 2.2005
R96 source.n1 source.t7 2.2005
R97 source.n3 source.t10 2.2005
R98 source.n3 source.t2 2.2005
R99 source.n7 source.t21 2.2005
R100 source.n7 source.t15 2.2005
R101 source.n9 source.t13 2.2005
R102 source.n9 source.t12 2.2005
R103 source.n6 source.n5 0.470328
R104 source.n18 source.n17 0.470328
R105 source.n11 source.n10 0.457397
R106 source.n10 source.n8 0.457397
R107 source.n8 source.n6 0.457397
R108 source.n5 source.n4 0.457397
R109 source.n4 source.n2 0.457397
R110 source.n2 source.n0 0.457397
R111 source.n14 source.n12 0.457397
R112 source.n16 source.n14 0.457397
R113 source.n17 source.n16 0.457397
R114 source.n20 source.n18 0.457397
R115 source.n22 source.n20 0.457397
R116 source.n23 source.n22 0.457397
R117 source source.n24 0.188
R118 plus.n2 plus.t2 1288.62
R119 plus.n11 plus.t1 1288.62
R120 plus.n15 plus.t6 1288.62
R121 plus.n24 plus.t4 1288.62
R122 plus.n3 plus.t0 1241.15
R123 plus.n1 plus.t11 1241.15
R124 plus.n8 plus.t9 1241.15
R125 plus.n10 plus.t8 1241.15
R126 plus.n16 plus.t10 1241.15
R127 plus.n14 plus.t7 1241.15
R128 plus.n21 plus.t3 1241.15
R129 plus.n23 plus.t5 1241.15
R130 plus.n5 plus.n2 161.489
R131 plus.n18 plus.n15 161.489
R132 plus.n5 plus.n4 161.3
R133 plus.n7 plus.n6 161.3
R134 plus.n9 plus.n0 161.3
R135 plus.n12 plus.n11 161.3
R136 plus.n18 plus.n17 161.3
R137 plus.n20 plus.n19 161.3
R138 plus.n22 plus.n13 161.3
R139 plus.n25 plus.n24 161.3
R140 plus.n4 plus.n3 43.0884
R141 plus.n10 plus.n9 43.0884
R142 plus.n23 plus.n22 43.0884
R143 plus.n17 plus.n16 43.0884
R144 plus.n7 plus.n1 38.7066
R145 plus.n8 plus.n7 38.7066
R146 plus.n21 plus.n20 38.7066
R147 plus.n20 plus.n14 38.7066
R148 plus.n4 plus.n1 34.3247
R149 plus.n9 plus.n8 34.3247
R150 plus.n22 plus.n21 34.3247
R151 plus.n17 plus.n14 34.3247
R152 plus.n3 plus.n2 29.9429
R153 plus.n11 plus.n10 29.9429
R154 plus.n24 plus.n23 29.9429
R155 plus.n16 plus.n15 29.9429
R156 plus plus.n25 27.3437
R157 plus plus.n12 10.9626
R158 plus.n6 plus.n5 0.189894
R159 plus.n6 plus.n0 0.189894
R160 plus.n12 plus.n0 0.189894
R161 plus.n25 plus.n13 0.189894
R162 plus.n19 plus.n13 0.189894
R163 plus.n19 plus.n18 0.189894
R164 drain_left.n6 drain_left.n4 65.9945
R165 drain_left.n3 drain_left.n2 65.9389
R166 drain_left.n3 drain_left.n0 65.9389
R167 drain_left.n6 drain_left.n5 65.5376
R168 drain_left.n8 drain_left.n7 65.5374
R169 drain_left.n3 drain_left.n1 65.5373
R170 drain_left drain_left.n3 27.3788
R171 drain_left drain_left.n8 6.11011
R172 drain_left.n1 drain_left.t8 2.2005
R173 drain_left.n1 drain_left.t4 2.2005
R174 drain_left.n2 drain_left.t1 2.2005
R175 drain_left.n2 drain_left.t5 2.2005
R176 drain_left.n0 drain_left.t7 2.2005
R177 drain_left.n0 drain_left.t6 2.2005
R178 drain_left.n7 drain_left.t3 2.2005
R179 drain_left.n7 drain_left.t10 2.2005
R180 drain_left.n5 drain_left.t0 2.2005
R181 drain_left.n5 drain_left.t2 2.2005
R182 drain_left.n4 drain_left.t9 2.2005
R183 drain_left.n4 drain_left.t11 2.2005
R184 drain_left.n8 drain_left.n6 0.457397
C0 plus minus 4.41722f
C1 plus drain_left 2.88872f
C2 drain_left minus 0.17046f
C3 source drain_right 21.6828f
C4 plus drain_right 0.292203f
C5 drain_right minus 2.74984f
C6 drain_left drain_right 0.711832f
C7 plus source 2.44333f
C8 source minus 2.42929f
C9 source drain_left 21.683699f
C10 drain_right a_n1458_n2688# 5.65497f
C11 drain_left a_n1458_n2688# 5.90442f
C12 source a_n1458_n2688# 6.849774f
C13 minus a_n1458_n2688# 5.430179f
C14 plus a_n1458_n2688# 7.26515f
C15 drain_left.t7 a_n1458_n2688# 0.268206f
C16 drain_left.t6 a_n1458_n2688# 0.268206f
C17 drain_left.n0 a_n1458_n2688# 2.34849f
C18 drain_left.t8 a_n1458_n2688# 0.268206f
C19 drain_left.t4 a_n1458_n2688# 0.268206f
C20 drain_left.n1 a_n1458_n2688# 2.34591f
C21 drain_left.t1 a_n1458_n2688# 0.268206f
C22 drain_left.t5 a_n1458_n2688# 0.268206f
C23 drain_left.n2 a_n1458_n2688# 2.34849f
C24 drain_left.n3 a_n1458_n2688# 2.63701f
C25 drain_left.t9 a_n1458_n2688# 0.268206f
C26 drain_left.t11 a_n1458_n2688# 0.268206f
C27 drain_left.n4 a_n1458_n2688# 2.34888f
C28 drain_left.t0 a_n1458_n2688# 0.268206f
C29 drain_left.t2 a_n1458_n2688# 0.268206f
C30 drain_left.n5 a_n1458_n2688# 2.34591f
C31 drain_left.n6 a_n1458_n2688# 0.838439f
C32 drain_left.t3 a_n1458_n2688# 0.268206f
C33 drain_left.t10 a_n1458_n2688# 0.268206f
C34 drain_left.n7 a_n1458_n2688# 2.3459f
C35 drain_left.n8 a_n1458_n2688# 0.72175f
C36 plus.n0 a_n1458_n2688# 0.056825f
C37 plus.t8 a_n1458_n2688# 0.289836f
C38 plus.t9 a_n1458_n2688# 0.289836f
C39 plus.t11 a_n1458_n2688# 0.289836f
C40 plus.n1 a_n1458_n2688# 0.12687f
C41 plus.t2 a_n1458_n2688# 0.294542f
C42 plus.n2 a_n1458_n2688# 0.143023f
C43 plus.t0 a_n1458_n2688# 0.289836f
C44 plus.n3 a_n1458_n2688# 0.12687f
C45 plus.n4 a_n1458_n2688# 0.019902f
C46 plus.n5 a_n1458_n2688# 0.125832f
C47 plus.n6 a_n1458_n2688# 0.056825f
C48 plus.n7 a_n1458_n2688# 0.019902f
C49 plus.n8 a_n1458_n2688# 0.12687f
C50 plus.n9 a_n1458_n2688# 0.019902f
C51 plus.n10 a_n1458_n2688# 0.12687f
C52 plus.t1 a_n1458_n2688# 0.294542f
C53 plus.n11 a_n1458_n2688# 0.142942f
C54 plus.n12 a_n1458_n2688# 0.551987f
C55 plus.n13 a_n1458_n2688# 0.056825f
C56 plus.t4 a_n1458_n2688# 0.294542f
C57 plus.t5 a_n1458_n2688# 0.289836f
C58 plus.t3 a_n1458_n2688# 0.289836f
C59 plus.t7 a_n1458_n2688# 0.289836f
C60 plus.n14 a_n1458_n2688# 0.12687f
C61 plus.t6 a_n1458_n2688# 0.294542f
C62 plus.n15 a_n1458_n2688# 0.143023f
C63 plus.t10 a_n1458_n2688# 0.289836f
C64 plus.n16 a_n1458_n2688# 0.12687f
C65 plus.n17 a_n1458_n2688# 0.019902f
C66 plus.n18 a_n1458_n2688# 0.125832f
C67 plus.n19 a_n1458_n2688# 0.056825f
C68 plus.n20 a_n1458_n2688# 0.019902f
C69 plus.n21 a_n1458_n2688# 0.12687f
C70 plus.n22 a_n1458_n2688# 0.019902f
C71 plus.n23 a_n1458_n2688# 0.12687f
C72 plus.n24 a_n1458_n2688# 0.142942f
C73 plus.n25 a_n1458_n2688# 1.45658f
C74 source.t1 a_n1458_n2688# 2.3001f
C75 source.n0 a_n1458_n2688# 1.30851f
C76 source.t9 a_n1458_n2688# 0.215699f
C77 source.t7 a_n1458_n2688# 0.215699f
C78 source.n1 a_n1458_n2688# 1.80569f
C79 source.n2 a_n1458_n2688# 0.371968f
C80 source.t10 a_n1458_n2688# 0.215699f
C81 source.t2 a_n1458_n2688# 0.215699f
C82 source.n3 a_n1458_n2688# 1.80569f
C83 source.n4 a_n1458_n2688# 0.371968f
C84 source.t5 a_n1458_n2688# 2.3001f
C85 source.n5 a_n1458_n2688# 0.467089f
C86 source.t14 a_n1458_n2688# 2.3001f
C87 source.n6 a_n1458_n2688# 0.467089f
C88 source.t21 a_n1458_n2688# 0.215699f
C89 source.t15 a_n1458_n2688# 0.215699f
C90 source.n7 a_n1458_n2688# 1.80569f
C91 source.n8 a_n1458_n2688# 0.371968f
C92 source.t13 a_n1458_n2688# 0.215699f
C93 source.t12 a_n1458_n2688# 0.215699f
C94 source.n9 a_n1458_n2688# 1.80569f
C95 source.n10 a_n1458_n2688# 0.371968f
C96 source.t16 a_n1458_n2688# 2.3001f
C97 source.n11 a_n1458_n2688# 1.74644f
C98 source.t4 a_n1458_n2688# 2.3001f
C99 source.n12 a_n1458_n2688# 1.74644f
C100 source.t6 a_n1458_n2688# 0.215699f
C101 source.t8 a_n1458_n2688# 0.215699f
C102 source.n13 a_n1458_n2688# 1.80568f
C103 source.n14 a_n1458_n2688# 0.371974f
C104 source.t3 a_n1458_n2688# 0.215699f
C105 source.t0 a_n1458_n2688# 0.215699f
C106 source.n15 a_n1458_n2688# 1.80568f
C107 source.n16 a_n1458_n2688# 0.371974f
C108 source.t11 a_n1458_n2688# 2.3001f
C109 source.n17 a_n1458_n2688# 0.467094f
C110 source.t22 a_n1458_n2688# 2.3001f
C111 source.n18 a_n1458_n2688# 0.467094f
C112 source.t19 a_n1458_n2688# 0.215699f
C113 source.t23 a_n1458_n2688# 0.215699f
C114 source.n19 a_n1458_n2688# 1.80568f
C115 source.n20 a_n1458_n2688# 0.371974f
C116 source.t20 a_n1458_n2688# 0.215699f
C117 source.t17 a_n1458_n2688# 0.215699f
C118 source.n21 a_n1458_n2688# 1.80568f
C119 source.n22 a_n1458_n2688# 0.371974f
C120 source.t18 a_n1458_n2688# 2.3001f
C121 source.n23 a_n1458_n2688# 0.631545f
C122 source.n24 a_n1458_n2688# 1.5744f
C123 drain_right.t11 a_n1458_n2688# 0.267631f
C124 drain_right.t9 a_n1458_n2688# 0.267631f
C125 drain_right.n0 a_n1458_n2688# 2.34345f
C126 drain_right.t4 a_n1458_n2688# 0.267631f
C127 drain_right.t3 a_n1458_n2688# 0.267631f
C128 drain_right.n1 a_n1458_n2688# 2.34088f
C129 drain_right.t6 a_n1458_n2688# 0.267631f
C130 drain_right.t0 a_n1458_n2688# 0.267631f
C131 drain_right.n2 a_n1458_n2688# 2.34345f
C132 drain_right.n3 a_n1458_n2688# 2.55334f
C133 drain_right.t7 a_n1458_n2688# 0.267631f
C134 drain_right.t5 a_n1458_n2688# 0.267631f
C135 drain_right.n4 a_n1458_n2688# 2.34383f
C136 drain_right.t1 a_n1458_n2688# 0.267631f
C137 drain_right.t8 a_n1458_n2688# 0.267631f
C138 drain_right.n5 a_n1458_n2688# 2.34088f
C139 drain_right.n6 a_n1458_n2688# 0.836649f
C140 drain_right.t10 a_n1458_n2688# 0.267631f
C141 drain_right.t2 a_n1458_n2688# 0.267631f
C142 drain_right.n7 a_n1458_n2688# 2.34088f
C143 drain_right.n8 a_n1458_n2688# 0.720191f
C144 minus.n0 a_n1458_n2688# 0.055002f
C145 minus.t7 a_n1458_n2688# 0.285092f
C146 minus.t10 a_n1458_n2688# 0.280537f
C147 minus.t11 a_n1458_n2688# 0.280537f
C148 minus.t2 a_n1458_n2688# 0.280537f
C149 minus.n1 a_n1458_n2688# 0.122799f
C150 minus.t9 a_n1458_n2688# 0.285092f
C151 minus.n2 a_n1458_n2688# 0.138434f
C152 minus.t8 a_n1458_n2688# 0.280537f
C153 minus.n3 a_n1458_n2688# 0.122799f
C154 minus.n4 a_n1458_n2688# 0.019263f
C155 minus.n5 a_n1458_n2688# 0.121794f
C156 minus.n6 a_n1458_n2688# 0.055002f
C157 minus.n7 a_n1458_n2688# 0.019263f
C158 minus.n8 a_n1458_n2688# 0.122799f
C159 minus.n9 a_n1458_n2688# 0.019263f
C160 minus.n10 a_n1458_n2688# 0.122799f
C161 minus.n11 a_n1458_n2688# 0.138355f
C162 minus.n12 a_n1458_n2688# 1.6195f
C163 minus.n13 a_n1458_n2688# 0.055002f
C164 minus.t6 a_n1458_n2688# 0.280537f
C165 minus.t3 a_n1458_n2688# 0.280537f
C166 minus.t0 a_n1458_n2688# 0.280537f
C167 minus.n14 a_n1458_n2688# 0.122799f
C168 minus.t1 a_n1458_n2688# 0.285092f
C169 minus.n15 a_n1458_n2688# 0.138434f
C170 minus.t4 a_n1458_n2688# 0.280537f
C171 minus.n16 a_n1458_n2688# 0.122799f
C172 minus.n17 a_n1458_n2688# 0.019263f
C173 minus.n18 a_n1458_n2688# 0.121794f
C174 minus.n19 a_n1458_n2688# 0.055002f
C175 minus.n20 a_n1458_n2688# 0.019263f
C176 minus.n21 a_n1458_n2688# 0.122799f
C177 minus.n22 a_n1458_n2688# 0.019263f
C178 minus.n23 a_n1458_n2688# 0.122799f
C179 minus.t5 a_n1458_n2688# 0.285092f
C180 minus.n24 a_n1458_n2688# 0.138355f
C181 minus.n25 a_n1458_n2688# 0.35375f
C182 minus.n26 a_n1458_n2688# 1.99082f
.ends

