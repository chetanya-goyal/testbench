* NGSPICE file created from diffpair513.ext - technology: sky130A

.subckt diffpair513 minus drain_right drain_left source plus
X0 drain_left.t7 plus.t0 source.t9 a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X1 drain_left.t6 plus.t1 source.t11 a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X2 drain_right.t7 minus.t0 source.t0 a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X3 source.t8 plus.t2 drain_left.t5 a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X4 source.t7 minus.t1 drain_right.t6 a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X5 source.t2 minus.t2 drain_right.t5 a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X6 a_n1346_n3888# a_n1346_n3888# a_n1346_n3888# a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.3
X7 a_n1346_n3888# a_n1346_n3888# a_n1346_n3888# a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X8 drain_left.t4 plus.t3 source.t13 a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X9 a_n1346_n3888# a_n1346_n3888# a_n1346_n3888# a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X10 source.t3 minus.t3 drain_right.t4 a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X11 drain_right.t3 minus.t4 source.t5 a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X12 source.t10 plus.t4 drain_left.t3 a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X13 source.t14 plus.t5 drain_left.t2 a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X14 source.t15 plus.t6 drain_left.t1 a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.3
X15 drain_right.t2 minus.t5 source.t1 a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
X16 drain_right.t1 minus.t6 source.t6 a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X17 source.t4 minus.t7 drain_right.t0 a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.3
X18 a_n1346_n3888# a_n1346_n3888# a_n1346_n3888# a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.3
X19 drain_left.t0 plus.t7 source.t12 a_n1346_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.3
R0 plus.n2 plus.t2 1337.92
R1 plus.n7 plus.t7 1337.92
R2 plus.n11 plus.t0 1337.92
R3 plus.n16 plus.t6 1337.92
R4 plus.n1 plus.t3 1309.43
R5 plus.n6 plus.t5 1309.43
R6 plus.n10 plus.t4 1309.43
R7 plus.n15 plus.t1 1309.43
R8 plus.n3 plus.n2 161.489
R9 plus.n12 plus.n11 161.489
R10 plus.n4 plus.n3 161.3
R11 plus.n5 plus.n0 161.3
R12 plus.n8 plus.n7 161.3
R13 plus.n13 plus.n12 161.3
R14 plus.n14 plus.n9 161.3
R15 plus.n17 plus.n16 161.3
R16 plus.n5 plus.n4 73.0308
R17 plus.n14 plus.n13 73.0308
R18 plus.n2 plus.n1 63.5369
R19 plus.n7 plus.n6 63.5369
R20 plus.n16 plus.n15 63.5369
R21 plus.n11 plus.n10 63.5369
R22 plus plus.n17 29.1998
R23 plus plus.n8 13.2429
R24 plus.n4 plus.n1 9.49444
R25 plus.n6 plus.n5 9.49444
R26 plus.n15 plus.n14 9.49444
R27 plus.n13 plus.n10 9.49444
R28 plus.n3 plus.n0 0.189894
R29 plus.n8 plus.n0 0.189894
R30 plus.n17 plus.n9 0.189894
R31 plus.n12 plus.n9 0.189894
R32 source.n3 source.t8 45.521
R33 source.n4 source.t5 45.521
R34 source.n7 source.t3 45.521
R35 source.n15 source.t1 45.5208
R36 source.n12 source.t2 45.5208
R37 source.n11 source.t9 45.5208
R38 source.n8 source.t15 45.5208
R39 source.n0 source.t12 45.5208
R40 source.n2 source.n1 44.201
R41 source.n6 source.n5 44.201
R42 source.n14 source.n13 44.2008
R43 source.n10 source.n9 44.2008
R44 source.n8 source.n7 24.1036
R45 source.n16 source.n0 18.5691
R46 source.n16 source.n15 5.53498
R47 source.n13 source.t6 1.3205
R48 source.n13 source.t7 1.3205
R49 source.n9 source.t11 1.3205
R50 source.n9 source.t10 1.3205
R51 source.n1 source.t13 1.3205
R52 source.n1 source.t14 1.3205
R53 source.n5 source.t0 1.3205
R54 source.n5 source.t4 1.3205
R55 source.n7 source.n6 0.543603
R56 source.n6 source.n4 0.543603
R57 source.n3 source.n2 0.543603
R58 source.n2 source.n0 0.543603
R59 source.n10 source.n8 0.543603
R60 source.n11 source.n10 0.543603
R61 source.n14 source.n12 0.543603
R62 source.n15 source.n14 0.543603
R63 source.n4 source.n3 0.470328
R64 source.n12 source.n11 0.470328
R65 source source.n16 0.188
R66 drain_left.n5 drain_left.n3 61.4229
R67 drain_left.n2 drain_left.n1 61.0958
R68 drain_left.n2 drain_left.n0 61.0958
R69 drain_left.n5 drain_left.n4 60.8796
R70 drain_left drain_left.n2 31.5407
R71 drain_left drain_left.n5 6.19632
R72 drain_left.n1 drain_left.t3 1.3205
R73 drain_left.n1 drain_left.t7 1.3205
R74 drain_left.n0 drain_left.t1 1.3205
R75 drain_left.n0 drain_left.t6 1.3205
R76 drain_left.n4 drain_left.t2 1.3205
R77 drain_left.n4 drain_left.t0 1.3205
R78 drain_left.n3 drain_left.t5 1.3205
R79 drain_left.n3 drain_left.t4 1.3205
R80 minus.n7 minus.t3 1337.92
R81 minus.n2 minus.t4 1337.92
R82 minus.n16 minus.t5 1337.92
R83 minus.n11 minus.t2 1337.92
R84 minus.n6 minus.t0 1309.43
R85 minus.n1 minus.t7 1309.43
R86 minus.n15 minus.t1 1309.43
R87 minus.n10 minus.t6 1309.43
R88 minus.n3 minus.n2 161.489
R89 minus.n12 minus.n11 161.489
R90 minus.n8 minus.n7 161.3
R91 minus.n5 minus.n0 161.3
R92 minus.n4 minus.n3 161.3
R93 minus.n17 minus.n16 161.3
R94 minus.n14 minus.n9 161.3
R95 minus.n13 minus.n12 161.3
R96 minus.n5 minus.n4 73.0308
R97 minus.n14 minus.n13 73.0308
R98 minus.n7 minus.n6 63.5369
R99 minus.n2 minus.n1 63.5369
R100 minus.n11 minus.n10 63.5369
R101 minus.n16 minus.n15 63.5369
R102 minus.n18 minus.n8 36.455
R103 minus.n6 minus.n5 9.49444
R104 minus.n4 minus.n1 9.49444
R105 minus.n13 minus.n10 9.49444
R106 minus.n15 minus.n14 9.49444
R107 minus.n18 minus.n17 6.46262
R108 minus.n8 minus.n0 0.189894
R109 minus.n3 minus.n0 0.189894
R110 minus.n12 minus.n9 0.189894
R111 minus.n17 minus.n9 0.189894
R112 minus minus.n18 0.188
R113 drain_right.n5 drain_right.n3 61.4227
R114 drain_right.n2 drain_right.n1 61.0958
R115 drain_right.n2 drain_right.n0 61.0958
R116 drain_right.n5 drain_right.n4 60.8798
R117 drain_right drain_right.n2 30.9874
R118 drain_right drain_right.n5 6.19632
R119 drain_right.n1 drain_right.t6 1.3205
R120 drain_right.n1 drain_right.t2 1.3205
R121 drain_right.n0 drain_right.t5 1.3205
R122 drain_right.n0 drain_right.t1 1.3205
R123 drain_right.n3 drain_right.t0 1.3205
R124 drain_right.n3 drain_right.t3 1.3205
R125 drain_right.n4 drain_right.t4 1.3205
R126 drain_right.n4 drain_right.t7 1.3205
C0 plus source 3.56353f
C1 plus drain_left 4.24035f
C2 drain_left source 20.249802f
C3 plus drain_right 0.280736f
C4 drain_right source 20.249f
C5 drain_right drain_left 0.630082f
C6 plus minus 5.387721f
C7 source minus 3.54949f
C8 drain_left minus 0.170671f
C9 drain_right minus 4.11315f
C10 drain_right a_n1346_n3888# 6.408319f
C11 drain_left a_n1346_n3888# 6.60581f
C12 source a_n1346_n3888# 10.173094f
C13 minus a_n1346_n3888# 5.388625f
C14 plus a_n1346_n3888# 7.60897f
C15 drain_right.t5 a_n1346_n3888# 0.39458f
C16 drain_right.t1 a_n1346_n3888# 0.39458f
C17 drain_right.n0 a_n1346_n3888# 3.56785f
C18 drain_right.t6 a_n1346_n3888# 0.39458f
C19 drain_right.t2 a_n1346_n3888# 0.39458f
C20 drain_right.n1 a_n1346_n3888# 3.56785f
C21 drain_right.n2 a_n1346_n3888# 2.36389f
C22 drain_right.t0 a_n1346_n3888# 0.39458f
C23 drain_right.t3 a_n1346_n3888# 0.39458f
C24 drain_right.n3 a_n1346_n3888# 3.57009f
C25 drain_right.t4 a_n1346_n3888# 0.39458f
C26 drain_right.t7 a_n1346_n3888# 0.39458f
C27 drain_right.n4 a_n1346_n3888# 3.56654f
C28 drain_right.n5 a_n1346_n3888# 1.06525f
C29 minus.n0 a_n1346_n3888# 0.055056f
C30 minus.t3 a_n1346_n3888# 0.704661f
C31 minus.t0 a_n1346_n3888# 0.698949f
C32 minus.t7 a_n1346_n3888# 0.698949f
C33 minus.n1 a_n1346_n3888# 0.26847f
C34 minus.t4 a_n1346_n3888# 0.704661f
C35 minus.n2 a_n1346_n3888# 0.285338f
C36 minus.n3 a_n1346_n3888# 0.11649f
C37 minus.n4 a_n1346_n3888# 0.02047f
C38 minus.n5 a_n1346_n3888# 0.02047f
C39 minus.n6 a_n1346_n3888# 0.26847f
C40 minus.n7 a_n1346_n3888# 0.285266f
C41 minus.n8 a_n1346_n3888# 1.96614f
C42 minus.n9 a_n1346_n3888# 0.055056f
C43 minus.t1 a_n1346_n3888# 0.698949f
C44 minus.t6 a_n1346_n3888# 0.698949f
C45 minus.n10 a_n1346_n3888# 0.26847f
C46 minus.t2 a_n1346_n3888# 0.704661f
C47 minus.n11 a_n1346_n3888# 0.285338f
C48 minus.n12 a_n1346_n3888# 0.11649f
C49 minus.n13 a_n1346_n3888# 0.02047f
C50 minus.n14 a_n1346_n3888# 0.02047f
C51 minus.n15 a_n1346_n3888# 0.26847f
C52 minus.t5 a_n1346_n3888# 0.704661f
C53 minus.n16 a_n1346_n3888# 0.285266f
C54 minus.n17 a_n1346_n3888# 0.355087f
C55 minus.n18 a_n1346_n3888# 2.38811f
C56 drain_left.t1 a_n1346_n3888# 0.394092f
C57 drain_left.t6 a_n1346_n3888# 0.394092f
C58 drain_left.n0 a_n1346_n3888# 3.56344f
C59 drain_left.t3 a_n1346_n3888# 0.394092f
C60 drain_left.t7 a_n1346_n3888# 0.394092f
C61 drain_left.n1 a_n1346_n3888# 3.56344f
C62 drain_left.n2 a_n1346_n3888# 2.43078f
C63 drain_left.t5 a_n1346_n3888# 0.394092f
C64 drain_left.t4 a_n1346_n3888# 0.394092f
C65 drain_left.n3 a_n1346_n3888# 3.56569f
C66 drain_left.t2 a_n1346_n3888# 0.394092f
C67 drain_left.t0 a_n1346_n3888# 0.394092f
C68 drain_left.n4 a_n1346_n3888# 3.56212f
C69 drain_left.n5 a_n1346_n3888# 1.06393f
C70 source.t12 a_n1346_n3888# 3.14023f
C71 source.n0 a_n1346_n3888# 1.45449f
C72 source.t13 a_n1346_n3888# 0.280212f
C73 source.t14 a_n1346_n3888# 0.280212f
C74 source.n1 a_n1346_n3888# 2.46143f
C75 source.n2 a_n1346_n3888# 0.315593f
C76 source.t8 a_n1346_n3888# 3.14023f
C77 source.n3 a_n1346_n3888# 0.395422f
C78 source.t5 a_n1346_n3888# 3.14023f
C79 source.n4 a_n1346_n3888# 0.395422f
C80 source.t0 a_n1346_n3888# 0.280212f
C81 source.t4 a_n1346_n3888# 0.280212f
C82 source.n5 a_n1346_n3888# 2.46143f
C83 source.n6 a_n1346_n3888# 0.315593f
C84 source.t3 a_n1346_n3888# 3.14023f
C85 source.n7 a_n1346_n3888# 1.84752f
C86 source.t15 a_n1346_n3888# 3.14023f
C87 source.n8 a_n1346_n3888# 1.84752f
C88 source.t11 a_n1346_n3888# 0.280212f
C89 source.t10 a_n1346_n3888# 0.280212f
C90 source.n9 a_n1346_n3888# 2.46142f
C91 source.n10 a_n1346_n3888# 0.315596f
C92 source.t9 a_n1346_n3888# 3.14023f
C93 source.n11 a_n1346_n3888# 0.395426f
C94 source.t2 a_n1346_n3888# 3.14023f
C95 source.n12 a_n1346_n3888# 0.395426f
C96 source.t6 a_n1346_n3888# 0.280212f
C97 source.t7 a_n1346_n3888# 0.280212f
C98 source.n13 a_n1346_n3888# 2.46142f
C99 source.n14 a_n1346_n3888# 0.315596f
C100 source.t1 a_n1346_n3888# 3.14023f
C101 source.n15 a_n1346_n3888# 0.528872f
C102 source.n16 a_n1346_n3888# 1.7285f
C103 plus.n0 a_n1346_n3888# 0.056386f
C104 plus.t5 a_n1346_n3888# 0.715833f
C105 plus.t3 a_n1346_n3888# 0.715833f
C106 plus.n1 a_n1346_n3888# 0.274956f
C107 plus.t2 a_n1346_n3888# 0.721682f
C108 plus.n2 a_n1346_n3888# 0.292231f
C109 plus.n3 a_n1346_n3888# 0.119304f
C110 plus.n4 a_n1346_n3888# 0.020965f
C111 plus.n5 a_n1346_n3888# 0.020965f
C112 plus.n6 a_n1346_n3888# 0.274956f
C113 plus.t7 a_n1346_n3888# 0.721682f
C114 plus.n7 a_n1346_n3888# 0.292157f
C115 plus.n8 a_n1346_n3888# 0.707573f
C116 plus.n9 a_n1346_n3888# 0.056386f
C117 plus.t6 a_n1346_n3888# 0.721682f
C118 plus.t1 a_n1346_n3888# 0.715833f
C119 plus.t4 a_n1346_n3888# 0.715833f
C120 plus.n10 a_n1346_n3888# 0.274956f
C121 plus.t0 a_n1346_n3888# 0.721682f
C122 plus.n11 a_n1346_n3888# 0.292231f
C123 plus.n12 a_n1346_n3888# 0.119304f
C124 plus.n13 a_n1346_n3888# 0.020965f
C125 plus.n14 a_n1346_n3888# 0.020965f
C126 plus.n15 a_n1346_n3888# 0.274956f
C127 plus.n16 a_n1346_n3888# 0.292157f
C128 plus.n17 a_n1346_n3888# 1.64741f
.ends

