* NGSPICE file created from diffpair549.ext - technology: sky130A

.subckt diffpair549 minus drain_right drain_left source plus
X0 a_n3394_n3888# a_n3394_n3888# a_n3394_n3888# a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.7
X1 source.t36 plus.t0 drain_left.t13 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X2 drain_left.t17 plus.t1 source.t35 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X3 source.t34 plus.t2 drain_left.t16 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X4 source.t40 minus.t0 drain_right.t23 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X5 drain_left.t23 plus.t3 source.t33 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X6 source.t32 plus.t4 drain_left.t22 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X7 source.t31 plus.t5 drain_left.t19 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X8 source.t9 minus.t1 drain_right.t22 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X9 drain_right.t21 minus.t2 source.t37 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X10 drain_left.t18 plus.t6 source.t30 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X11 source.t29 plus.t7 drain_left.t1 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X12 source.t28 plus.t8 drain_left.t0 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X13 drain_right.t20 minus.t3 source.t39 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X14 source.t8 minus.t4 drain_right.t19 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X15 source.t43 minus.t5 drain_right.t18 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X16 drain_right.t17 minus.t6 source.t1 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X17 source.t27 plus.t9 drain_left.t15 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X18 drain_left.t14 plus.t10 source.t26 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X19 drain_right.t16 minus.t7 source.t7 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X20 source.t38 minus.t8 drain_right.t15 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X21 drain_right.t14 minus.t9 source.t41 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X22 drain_right.t13 minus.t10 source.t0 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X23 drain_right.t12 minus.t11 source.t45 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X24 drain_right.t11 minus.t12 source.t5 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X25 drain_left.t5 plus.t11 source.t25 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X26 drain_right.t10 minus.t13 source.t11 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X27 a_n3394_n3888# a_n3394_n3888# a_n3394_n3888# a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.7
X28 drain_left.t4 plus.t12 source.t24 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X29 source.t23 plus.t13 drain_left.t8 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X30 drain_left.t7 plus.t14 source.t22 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X31 drain_right.t9 minus.t14 source.t4 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X32 a_n3394_n3888# a_n3394_n3888# a_n3394_n3888# a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.7
X33 source.t21 plus.t15 drain_left.t10 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X34 drain_left.t9 plus.t16 source.t20 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X35 drain_left.t3 plus.t17 source.t19 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X36 source.t47 minus.t15 drain_right.t8 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X37 source.t2 minus.t16 drain_right.t7 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X38 drain_right.t6 minus.t17 source.t46 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X39 source.t44 minus.t18 drain_right.t5 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X40 drain_left.t2 plus.t18 source.t18 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X41 source.t17 plus.t19 drain_left.t12 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X42 drain_left.t11 plus.t20 source.t16 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X43 source.t3 minus.t19 drain_right.t4 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X44 drain_left.t21 plus.t21 source.t15 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X45 source.t14 plus.t22 drain_left.t20 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X46 source.t10 minus.t20 drain_right.t3 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X47 source.t42 minus.t21 drain_right.t2 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X48 a_n3394_n3888# a_n3394_n3888# a_n3394_n3888# a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.7
X49 source.t13 plus.t23 drain_left.t6 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X50 source.t12 minus.t22 drain_right.t1 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X51 drain_right.t0 minus.t23 source.t6 a_n3394_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
R0 plus.n11 plus.t8 598.907
R1 plus.n53 plus.t3 598.907
R2 plus.n40 plus.t1 572.548
R3 plus.n38 plus.t13 572.548
R4 plus.n2 plus.t6 572.548
R5 plus.n32 plus.t23 572.548
R6 plus.n4 plus.t11 572.548
R7 plus.n26 plus.t2 572.548
R8 plus.n6 plus.t14 572.548
R9 plus.n20 plus.t7 572.548
R10 plus.n8 plus.t12 572.548
R11 plus.n14 plus.t5 572.548
R12 plus.n10 plus.t17 572.548
R13 plus.n82 plus.t22 572.548
R14 plus.n80 plus.t20 572.548
R15 plus.n44 plus.t19 572.548
R16 plus.n74 plus.t18 572.548
R17 plus.n46 plus.t0 572.548
R18 plus.n68 plus.t10 572.548
R19 plus.n48 plus.t9 572.548
R20 plus.n62 plus.t16 572.548
R21 plus.n50 plus.t15 572.548
R22 plus.n56 plus.t21 572.548
R23 plus.n52 plus.t4 572.548
R24 plus.n13 plus.n12 161.3
R25 plus.n14 plus.n9 161.3
R26 plus.n16 plus.n15 161.3
R27 plus.n17 plus.n8 161.3
R28 plus.n19 plus.n18 161.3
R29 plus.n20 plus.n7 161.3
R30 plus.n22 plus.n21 161.3
R31 plus.n23 plus.n6 161.3
R32 plus.n25 plus.n24 161.3
R33 plus.n26 plus.n5 161.3
R34 plus.n28 plus.n27 161.3
R35 plus.n29 plus.n4 161.3
R36 plus.n31 plus.n30 161.3
R37 plus.n32 plus.n3 161.3
R38 plus.n34 plus.n33 161.3
R39 plus.n35 plus.n2 161.3
R40 plus.n37 plus.n36 161.3
R41 plus.n38 plus.n1 161.3
R42 plus.n39 plus.n0 161.3
R43 plus.n41 plus.n40 161.3
R44 plus.n55 plus.n54 161.3
R45 plus.n56 plus.n51 161.3
R46 plus.n58 plus.n57 161.3
R47 plus.n59 plus.n50 161.3
R48 plus.n61 plus.n60 161.3
R49 plus.n62 plus.n49 161.3
R50 plus.n64 plus.n63 161.3
R51 plus.n65 plus.n48 161.3
R52 plus.n67 plus.n66 161.3
R53 plus.n68 plus.n47 161.3
R54 plus.n70 plus.n69 161.3
R55 plus.n71 plus.n46 161.3
R56 plus.n73 plus.n72 161.3
R57 plus.n74 plus.n45 161.3
R58 plus.n76 plus.n75 161.3
R59 plus.n77 plus.n44 161.3
R60 plus.n79 plus.n78 161.3
R61 plus.n80 plus.n43 161.3
R62 plus.n81 plus.n42 161.3
R63 plus.n83 plus.n82 161.3
R64 plus.n40 plus.n39 46.0096
R65 plus.n82 plus.n81 46.0096
R66 plus.n12 plus.n11 45.0871
R67 plus.n54 plus.n53 45.0871
R68 plus.n38 plus.n37 41.6278
R69 plus.n13 plus.n10 41.6278
R70 plus.n80 plus.n79 41.6278
R71 plus.n55 plus.n52 41.6278
R72 plus.n33 plus.n2 37.246
R73 plus.n15 plus.n14 37.246
R74 plus.n75 plus.n44 37.246
R75 plus.n57 plus.n56 37.246
R76 plus plus.n83 37.1733
R77 plus.n32 plus.n31 32.8641
R78 plus.n19 plus.n8 32.8641
R79 plus.n74 plus.n73 32.8641
R80 plus.n61 plus.n50 32.8641
R81 plus.n27 plus.n4 28.4823
R82 plus.n21 plus.n20 28.4823
R83 plus.n69 plus.n46 28.4823
R84 plus.n63 plus.n62 28.4823
R85 plus.n25 plus.n6 24.1005
R86 plus.n26 plus.n25 24.1005
R87 plus.n68 plus.n67 24.1005
R88 plus.n67 plus.n48 24.1005
R89 plus.n27 plus.n26 19.7187
R90 plus.n21 plus.n6 19.7187
R91 plus.n69 plus.n68 19.7187
R92 plus.n63 plus.n48 19.7187
R93 plus.n31 plus.n4 15.3369
R94 plus.n20 plus.n19 15.3369
R95 plus.n73 plus.n46 15.3369
R96 plus.n62 plus.n61 15.3369
R97 plus.n11 plus.n10 14.1472
R98 plus.n53 plus.n52 14.1472
R99 plus plus.n41 13.4588
R100 plus.n33 plus.n32 10.955
R101 plus.n15 plus.n8 10.955
R102 plus.n75 plus.n74 10.955
R103 plus.n57 plus.n50 10.955
R104 plus.n37 plus.n2 6.57323
R105 plus.n14 plus.n13 6.57323
R106 plus.n79 plus.n44 6.57323
R107 plus.n56 plus.n55 6.57323
R108 plus.n39 plus.n38 2.19141
R109 plus.n81 plus.n80 2.19141
R110 plus.n12 plus.n9 0.189894
R111 plus.n16 plus.n9 0.189894
R112 plus.n17 plus.n16 0.189894
R113 plus.n18 plus.n17 0.189894
R114 plus.n18 plus.n7 0.189894
R115 plus.n22 plus.n7 0.189894
R116 plus.n23 plus.n22 0.189894
R117 plus.n24 plus.n23 0.189894
R118 plus.n24 plus.n5 0.189894
R119 plus.n28 plus.n5 0.189894
R120 plus.n29 plus.n28 0.189894
R121 plus.n30 plus.n29 0.189894
R122 plus.n30 plus.n3 0.189894
R123 plus.n34 plus.n3 0.189894
R124 plus.n35 plus.n34 0.189894
R125 plus.n36 plus.n35 0.189894
R126 plus.n36 plus.n1 0.189894
R127 plus.n1 plus.n0 0.189894
R128 plus.n41 plus.n0 0.189894
R129 plus.n83 plus.n42 0.189894
R130 plus.n43 plus.n42 0.189894
R131 plus.n78 plus.n43 0.189894
R132 plus.n78 plus.n77 0.189894
R133 plus.n77 plus.n76 0.189894
R134 plus.n76 plus.n45 0.189894
R135 plus.n72 plus.n45 0.189894
R136 plus.n72 plus.n71 0.189894
R137 plus.n71 plus.n70 0.189894
R138 plus.n70 plus.n47 0.189894
R139 plus.n66 plus.n47 0.189894
R140 plus.n66 plus.n65 0.189894
R141 plus.n65 plus.n64 0.189894
R142 plus.n64 plus.n49 0.189894
R143 plus.n60 plus.n49 0.189894
R144 plus.n60 plus.n59 0.189894
R145 plus.n59 plus.n58 0.189894
R146 plus.n58 plus.n51 0.189894
R147 plus.n54 plus.n51 0.189894
R148 drain_left.n13 drain_left.n11 61.7677
R149 drain_left.n7 drain_left.n5 61.7675
R150 drain_left.n2 drain_left.n0 61.7675
R151 drain_left.n19 drain_left.n18 60.8798
R152 drain_left.n17 drain_left.n16 60.8798
R153 drain_left.n15 drain_left.n14 60.8798
R154 drain_left.n13 drain_left.n12 60.8798
R155 drain_left.n21 drain_left.n20 60.8796
R156 drain_left.n7 drain_left.n6 60.8796
R157 drain_left.n9 drain_left.n8 60.8796
R158 drain_left.n4 drain_left.n3 60.8796
R159 drain_left.n2 drain_left.n1 60.8796
R160 drain_left drain_left.n10 38.0751
R161 drain_left drain_left.n21 6.54115
R162 drain_left.n5 drain_left.t22 1.3205
R163 drain_left.n5 drain_left.t23 1.3205
R164 drain_left.n6 drain_left.t10 1.3205
R165 drain_left.n6 drain_left.t21 1.3205
R166 drain_left.n8 drain_left.t15 1.3205
R167 drain_left.n8 drain_left.t9 1.3205
R168 drain_left.n3 drain_left.t13 1.3205
R169 drain_left.n3 drain_left.t14 1.3205
R170 drain_left.n1 drain_left.t12 1.3205
R171 drain_left.n1 drain_left.t2 1.3205
R172 drain_left.n0 drain_left.t20 1.3205
R173 drain_left.n0 drain_left.t11 1.3205
R174 drain_left.n20 drain_left.t8 1.3205
R175 drain_left.n20 drain_left.t17 1.3205
R176 drain_left.n18 drain_left.t6 1.3205
R177 drain_left.n18 drain_left.t18 1.3205
R178 drain_left.n16 drain_left.t16 1.3205
R179 drain_left.n16 drain_left.t5 1.3205
R180 drain_left.n14 drain_left.t1 1.3205
R181 drain_left.n14 drain_left.t7 1.3205
R182 drain_left.n12 drain_left.t19 1.3205
R183 drain_left.n12 drain_left.t4 1.3205
R184 drain_left.n11 drain_left.t0 1.3205
R185 drain_left.n11 drain_left.t3 1.3205
R186 drain_left.n9 drain_left.n7 0.888431
R187 drain_left.n4 drain_left.n2 0.888431
R188 drain_left.n15 drain_left.n13 0.888431
R189 drain_left.n17 drain_left.n15 0.888431
R190 drain_left.n19 drain_left.n17 0.888431
R191 drain_left.n21 drain_left.n19 0.888431
R192 drain_left.n10 drain_left.n9 0.389119
R193 drain_left.n10 drain_left.n4 0.389119
R194 source.n11 source.t28 45.521
R195 source.n12 source.t4 45.521
R196 source.n23 source.t47 45.521
R197 source.n47 source.t1 45.5208
R198 source.n36 source.t38 45.5208
R199 source.n35 source.t33 45.5208
R200 source.n24 source.t14 45.5208
R201 source.n0 source.t35 45.5208
R202 source.n2 source.n1 44.201
R203 source.n4 source.n3 44.201
R204 source.n6 source.n5 44.201
R205 source.n8 source.n7 44.201
R206 source.n10 source.n9 44.201
R207 source.n14 source.n13 44.201
R208 source.n16 source.n15 44.201
R209 source.n18 source.n17 44.201
R210 source.n20 source.n19 44.201
R211 source.n22 source.n21 44.201
R212 source.n46 source.n45 44.2008
R213 source.n44 source.n43 44.2008
R214 source.n42 source.n41 44.2008
R215 source.n40 source.n39 44.2008
R216 source.n38 source.n37 44.2008
R217 source.n34 source.n33 44.2008
R218 source.n32 source.n31 44.2008
R219 source.n30 source.n29 44.2008
R220 source.n28 source.n27 44.2008
R221 source.n26 source.n25 44.2008
R222 source.n24 source.n23 24.4484
R223 source.n48 source.n0 18.7415
R224 source.n48 source.n47 5.7074
R225 source.n45 source.t5 1.3205
R226 source.n45 source.t8 1.3205
R227 source.n43 source.t46 1.3205
R228 source.n43 source.t44 1.3205
R229 source.n41 source.t6 1.3205
R230 source.n41 source.t12 1.3205
R231 source.n39 source.t37 1.3205
R232 source.n39 source.t43 1.3205
R233 source.n37 source.t41 1.3205
R234 source.n37 source.t40 1.3205
R235 source.n33 source.t15 1.3205
R236 source.n33 source.t32 1.3205
R237 source.n31 source.t20 1.3205
R238 source.n31 source.t21 1.3205
R239 source.n29 source.t26 1.3205
R240 source.n29 source.t27 1.3205
R241 source.n27 source.t18 1.3205
R242 source.n27 source.t36 1.3205
R243 source.n25 source.t16 1.3205
R244 source.n25 source.t17 1.3205
R245 source.n1 source.t30 1.3205
R246 source.n1 source.t23 1.3205
R247 source.n3 source.t25 1.3205
R248 source.n3 source.t13 1.3205
R249 source.n5 source.t22 1.3205
R250 source.n5 source.t34 1.3205
R251 source.n7 source.t24 1.3205
R252 source.n7 source.t29 1.3205
R253 source.n9 source.t19 1.3205
R254 source.n9 source.t31 1.3205
R255 source.n13 source.t11 1.3205
R256 source.n13 source.t9 1.3205
R257 source.n15 source.t45 1.3205
R258 source.n15 source.t10 1.3205
R259 source.n17 source.t0 1.3205
R260 source.n17 source.t42 1.3205
R261 source.n19 source.t7 1.3205
R262 source.n19 source.t3 1.3205
R263 source.n21 source.t39 1.3205
R264 source.n21 source.t2 1.3205
R265 source.n23 source.n22 0.888431
R266 source.n22 source.n20 0.888431
R267 source.n20 source.n18 0.888431
R268 source.n18 source.n16 0.888431
R269 source.n16 source.n14 0.888431
R270 source.n14 source.n12 0.888431
R271 source.n11 source.n10 0.888431
R272 source.n10 source.n8 0.888431
R273 source.n8 source.n6 0.888431
R274 source.n6 source.n4 0.888431
R275 source.n4 source.n2 0.888431
R276 source.n2 source.n0 0.888431
R277 source.n26 source.n24 0.888431
R278 source.n28 source.n26 0.888431
R279 source.n30 source.n28 0.888431
R280 source.n32 source.n30 0.888431
R281 source.n34 source.n32 0.888431
R282 source.n35 source.n34 0.888431
R283 source.n38 source.n36 0.888431
R284 source.n40 source.n38 0.888431
R285 source.n42 source.n40 0.888431
R286 source.n44 source.n42 0.888431
R287 source.n46 source.n44 0.888431
R288 source.n47 source.n46 0.888431
R289 source.n12 source.n11 0.470328
R290 source.n36 source.n35 0.470328
R291 source source.n48 0.188
R292 minus.n11 minus.t14 598.907
R293 minus.n53 minus.t8 598.907
R294 minus.n10 minus.t1 572.548
R295 minus.n14 minus.t13 572.548
R296 minus.n16 minus.t20 572.548
R297 minus.n20 minus.t11 572.548
R298 minus.n22 minus.t21 572.548
R299 minus.n26 minus.t10 572.548
R300 minus.n28 minus.t19 572.548
R301 minus.n32 minus.t7 572.548
R302 minus.n34 minus.t16 572.548
R303 minus.n38 minus.t3 572.548
R304 minus.n40 minus.t15 572.548
R305 minus.n52 minus.t9 572.548
R306 minus.n56 minus.t0 572.548
R307 minus.n58 minus.t2 572.548
R308 minus.n62 minus.t5 572.548
R309 minus.n64 minus.t23 572.548
R310 minus.n68 minus.t22 572.548
R311 minus.n70 minus.t17 572.548
R312 minus.n74 minus.t18 572.548
R313 minus.n76 minus.t12 572.548
R314 minus.n80 minus.t4 572.548
R315 minus.n82 minus.t6 572.548
R316 minus.n41 minus.n40 161.3
R317 minus.n39 minus.n0 161.3
R318 minus.n38 minus.n37 161.3
R319 minus.n36 minus.n1 161.3
R320 minus.n35 minus.n34 161.3
R321 minus.n33 minus.n2 161.3
R322 minus.n32 minus.n31 161.3
R323 minus.n30 minus.n3 161.3
R324 minus.n29 minus.n28 161.3
R325 minus.n27 minus.n4 161.3
R326 minus.n26 minus.n25 161.3
R327 minus.n24 minus.n5 161.3
R328 minus.n23 minus.n22 161.3
R329 minus.n21 minus.n6 161.3
R330 minus.n20 minus.n19 161.3
R331 minus.n18 minus.n7 161.3
R332 minus.n17 minus.n16 161.3
R333 minus.n15 minus.n8 161.3
R334 minus.n14 minus.n13 161.3
R335 minus.n12 minus.n9 161.3
R336 minus.n83 minus.n82 161.3
R337 minus.n81 minus.n42 161.3
R338 minus.n80 minus.n79 161.3
R339 minus.n78 minus.n43 161.3
R340 minus.n77 minus.n76 161.3
R341 minus.n75 minus.n44 161.3
R342 minus.n74 minus.n73 161.3
R343 minus.n72 minus.n45 161.3
R344 minus.n71 minus.n70 161.3
R345 minus.n69 minus.n46 161.3
R346 minus.n68 minus.n67 161.3
R347 minus.n66 minus.n47 161.3
R348 minus.n65 minus.n64 161.3
R349 minus.n63 minus.n48 161.3
R350 minus.n62 minus.n61 161.3
R351 minus.n60 minus.n49 161.3
R352 minus.n59 minus.n58 161.3
R353 minus.n57 minus.n50 161.3
R354 minus.n56 minus.n55 161.3
R355 minus.n54 minus.n51 161.3
R356 minus.n40 minus.n39 46.0096
R357 minus.n82 minus.n81 46.0096
R358 minus.n12 minus.n11 45.0871
R359 minus.n54 minus.n53 45.0871
R360 minus.n84 minus.n41 44.4285
R361 minus.n10 minus.n9 41.6278
R362 minus.n38 minus.n1 41.6278
R363 minus.n52 minus.n51 41.6278
R364 minus.n80 minus.n43 41.6278
R365 minus.n15 minus.n14 37.246
R366 minus.n34 minus.n33 37.246
R367 minus.n57 minus.n56 37.246
R368 minus.n76 minus.n75 37.246
R369 minus.n16 minus.n7 32.8641
R370 minus.n32 minus.n3 32.8641
R371 minus.n58 minus.n49 32.8641
R372 minus.n74 minus.n45 32.8641
R373 minus.n21 minus.n20 28.4823
R374 minus.n28 minus.n27 28.4823
R375 minus.n63 minus.n62 28.4823
R376 minus.n70 minus.n69 28.4823
R377 minus.n26 minus.n5 24.1005
R378 minus.n22 minus.n5 24.1005
R379 minus.n64 minus.n47 24.1005
R380 minus.n68 minus.n47 24.1005
R381 minus.n22 minus.n21 19.7187
R382 minus.n27 minus.n26 19.7187
R383 minus.n64 minus.n63 19.7187
R384 minus.n69 minus.n68 19.7187
R385 minus.n20 minus.n7 15.3369
R386 minus.n28 minus.n3 15.3369
R387 minus.n62 minus.n49 15.3369
R388 minus.n70 minus.n45 15.3369
R389 minus.n11 minus.n10 14.1472
R390 minus.n53 minus.n52 14.1472
R391 minus.n16 minus.n15 10.955
R392 minus.n33 minus.n32 10.955
R393 minus.n58 minus.n57 10.955
R394 minus.n75 minus.n74 10.955
R395 minus.n84 minus.n83 6.67853
R396 minus.n14 minus.n9 6.57323
R397 minus.n34 minus.n1 6.57323
R398 minus.n56 minus.n51 6.57323
R399 minus.n76 minus.n43 6.57323
R400 minus.n39 minus.n38 2.19141
R401 minus.n81 minus.n80 2.19141
R402 minus.n41 minus.n0 0.189894
R403 minus.n37 minus.n0 0.189894
R404 minus.n37 minus.n36 0.189894
R405 minus.n36 minus.n35 0.189894
R406 minus.n35 minus.n2 0.189894
R407 minus.n31 minus.n2 0.189894
R408 minus.n31 minus.n30 0.189894
R409 minus.n30 minus.n29 0.189894
R410 minus.n29 minus.n4 0.189894
R411 minus.n25 minus.n4 0.189894
R412 minus.n25 minus.n24 0.189894
R413 minus.n24 minus.n23 0.189894
R414 minus.n23 minus.n6 0.189894
R415 minus.n19 minus.n6 0.189894
R416 minus.n19 minus.n18 0.189894
R417 minus.n18 minus.n17 0.189894
R418 minus.n17 minus.n8 0.189894
R419 minus.n13 minus.n8 0.189894
R420 minus.n13 minus.n12 0.189894
R421 minus.n55 minus.n54 0.189894
R422 minus.n55 minus.n50 0.189894
R423 minus.n59 minus.n50 0.189894
R424 minus.n60 minus.n59 0.189894
R425 minus.n61 minus.n60 0.189894
R426 minus.n61 minus.n48 0.189894
R427 minus.n65 minus.n48 0.189894
R428 minus.n66 minus.n65 0.189894
R429 minus.n67 minus.n66 0.189894
R430 minus.n67 minus.n46 0.189894
R431 minus.n71 minus.n46 0.189894
R432 minus.n72 minus.n71 0.189894
R433 minus.n73 minus.n72 0.189894
R434 minus.n73 minus.n44 0.189894
R435 minus.n77 minus.n44 0.189894
R436 minus.n78 minus.n77 0.189894
R437 minus.n79 minus.n78 0.189894
R438 minus.n79 minus.n42 0.189894
R439 minus.n83 minus.n42 0.189894
R440 minus minus.n84 0.188
R441 drain_right.n13 drain_right.n11 61.7676
R442 drain_right.n7 drain_right.n5 61.7675
R443 drain_right.n2 drain_right.n0 61.7675
R444 drain_right.n13 drain_right.n12 60.8798
R445 drain_right.n15 drain_right.n14 60.8798
R446 drain_right.n17 drain_right.n16 60.8798
R447 drain_right.n19 drain_right.n18 60.8798
R448 drain_right.n21 drain_right.n20 60.8798
R449 drain_right.n7 drain_right.n6 60.8796
R450 drain_right.n9 drain_right.n8 60.8796
R451 drain_right.n4 drain_right.n3 60.8796
R452 drain_right.n2 drain_right.n1 60.8796
R453 drain_right drain_right.n10 37.5219
R454 drain_right drain_right.n21 6.54115
R455 drain_right.n5 drain_right.t19 1.3205
R456 drain_right.n5 drain_right.t17 1.3205
R457 drain_right.n6 drain_right.t5 1.3205
R458 drain_right.n6 drain_right.t11 1.3205
R459 drain_right.n8 drain_right.t1 1.3205
R460 drain_right.n8 drain_right.t6 1.3205
R461 drain_right.n3 drain_right.t18 1.3205
R462 drain_right.n3 drain_right.t0 1.3205
R463 drain_right.n1 drain_right.t23 1.3205
R464 drain_right.n1 drain_right.t21 1.3205
R465 drain_right.n0 drain_right.t15 1.3205
R466 drain_right.n0 drain_right.t14 1.3205
R467 drain_right.n11 drain_right.t22 1.3205
R468 drain_right.n11 drain_right.t9 1.3205
R469 drain_right.n12 drain_right.t3 1.3205
R470 drain_right.n12 drain_right.t10 1.3205
R471 drain_right.n14 drain_right.t2 1.3205
R472 drain_right.n14 drain_right.t12 1.3205
R473 drain_right.n16 drain_right.t4 1.3205
R474 drain_right.n16 drain_right.t13 1.3205
R475 drain_right.n18 drain_right.t7 1.3205
R476 drain_right.n18 drain_right.t16 1.3205
R477 drain_right.n20 drain_right.t8 1.3205
R478 drain_right.n20 drain_right.t20 1.3205
R479 drain_right.n9 drain_right.n7 0.888431
R480 drain_right.n4 drain_right.n2 0.888431
R481 drain_right.n21 drain_right.n19 0.888431
R482 drain_right.n19 drain_right.n17 0.888431
R483 drain_right.n17 drain_right.n15 0.888431
R484 drain_right.n15 drain_right.n13 0.888431
R485 drain_right.n10 drain_right.n9 0.389119
R486 drain_right.n10 drain_right.n4 0.389119
C0 drain_left minus 0.174517f
C1 drain_right plus 0.498726f
C2 drain_left source 34.254803f
C3 drain_right minus 18.478699f
C4 drain_right source 34.2573f
C5 minus plus 7.93645f
C6 drain_right drain_left 1.87044f
C7 source plus 18.6661f
C8 drain_left plus 18.819199f
C9 source minus 18.6521f
C10 drain_right a_n3394_n3888# 8.4403f
C11 drain_left a_n3394_n3888# 8.906859f
C12 source a_n3394_n3888# 11.256248f
C13 minus a_n3394_n3888# 13.948141f
C14 plus a_n3394_n3888# 15.979861f
C15 drain_right.t15 a_n3394_n3888# 0.322578f
C16 drain_right.t14 a_n3394_n3888# 0.322578f
C17 drain_right.n0 a_n3394_n3888# 2.92133f
C18 drain_right.t23 a_n3394_n3888# 0.322578f
C19 drain_right.t21 a_n3394_n3888# 0.322578f
C20 drain_right.n1 a_n3394_n3888# 2.91573f
C21 drain_right.n2 a_n3394_n3888# 0.762604f
C22 drain_right.t18 a_n3394_n3888# 0.322578f
C23 drain_right.t0 a_n3394_n3888# 0.322578f
C24 drain_right.n3 a_n3394_n3888# 2.91573f
C25 drain_right.n4 a_n3394_n3888# 0.336461f
C26 drain_right.t19 a_n3394_n3888# 0.322578f
C27 drain_right.t17 a_n3394_n3888# 0.322578f
C28 drain_right.n5 a_n3394_n3888# 2.92133f
C29 drain_right.t5 a_n3394_n3888# 0.322578f
C30 drain_right.t11 a_n3394_n3888# 0.322578f
C31 drain_right.n6 a_n3394_n3888# 2.91573f
C32 drain_right.n7 a_n3394_n3888# 0.762604f
C33 drain_right.t1 a_n3394_n3888# 0.322578f
C34 drain_right.t6 a_n3394_n3888# 0.322578f
C35 drain_right.n8 a_n3394_n3888# 2.91573f
C36 drain_right.n9 a_n3394_n3888# 0.336461f
C37 drain_right.n10 a_n3394_n3888# 1.93527f
C38 drain_right.t22 a_n3394_n3888# 0.322578f
C39 drain_right.t9 a_n3394_n3888# 0.322578f
C40 drain_right.n11 a_n3394_n3888# 2.92132f
C41 drain_right.t3 a_n3394_n3888# 0.322578f
C42 drain_right.t10 a_n3394_n3888# 0.322578f
C43 drain_right.n12 a_n3394_n3888# 2.91573f
C44 drain_right.n13 a_n3394_n3888# 0.762609f
C45 drain_right.t2 a_n3394_n3888# 0.322578f
C46 drain_right.t12 a_n3394_n3888# 0.322578f
C47 drain_right.n14 a_n3394_n3888# 2.91573f
C48 drain_right.n15 a_n3394_n3888# 0.378619f
C49 drain_right.t4 a_n3394_n3888# 0.322578f
C50 drain_right.t13 a_n3394_n3888# 0.322578f
C51 drain_right.n16 a_n3394_n3888# 2.91573f
C52 drain_right.n17 a_n3394_n3888# 0.378619f
C53 drain_right.t7 a_n3394_n3888# 0.322578f
C54 drain_right.t16 a_n3394_n3888# 0.322578f
C55 drain_right.n18 a_n3394_n3888# 2.91573f
C56 drain_right.n19 a_n3394_n3888# 0.378619f
C57 drain_right.t8 a_n3394_n3888# 0.322578f
C58 drain_right.t20 a_n3394_n3888# 0.322578f
C59 drain_right.n20 a_n3394_n3888# 2.91573f
C60 drain_right.n21 a_n3394_n3888# 0.619327f
C61 minus.n0 a_n3394_n3888# 0.039048f
C62 minus.n1 a_n3394_n3888# 0.008861f
C63 minus.t3 a_n3394_n3888# 1.1651f
C64 minus.n2 a_n3394_n3888# 0.039048f
C65 minus.n3 a_n3394_n3888# 0.008861f
C66 minus.t7 a_n3394_n3888# 1.1651f
C67 minus.n4 a_n3394_n3888# 0.039048f
C68 minus.n5 a_n3394_n3888# 0.008861f
C69 minus.t10 a_n3394_n3888# 1.1651f
C70 minus.n6 a_n3394_n3888# 0.039048f
C71 minus.n7 a_n3394_n3888# 0.008861f
C72 minus.t11 a_n3394_n3888# 1.1651f
C73 minus.n8 a_n3394_n3888# 0.039048f
C74 minus.n9 a_n3394_n3888# 0.008861f
C75 minus.t13 a_n3394_n3888# 1.1651f
C76 minus.t14 a_n3394_n3888# 1.18492f
C77 minus.t1 a_n3394_n3888# 1.1651f
C78 minus.n10 a_n3394_n3888# 0.457608f
C79 minus.n11 a_n3394_n3888# 0.431878f
C80 minus.n12 a_n3394_n3888# 0.168103f
C81 minus.n13 a_n3394_n3888# 0.039048f
C82 minus.n14 a_n3394_n3888# 0.449617f
C83 minus.n15 a_n3394_n3888# 0.008861f
C84 minus.t20 a_n3394_n3888# 1.1651f
C85 minus.n16 a_n3394_n3888# 0.449617f
C86 minus.n17 a_n3394_n3888# 0.039048f
C87 minus.n18 a_n3394_n3888# 0.039048f
C88 minus.n19 a_n3394_n3888# 0.039048f
C89 minus.n20 a_n3394_n3888# 0.449617f
C90 minus.n21 a_n3394_n3888# 0.008861f
C91 minus.t21 a_n3394_n3888# 1.1651f
C92 minus.n22 a_n3394_n3888# 0.449617f
C93 minus.n23 a_n3394_n3888# 0.039048f
C94 minus.n24 a_n3394_n3888# 0.039048f
C95 minus.n25 a_n3394_n3888# 0.039048f
C96 minus.n26 a_n3394_n3888# 0.449617f
C97 minus.n27 a_n3394_n3888# 0.008861f
C98 minus.t19 a_n3394_n3888# 1.1651f
C99 minus.n28 a_n3394_n3888# 0.449617f
C100 minus.n29 a_n3394_n3888# 0.039048f
C101 minus.n30 a_n3394_n3888# 0.039048f
C102 minus.n31 a_n3394_n3888# 0.039048f
C103 minus.n32 a_n3394_n3888# 0.449617f
C104 minus.n33 a_n3394_n3888# 0.008861f
C105 minus.t16 a_n3394_n3888# 1.1651f
C106 minus.n34 a_n3394_n3888# 0.449617f
C107 minus.n35 a_n3394_n3888# 0.039048f
C108 minus.n36 a_n3394_n3888# 0.039048f
C109 minus.n37 a_n3394_n3888# 0.039048f
C110 minus.n38 a_n3394_n3888# 0.449617f
C111 minus.n39 a_n3394_n3888# 0.008861f
C112 minus.t15 a_n3394_n3888# 1.1651f
C113 minus.n40 a_n3394_n3888# 0.449978f
C114 minus.n41 a_n3394_n3888# 1.8813f
C115 minus.n42 a_n3394_n3888# 0.039048f
C116 minus.n43 a_n3394_n3888# 0.008861f
C117 minus.n44 a_n3394_n3888# 0.039048f
C118 minus.n45 a_n3394_n3888# 0.008861f
C119 minus.n46 a_n3394_n3888# 0.039048f
C120 minus.n47 a_n3394_n3888# 0.008861f
C121 minus.n48 a_n3394_n3888# 0.039048f
C122 minus.n49 a_n3394_n3888# 0.008861f
C123 minus.n50 a_n3394_n3888# 0.039048f
C124 minus.n51 a_n3394_n3888# 0.008861f
C125 minus.t8 a_n3394_n3888# 1.18492f
C126 minus.t9 a_n3394_n3888# 1.1651f
C127 minus.n52 a_n3394_n3888# 0.457608f
C128 minus.n53 a_n3394_n3888# 0.431878f
C129 minus.n54 a_n3394_n3888# 0.168103f
C130 minus.n55 a_n3394_n3888# 0.039048f
C131 minus.t0 a_n3394_n3888# 1.1651f
C132 minus.n56 a_n3394_n3888# 0.449617f
C133 minus.n57 a_n3394_n3888# 0.008861f
C134 minus.t2 a_n3394_n3888# 1.1651f
C135 minus.n58 a_n3394_n3888# 0.449617f
C136 minus.n59 a_n3394_n3888# 0.039048f
C137 minus.n60 a_n3394_n3888# 0.039048f
C138 minus.n61 a_n3394_n3888# 0.039048f
C139 minus.t5 a_n3394_n3888# 1.1651f
C140 minus.n62 a_n3394_n3888# 0.449617f
C141 minus.n63 a_n3394_n3888# 0.008861f
C142 minus.t23 a_n3394_n3888# 1.1651f
C143 minus.n64 a_n3394_n3888# 0.449617f
C144 minus.n65 a_n3394_n3888# 0.039048f
C145 minus.n66 a_n3394_n3888# 0.039048f
C146 minus.n67 a_n3394_n3888# 0.039048f
C147 minus.t22 a_n3394_n3888# 1.1651f
C148 minus.n68 a_n3394_n3888# 0.449617f
C149 minus.n69 a_n3394_n3888# 0.008861f
C150 minus.t17 a_n3394_n3888# 1.1651f
C151 minus.n70 a_n3394_n3888# 0.449617f
C152 minus.n71 a_n3394_n3888# 0.039048f
C153 minus.n72 a_n3394_n3888# 0.039048f
C154 minus.n73 a_n3394_n3888# 0.039048f
C155 minus.t18 a_n3394_n3888# 1.1651f
C156 minus.n74 a_n3394_n3888# 0.449617f
C157 minus.n75 a_n3394_n3888# 0.008861f
C158 minus.t12 a_n3394_n3888# 1.1651f
C159 minus.n76 a_n3394_n3888# 0.449617f
C160 minus.n77 a_n3394_n3888# 0.039048f
C161 minus.n78 a_n3394_n3888# 0.039048f
C162 minus.n79 a_n3394_n3888# 0.039048f
C163 minus.t4 a_n3394_n3888# 1.1651f
C164 minus.n80 a_n3394_n3888# 0.449617f
C165 minus.n81 a_n3394_n3888# 0.008861f
C166 minus.t6 a_n3394_n3888# 1.1651f
C167 minus.n82 a_n3394_n3888# 0.449978f
C168 minus.n83 a_n3394_n3888# 0.271573f
C169 minus.n84 a_n3394_n3888# 2.22815f
C170 source.t35 a_n3394_n3888# 3.25492f
C171 source.n0 a_n3394_n3888# 1.5515f
C172 source.t30 a_n3394_n3888# 0.290446f
C173 source.t23 a_n3394_n3888# 0.290446f
C174 source.n1 a_n3394_n3888# 2.55133f
C175 source.n2 a_n3394_n3888# 0.381571f
C176 source.t25 a_n3394_n3888# 0.290446f
C177 source.t13 a_n3394_n3888# 0.290446f
C178 source.n3 a_n3394_n3888# 2.55133f
C179 source.n4 a_n3394_n3888# 0.381571f
C180 source.t22 a_n3394_n3888# 0.290446f
C181 source.t34 a_n3394_n3888# 0.290446f
C182 source.n5 a_n3394_n3888# 2.55133f
C183 source.n6 a_n3394_n3888# 0.381571f
C184 source.t24 a_n3394_n3888# 0.290446f
C185 source.t29 a_n3394_n3888# 0.290446f
C186 source.n7 a_n3394_n3888# 2.55133f
C187 source.n8 a_n3394_n3888# 0.381571f
C188 source.t19 a_n3394_n3888# 0.290446f
C189 source.t31 a_n3394_n3888# 0.290446f
C190 source.n9 a_n3394_n3888# 2.55133f
C191 source.n10 a_n3394_n3888# 0.381571f
C192 source.t28 a_n3394_n3888# 3.25492f
C193 source.n11 a_n3394_n3888# 0.43709f
C194 source.t4 a_n3394_n3888# 3.25492f
C195 source.n12 a_n3394_n3888# 0.43709f
C196 source.t11 a_n3394_n3888# 0.290446f
C197 source.t9 a_n3394_n3888# 0.290446f
C198 source.n13 a_n3394_n3888# 2.55133f
C199 source.n14 a_n3394_n3888# 0.381571f
C200 source.t45 a_n3394_n3888# 0.290446f
C201 source.t10 a_n3394_n3888# 0.290446f
C202 source.n15 a_n3394_n3888# 2.55133f
C203 source.n16 a_n3394_n3888# 0.381571f
C204 source.t0 a_n3394_n3888# 0.290446f
C205 source.t42 a_n3394_n3888# 0.290446f
C206 source.n17 a_n3394_n3888# 2.55133f
C207 source.n18 a_n3394_n3888# 0.381571f
C208 source.t7 a_n3394_n3888# 0.290446f
C209 source.t3 a_n3394_n3888# 0.290446f
C210 source.n19 a_n3394_n3888# 2.55133f
C211 source.n20 a_n3394_n3888# 0.381571f
C212 source.t39 a_n3394_n3888# 0.290446f
C213 source.t2 a_n3394_n3888# 0.290446f
C214 source.n21 a_n3394_n3888# 2.55133f
C215 source.n22 a_n3394_n3888# 0.381571f
C216 source.t47 a_n3394_n3888# 3.25492f
C217 source.n23 a_n3394_n3888# 1.96945f
C218 source.t14 a_n3394_n3888# 3.25492f
C219 source.n24 a_n3394_n3888# 1.96945f
C220 source.t16 a_n3394_n3888# 0.290446f
C221 source.t17 a_n3394_n3888# 0.290446f
C222 source.n25 a_n3394_n3888# 2.55132f
C223 source.n26 a_n3394_n3888# 0.381574f
C224 source.t18 a_n3394_n3888# 0.290446f
C225 source.t36 a_n3394_n3888# 0.290446f
C226 source.n27 a_n3394_n3888# 2.55132f
C227 source.n28 a_n3394_n3888# 0.381574f
C228 source.t26 a_n3394_n3888# 0.290446f
C229 source.t27 a_n3394_n3888# 0.290446f
C230 source.n29 a_n3394_n3888# 2.55132f
C231 source.n30 a_n3394_n3888# 0.381574f
C232 source.t20 a_n3394_n3888# 0.290446f
C233 source.t21 a_n3394_n3888# 0.290446f
C234 source.n31 a_n3394_n3888# 2.55132f
C235 source.n32 a_n3394_n3888# 0.381574f
C236 source.t15 a_n3394_n3888# 0.290446f
C237 source.t32 a_n3394_n3888# 0.290446f
C238 source.n33 a_n3394_n3888# 2.55132f
C239 source.n34 a_n3394_n3888# 0.381574f
C240 source.t33 a_n3394_n3888# 3.25492f
C241 source.n35 a_n3394_n3888# 0.437094f
C242 source.t38 a_n3394_n3888# 3.25492f
C243 source.n36 a_n3394_n3888# 0.437094f
C244 source.t41 a_n3394_n3888# 0.290446f
C245 source.t40 a_n3394_n3888# 0.290446f
C246 source.n37 a_n3394_n3888# 2.55132f
C247 source.n38 a_n3394_n3888# 0.381574f
C248 source.t37 a_n3394_n3888# 0.290446f
C249 source.t43 a_n3394_n3888# 0.290446f
C250 source.n39 a_n3394_n3888# 2.55132f
C251 source.n40 a_n3394_n3888# 0.381574f
C252 source.t6 a_n3394_n3888# 0.290446f
C253 source.t12 a_n3394_n3888# 0.290446f
C254 source.n41 a_n3394_n3888# 2.55132f
C255 source.n42 a_n3394_n3888# 0.381574f
C256 source.t46 a_n3394_n3888# 0.290446f
C257 source.t44 a_n3394_n3888# 0.290446f
C258 source.n43 a_n3394_n3888# 2.55132f
C259 source.n44 a_n3394_n3888# 0.381574f
C260 source.t5 a_n3394_n3888# 0.290446f
C261 source.t8 a_n3394_n3888# 0.290446f
C262 source.n45 a_n3394_n3888# 2.55132f
C263 source.n46 a_n3394_n3888# 0.381574f
C264 source.t1 a_n3394_n3888# 3.25492f
C265 source.n47 a_n3394_n3888# 0.596929f
C266 source.n48 a_n3394_n3888# 1.80791f
C267 drain_left.t20 a_n3394_n3888# 0.323758f
C268 drain_left.t11 a_n3394_n3888# 0.323758f
C269 drain_left.n0 a_n3394_n3888# 2.93202f
C270 drain_left.t12 a_n3394_n3888# 0.323758f
C271 drain_left.t2 a_n3394_n3888# 0.323758f
C272 drain_left.n1 a_n3394_n3888# 2.92639f
C273 drain_left.n2 a_n3394_n3888# 0.765394f
C274 drain_left.t13 a_n3394_n3888# 0.323758f
C275 drain_left.t14 a_n3394_n3888# 0.323758f
C276 drain_left.n3 a_n3394_n3888# 2.92639f
C277 drain_left.n4 a_n3394_n3888# 0.337692f
C278 drain_left.t22 a_n3394_n3888# 0.323758f
C279 drain_left.t23 a_n3394_n3888# 0.323758f
C280 drain_left.n5 a_n3394_n3888# 2.93202f
C281 drain_left.t10 a_n3394_n3888# 0.323758f
C282 drain_left.t21 a_n3394_n3888# 0.323758f
C283 drain_left.n6 a_n3394_n3888# 2.92639f
C284 drain_left.n7 a_n3394_n3888# 0.765394f
C285 drain_left.t15 a_n3394_n3888# 0.323758f
C286 drain_left.t9 a_n3394_n3888# 0.323758f
C287 drain_left.n8 a_n3394_n3888# 2.92639f
C288 drain_left.n9 a_n3394_n3888# 0.337692f
C289 drain_left.n10 a_n3394_n3888# 1.99789f
C290 drain_left.t0 a_n3394_n3888# 0.323758f
C291 drain_left.t3 a_n3394_n3888# 0.323758f
C292 drain_left.n11 a_n3394_n3888# 2.93202f
C293 drain_left.t19 a_n3394_n3888# 0.323758f
C294 drain_left.t4 a_n3394_n3888# 0.323758f
C295 drain_left.n12 a_n3394_n3888# 2.9264f
C296 drain_left.n13 a_n3394_n3888# 0.765389f
C297 drain_left.t1 a_n3394_n3888# 0.323758f
C298 drain_left.t7 a_n3394_n3888# 0.323758f
C299 drain_left.n14 a_n3394_n3888# 2.9264f
C300 drain_left.n15 a_n3394_n3888# 0.380004f
C301 drain_left.t16 a_n3394_n3888# 0.323758f
C302 drain_left.t5 a_n3394_n3888# 0.323758f
C303 drain_left.n16 a_n3394_n3888# 2.9264f
C304 drain_left.n17 a_n3394_n3888# 0.380004f
C305 drain_left.t6 a_n3394_n3888# 0.323758f
C306 drain_left.t18 a_n3394_n3888# 0.323758f
C307 drain_left.n18 a_n3394_n3888# 2.9264f
C308 drain_left.n19 a_n3394_n3888# 0.380004f
C309 drain_left.t8 a_n3394_n3888# 0.323758f
C310 drain_left.t17 a_n3394_n3888# 0.323758f
C311 drain_left.n20 a_n3394_n3888# 2.92639f
C312 drain_left.n21 a_n3394_n3888# 0.621603f
C313 plus.n0 a_n3394_n3888# 0.039377f
C314 plus.t1 a_n3394_n3888# 1.17491f
C315 plus.t13 a_n3394_n3888# 1.17491f
C316 plus.n1 a_n3394_n3888# 0.039377f
C317 plus.t6 a_n3394_n3888# 1.17491f
C318 plus.n2 a_n3394_n3888# 0.453402f
C319 plus.n3 a_n3394_n3888# 0.039377f
C320 plus.t23 a_n3394_n3888# 1.17491f
C321 plus.t11 a_n3394_n3888# 1.17491f
C322 plus.n4 a_n3394_n3888# 0.453402f
C323 plus.n5 a_n3394_n3888# 0.039377f
C324 plus.t2 a_n3394_n3888# 1.17491f
C325 plus.t14 a_n3394_n3888# 1.17491f
C326 plus.n6 a_n3394_n3888# 0.453402f
C327 plus.n7 a_n3394_n3888# 0.039377f
C328 plus.t7 a_n3394_n3888# 1.17491f
C329 plus.t12 a_n3394_n3888# 1.17491f
C330 plus.n8 a_n3394_n3888# 0.453402f
C331 plus.n9 a_n3394_n3888# 0.039377f
C332 plus.t5 a_n3394_n3888# 1.17491f
C333 plus.t17 a_n3394_n3888# 1.17491f
C334 plus.n10 a_n3394_n3888# 0.46146f
C335 plus.t8 a_n3394_n3888# 1.1949f
C336 plus.n11 a_n3394_n3888# 0.435513f
C337 plus.n12 a_n3394_n3888# 0.169518f
C338 plus.n13 a_n3394_n3888# 0.008935f
C339 plus.n14 a_n3394_n3888# 0.453402f
C340 plus.n15 a_n3394_n3888# 0.008935f
C341 plus.n16 a_n3394_n3888# 0.039377f
C342 plus.n17 a_n3394_n3888# 0.039377f
C343 plus.n18 a_n3394_n3888# 0.039377f
C344 plus.n19 a_n3394_n3888# 0.008935f
C345 plus.n20 a_n3394_n3888# 0.453402f
C346 plus.n21 a_n3394_n3888# 0.008935f
C347 plus.n22 a_n3394_n3888# 0.039377f
C348 plus.n23 a_n3394_n3888# 0.039377f
C349 plus.n24 a_n3394_n3888# 0.039377f
C350 plus.n25 a_n3394_n3888# 0.008935f
C351 plus.n26 a_n3394_n3888# 0.453402f
C352 plus.n27 a_n3394_n3888# 0.008935f
C353 plus.n28 a_n3394_n3888# 0.039377f
C354 plus.n29 a_n3394_n3888# 0.039377f
C355 plus.n30 a_n3394_n3888# 0.039377f
C356 plus.n31 a_n3394_n3888# 0.008935f
C357 plus.n32 a_n3394_n3888# 0.453402f
C358 plus.n33 a_n3394_n3888# 0.008935f
C359 plus.n34 a_n3394_n3888# 0.039377f
C360 plus.n35 a_n3394_n3888# 0.039377f
C361 plus.n36 a_n3394_n3888# 0.039377f
C362 plus.n37 a_n3394_n3888# 0.008935f
C363 plus.n38 a_n3394_n3888# 0.453402f
C364 plus.n39 a_n3394_n3888# 0.008935f
C365 plus.n40 a_n3394_n3888# 0.453766f
C366 plus.n41 a_n3394_n3888# 0.514088f
C367 plus.n42 a_n3394_n3888# 0.039377f
C368 plus.t22 a_n3394_n3888# 1.17491f
C369 plus.n43 a_n3394_n3888# 0.039377f
C370 plus.t20 a_n3394_n3888# 1.17491f
C371 plus.t19 a_n3394_n3888# 1.17491f
C372 plus.n44 a_n3394_n3888# 0.453402f
C373 plus.n45 a_n3394_n3888# 0.039377f
C374 plus.t18 a_n3394_n3888# 1.17491f
C375 plus.t0 a_n3394_n3888# 1.17491f
C376 plus.n46 a_n3394_n3888# 0.453402f
C377 plus.n47 a_n3394_n3888# 0.039377f
C378 plus.t10 a_n3394_n3888# 1.17491f
C379 plus.t9 a_n3394_n3888# 1.17491f
C380 plus.n48 a_n3394_n3888# 0.453402f
C381 plus.n49 a_n3394_n3888# 0.039377f
C382 plus.t16 a_n3394_n3888# 1.17491f
C383 plus.t15 a_n3394_n3888# 1.17491f
C384 plus.n50 a_n3394_n3888# 0.453402f
C385 plus.n51 a_n3394_n3888# 0.039377f
C386 plus.t21 a_n3394_n3888# 1.17491f
C387 plus.t4 a_n3394_n3888# 1.17491f
C388 plus.n52 a_n3394_n3888# 0.46146f
C389 plus.t3 a_n3394_n3888# 1.1949f
C390 plus.n53 a_n3394_n3888# 0.435513f
C391 plus.n54 a_n3394_n3888# 0.169518f
C392 plus.n55 a_n3394_n3888# 0.008935f
C393 plus.n56 a_n3394_n3888# 0.453402f
C394 plus.n57 a_n3394_n3888# 0.008935f
C395 plus.n58 a_n3394_n3888# 0.039377f
C396 plus.n59 a_n3394_n3888# 0.039377f
C397 plus.n60 a_n3394_n3888# 0.039377f
C398 plus.n61 a_n3394_n3888# 0.008935f
C399 plus.n62 a_n3394_n3888# 0.453402f
C400 plus.n63 a_n3394_n3888# 0.008935f
C401 plus.n64 a_n3394_n3888# 0.039377f
C402 plus.n65 a_n3394_n3888# 0.039377f
C403 plus.n66 a_n3394_n3888# 0.039377f
C404 plus.n67 a_n3394_n3888# 0.008935f
C405 plus.n68 a_n3394_n3888# 0.453402f
C406 plus.n69 a_n3394_n3888# 0.008935f
C407 plus.n70 a_n3394_n3888# 0.039377f
C408 plus.n71 a_n3394_n3888# 0.039377f
C409 plus.n72 a_n3394_n3888# 0.039377f
C410 plus.n73 a_n3394_n3888# 0.008935f
C411 plus.n74 a_n3394_n3888# 0.453402f
C412 plus.n75 a_n3394_n3888# 0.008935f
C413 plus.n76 a_n3394_n3888# 0.039377f
C414 plus.n77 a_n3394_n3888# 0.039377f
C415 plus.n78 a_n3394_n3888# 0.039377f
C416 plus.n79 a_n3394_n3888# 0.008935f
C417 plus.n80 a_n3394_n3888# 0.453402f
C418 plus.n81 a_n3394_n3888# 0.008935f
C419 plus.n82 a_n3394_n3888# 0.453766f
C420 plus.n83 a_n3394_n3888# 1.59258f
.ends

