* NGSPICE file created from diffpair216.ext - technology: sky130A

.subckt diffpair216 minus drain_right drain_left source plus
X0 drain_right.t13 minus.t0 source.t16 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X1 a_n2204_n1488# a_n2204_n1488# a_n2204_n1488# a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.6
X2 drain_left.t13 plus.t0 source.t9 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X3 source.t0 plus.t1 drain_left.t12 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X4 drain_right.t12 minus.t1 source.t25 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X5 source.t26 minus.t2 drain_right.t11 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X6 source.t8 plus.t2 drain_left.t11 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X7 drain_right.t10 minus.t3 source.t21 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X8 drain_right.t9 minus.t4 source.t24 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X9 source.t23 minus.t5 drain_right.t8 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X10 drain_left.t10 plus.t3 source.t11 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X11 drain_left.t9 plus.t4 source.t1 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X12 a_n2204_n1488# a_n2204_n1488# a_n2204_n1488# a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X13 drain_left.t8 plus.t5 source.t2 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X14 source.t13 minus.t6 drain_right.t7 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X15 drain_right.t6 minus.t7 source.t19 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X16 drain_right.t5 minus.t8 source.t15 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X17 source.t3 plus.t6 drain_left.t7 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X18 source.t7 plus.t7 drain_left.t6 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X19 source.t14 minus.t9 drain_right.t4 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X20 source.t17 minus.t10 drain_right.t3 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X21 source.t20 minus.t11 drain_right.t2 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X22 a_n2204_n1488# a_n2204_n1488# a_n2204_n1488# a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X23 drain_left.t5 plus.t8 source.t10 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X24 drain_right.t1 minus.t12 source.t22 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X25 drain_right.t0 minus.t13 source.t18 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X26 source.t4 plus.t9 drain_left.t4 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X27 drain_left.t3 plus.t10 source.t27 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X28 a_n2204_n1488# a_n2204_n1488# a_n2204_n1488# a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X29 drain_left.t2 plus.t11 source.t6 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X30 drain_left.t1 plus.t12 source.t12 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X31 source.t5 plus.t13 drain_left.t0 a_n2204_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
R0 minus.n5 minus.t12 209.819
R1 minus.n23 minus.t13 209.819
R2 minus.n4 minus.t9 185.972
R3 minus.n8 minus.t8 185.972
R4 minus.n9 minus.t6 185.972
R5 minus.n10 minus.t3 185.972
R6 minus.n14 minus.t5 185.972
R7 minus.n16 minus.t4 185.972
R8 minus.n22 minus.t2 185.972
R9 minus.n26 minus.t0 185.972
R10 minus.n27 minus.t11 185.972
R11 minus.n28 minus.t7 185.972
R12 minus.n32 minus.t10 185.972
R13 minus.n34 minus.t1 185.972
R14 minus.n17 minus.n16 161.3
R15 minus.n15 minus.n0 161.3
R16 minus.n14 minus.n13 161.3
R17 minus.n12 minus.n1 161.3
R18 minus.n11 minus.n10 161.3
R19 minus.n8 minus.n7 161.3
R20 minus.n6 minus.n3 161.3
R21 minus.n35 minus.n34 161.3
R22 minus.n33 minus.n18 161.3
R23 minus.n32 minus.n31 161.3
R24 minus.n30 minus.n19 161.3
R25 minus.n29 minus.n28 161.3
R26 minus.n26 minus.n25 161.3
R27 minus.n24 minus.n21 161.3
R28 minus.n9 minus.n2 80.6037
R29 minus.n27 minus.n20 80.6037
R30 minus.n9 minus.n8 48.2005
R31 minus.n10 minus.n9 48.2005
R32 minus.n27 minus.n26 48.2005
R33 minus.n28 minus.n27 48.2005
R34 minus.n4 minus.n3 45.2793
R35 minus.n14 minus.n1 45.2793
R36 minus.n22 minus.n21 45.2793
R37 minus.n32 minus.n19 45.2793
R38 minus.n6 minus.n5 44.9119
R39 minus.n24 minus.n23 44.9119
R40 minus.n16 minus.n15 35.055
R41 minus.n34 minus.n33 35.055
R42 minus.n36 minus.n17 30.7259
R43 minus.n5 minus.n4 17.739
R44 minus.n23 minus.n22 17.739
R45 minus.n15 minus.n14 13.146
R46 minus.n33 minus.n32 13.146
R47 minus.n36 minus.n35 6.57436
R48 minus.n8 minus.n3 2.92171
R49 minus.n10 minus.n1 2.92171
R50 minus.n26 minus.n21 2.92171
R51 minus.n28 minus.n19 2.92171
R52 minus.n11 minus.n2 0.285035
R53 minus.n7 minus.n2 0.285035
R54 minus.n25 minus.n20 0.285035
R55 minus.n29 minus.n20 0.285035
R56 minus.n17 minus.n0 0.189894
R57 minus.n13 minus.n0 0.189894
R58 minus.n13 minus.n12 0.189894
R59 minus.n12 minus.n11 0.189894
R60 minus.n7 minus.n6 0.189894
R61 minus.n25 minus.n24 0.189894
R62 minus.n30 minus.n29 0.189894
R63 minus.n31 minus.n30 0.189894
R64 minus.n31 minus.n18 0.189894
R65 minus.n35 minus.n18 0.189894
R66 minus minus.n36 0.188
R67 source.n0 source.t9 69.6943
R68 source.n7 source.t22 69.6943
R69 source.n27 source.t25 69.6942
R70 source.n20 source.t11 69.6942
R71 source.n2 source.n1 63.0943
R72 source.n4 source.n3 63.0943
R73 source.n6 source.n5 63.0943
R74 source.n9 source.n8 63.0943
R75 source.n11 source.n10 63.0943
R76 source.n13 source.n12 63.0943
R77 source.n26 source.n25 63.0942
R78 source.n24 source.n23 63.0942
R79 source.n22 source.n21 63.0942
R80 source.n19 source.n18 63.0942
R81 source.n17 source.n16 63.0942
R82 source.n15 source.n14 63.0942
R83 source.n15 source.n13 16.073
R84 source.n28 source.n0 9.60747
R85 source.n25 source.t19 6.6005
R86 source.n25 source.t17 6.6005
R87 source.n23 source.t16 6.6005
R88 source.n23 source.t20 6.6005
R89 source.n21 source.t18 6.6005
R90 source.n21 source.t26 6.6005
R91 source.n18 source.t6 6.6005
R92 source.n18 source.t5 6.6005
R93 source.n16 source.t1 6.6005
R94 source.n16 source.t3 6.6005
R95 source.n14 source.t12 6.6005
R96 source.n14 source.t8 6.6005
R97 source.n1 source.t2 6.6005
R98 source.n1 source.t0 6.6005
R99 source.n3 source.t10 6.6005
R100 source.n3 source.t7 6.6005
R101 source.n5 source.t27 6.6005
R102 source.n5 source.t4 6.6005
R103 source.n8 source.t15 6.6005
R104 source.n8 source.t14 6.6005
R105 source.n10 source.t21 6.6005
R106 source.n10 source.t13 6.6005
R107 source.n12 source.t24 6.6005
R108 source.n12 source.t23 6.6005
R109 source.n28 source.n27 5.66429
R110 source.n7 source.n6 0.87119
R111 source.n22 source.n20 0.87119
R112 source.n13 source.n11 0.802224
R113 source.n11 source.n9 0.802224
R114 source.n9 source.n7 0.802224
R115 source.n6 source.n4 0.802224
R116 source.n4 source.n2 0.802224
R117 source.n2 source.n0 0.802224
R118 source.n17 source.n15 0.802224
R119 source.n19 source.n17 0.802224
R120 source.n20 source.n19 0.802224
R121 source.n24 source.n22 0.802224
R122 source.n26 source.n24 0.802224
R123 source.n27 source.n26 0.802224
R124 source source.n28 0.188
R125 drain_right.n1 drain_right.t0 87.1747
R126 drain_right.n11 drain_right.t9 86.3731
R127 drain_right.n8 drain_right.n6 80.5748
R128 drain_right.n4 drain_right.n2 80.5747
R129 drain_right.n8 drain_right.n7 79.7731
R130 drain_right.n10 drain_right.n9 79.7731
R131 drain_right.n4 drain_right.n3 79.773
R132 drain_right.n1 drain_right.n0 79.773
R133 drain_right drain_right.n5 24.6056
R134 drain_right.n2 drain_right.t3 6.6005
R135 drain_right.n2 drain_right.t12 6.6005
R136 drain_right.n3 drain_right.t2 6.6005
R137 drain_right.n3 drain_right.t6 6.6005
R138 drain_right.n0 drain_right.t11 6.6005
R139 drain_right.n0 drain_right.t13 6.6005
R140 drain_right.n6 drain_right.t4 6.6005
R141 drain_right.n6 drain_right.t1 6.6005
R142 drain_right.n7 drain_right.t7 6.6005
R143 drain_right.n7 drain_right.t5 6.6005
R144 drain_right.n9 drain_right.t8 6.6005
R145 drain_right.n9 drain_right.t10 6.6005
R146 drain_right drain_right.n11 6.05408
R147 drain_right.n11 drain_right.n10 0.802224
R148 drain_right.n10 drain_right.n8 0.802224
R149 drain_right.n5 drain_right.n1 0.546447
R150 drain_right.n5 drain_right.n4 0.145585
R151 plus.n5 plus.t10 209.819
R152 plus.n23 plus.t3 209.819
R153 plus.n16 plus.t0 185.972
R154 plus.n14 plus.t1 185.972
R155 plus.n2 plus.t5 185.972
R156 plus.n9 plus.t7 185.972
R157 plus.n8 plus.t8 185.972
R158 plus.n4 plus.t9 185.972
R159 plus.n34 plus.t12 185.972
R160 plus.n32 plus.t2 185.972
R161 plus.n20 plus.t4 185.972
R162 plus.n27 plus.t6 185.972
R163 plus.n26 plus.t11 185.972
R164 plus.n22 plus.t13 185.972
R165 plus.n7 plus.n6 161.3
R166 plus.n8 plus.n3 161.3
R167 plus.n11 plus.n2 161.3
R168 plus.n13 plus.n12 161.3
R169 plus.n14 plus.n1 161.3
R170 plus.n15 plus.n0 161.3
R171 plus.n17 plus.n16 161.3
R172 plus.n25 plus.n24 161.3
R173 plus.n26 plus.n21 161.3
R174 plus.n29 plus.n20 161.3
R175 plus.n31 plus.n30 161.3
R176 plus.n32 plus.n19 161.3
R177 plus.n33 plus.n18 161.3
R178 plus.n35 plus.n34 161.3
R179 plus.n10 plus.n9 80.6037
R180 plus.n28 plus.n27 80.6037
R181 plus.n9 plus.n2 48.2005
R182 plus.n9 plus.n8 48.2005
R183 plus.n27 plus.n20 48.2005
R184 plus.n27 plus.n26 48.2005
R185 plus.n14 plus.n13 45.2793
R186 plus.n7 plus.n4 45.2793
R187 plus.n32 plus.n31 45.2793
R188 plus.n25 plus.n22 45.2793
R189 plus.n24 plus.n23 44.9119
R190 plus.n6 plus.n5 44.9119
R191 plus.n16 plus.n15 35.055
R192 plus.n34 plus.n33 35.055
R193 plus plus.n35 28.0161
R194 plus.n23 plus.n22 17.739
R195 plus.n5 plus.n4 17.739
R196 plus.n15 plus.n14 13.146
R197 plus.n33 plus.n32 13.146
R198 plus plus.n17 8.80921
R199 plus.n13 plus.n2 2.92171
R200 plus.n8 plus.n7 2.92171
R201 plus.n31 plus.n20 2.92171
R202 plus.n26 plus.n25 2.92171
R203 plus.n10 plus.n3 0.285035
R204 plus.n11 plus.n10 0.285035
R205 plus.n29 plus.n28 0.285035
R206 plus.n28 plus.n21 0.285035
R207 plus.n6 plus.n3 0.189894
R208 plus.n12 plus.n11 0.189894
R209 plus.n12 plus.n1 0.189894
R210 plus.n1 plus.n0 0.189894
R211 plus.n17 plus.n0 0.189894
R212 plus.n35 plus.n18 0.189894
R213 plus.n19 plus.n18 0.189894
R214 plus.n30 plus.n19 0.189894
R215 plus.n30 plus.n29 0.189894
R216 plus.n24 plus.n21 0.189894
R217 drain_left.n7 drain_left.t3 87.1748
R218 drain_left.n1 drain_left.t1 87.1747
R219 drain_left.n4 drain_left.n2 80.5747
R220 drain_left.n11 drain_left.n10 79.7731
R221 drain_left.n9 drain_left.n8 79.7731
R222 drain_left.n7 drain_left.n6 79.7731
R223 drain_left.n4 drain_left.n3 79.773
R224 drain_left.n1 drain_left.n0 79.773
R225 drain_left drain_left.n5 25.1588
R226 drain_left.n2 drain_left.t0 6.6005
R227 drain_left.n2 drain_left.t10 6.6005
R228 drain_left.n3 drain_left.t7 6.6005
R229 drain_left.n3 drain_left.t2 6.6005
R230 drain_left.n0 drain_left.t11 6.6005
R231 drain_left.n0 drain_left.t9 6.6005
R232 drain_left.n10 drain_left.t12 6.6005
R233 drain_left.n10 drain_left.t13 6.6005
R234 drain_left.n8 drain_left.t6 6.6005
R235 drain_left.n8 drain_left.t8 6.6005
R236 drain_left.n6 drain_left.t4 6.6005
R237 drain_left.n6 drain_left.t5 6.6005
R238 drain_left drain_left.n11 6.45494
R239 drain_left.n9 drain_left.n7 0.802224
R240 drain_left.n11 drain_left.n9 0.802224
R241 drain_left.n5 drain_left.n1 0.546447
R242 drain_left.n5 drain_left.n4 0.145585
C0 drain_right minus 2.46507f
C1 source drain_right 7.30952f
C2 drain_left drain_right 1.14527f
C3 source minus 2.83304f
C4 drain_left minus 0.178018f
C5 source drain_left 7.31078f
C6 drain_right plus 0.378841f
C7 plus minus 4.23822f
C8 source plus 2.84717f
C9 drain_left plus 2.68089f
C10 drain_right a_n2204_n1488# 4.85671f
C11 drain_left a_n2204_n1488# 5.19847f
C12 source a_n2204_n1488# 3.117502f
C13 minus a_n2204_n1488# 7.985787f
C14 plus a_n2204_n1488# 9.28651f
C15 drain_left.t1 a_n2204_n1488# 0.573659f
C16 drain_left.t11 a_n2204_n1488# 0.06165f
C17 drain_left.t9 a_n2204_n1488# 0.06165f
C18 drain_left.n0 a_n2204_n1488# 0.444617f
C19 drain_left.n1 a_n2204_n1488# 0.647119f
C20 drain_left.t0 a_n2204_n1488# 0.06165f
C21 drain_left.t10 a_n2204_n1488# 0.06165f
C22 drain_left.n2 a_n2204_n1488# 0.44813f
C23 drain_left.t7 a_n2204_n1488# 0.06165f
C24 drain_left.t2 a_n2204_n1488# 0.06165f
C25 drain_left.n3 a_n2204_n1488# 0.444617f
C26 drain_left.n4 a_n2204_n1488# 0.641153f
C27 drain_left.n5 a_n2204_n1488# 0.896484f
C28 drain_left.t3 a_n2204_n1488# 0.573661f
C29 drain_left.t4 a_n2204_n1488# 0.06165f
C30 drain_left.t5 a_n2204_n1488# 0.06165f
C31 drain_left.n6 a_n2204_n1488# 0.444619f
C32 drain_left.n7 a_n2204_n1488# 0.667444f
C33 drain_left.t6 a_n2204_n1488# 0.06165f
C34 drain_left.t8 a_n2204_n1488# 0.06165f
C35 drain_left.n8 a_n2204_n1488# 0.444619f
C36 drain_left.n9 a_n2204_n1488# 0.342527f
C37 drain_left.t12 a_n2204_n1488# 0.06165f
C38 drain_left.t13 a_n2204_n1488# 0.06165f
C39 drain_left.n10 a_n2204_n1488# 0.444619f
C40 drain_left.n11 a_n2204_n1488# 0.569291f
C41 plus.n0 a_n2204_n1488# 0.046053f
C42 plus.t0 a_n2204_n1488# 0.248571f
C43 plus.t1 a_n2204_n1488# 0.248571f
C44 plus.n1 a_n2204_n1488# 0.046053f
C45 plus.t5 a_n2204_n1488# 0.248571f
C46 plus.n2 a_n2204_n1488# 0.147565f
C47 plus.n3 a_n2204_n1488# 0.061451f
C48 plus.t7 a_n2204_n1488# 0.248571f
C49 plus.t8 a_n2204_n1488# 0.248571f
C50 plus.t9 a_n2204_n1488# 0.248571f
C51 plus.n4 a_n2204_n1488# 0.154689f
C52 plus.t10 a_n2204_n1488# 0.265186f
C53 plus.n5 a_n2204_n1488# 0.133488f
C54 plus.n6 a_n2204_n1488# 0.188406f
C55 plus.n7 a_n2204_n1488# 0.01045f
C56 plus.n8 a_n2204_n1488# 0.147565f
C57 plus.n9 a_n2204_n1488# 0.157447f
C58 plus.n10 a_n2204_n1488# 0.061308f
C59 plus.n11 a_n2204_n1488# 0.061451f
C60 plus.n12 a_n2204_n1488# 0.046053f
C61 plus.n13 a_n2204_n1488# 0.01045f
C62 plus.n14 a_n2204_n1488# 0.148984f
C63 plus.n15 a_n2204_n1488# 0.01045f
C64 plus.n16 a_n2204_n1488# 0.144441f
C65 plus.n17 a_n2204_n1488# 0.352474f
C66 plus.n18 a_n2204_n1488# 0.046053f
C67 plus.t12 a_n2204_n1488# 0.248571f
C68 plus.n19 a_n2204_n1488# 0.046053f
C69 plus.t2 a_n2204_n1488# 0.248571f
C70 plus.t4 a_n2204_n1488# 0.248571f
C71 plus.n20 a_n2204_n1488# 0.147565f
C72 plus.n21 a_n2204_n1488# 0.061451f
C73 plus.t6 a_n2204_n1488# 0.248571f
C74 plus.t11 a_n2204_n1488# 0.248571f
C75 plus.t13 a_n2204_n1488# 0.248571f
C76 plus.n22 a_n2204_n1488# 0.154689f
C77 plus.t3 a_n2204_n1488# 0.265186f
C78 plus.n23 a_n2204_n1488# 0.133488f
C79 plus.n24 a_n2204_n1488# 0.188406f
C80 plus.n25 a_n2204_n1488# 0.01045f
C81 plus.n26 a_n2204_n1488# 0.147565f
C82 plus.n27 a_n2204_n1488# 0.157447f
C83 plus.n28 a_n2204_n1488# 0.061308f
C84 plus.n29 a_n2204_n1488# 0.061451f
C85 plus.n30 a_n2204_n1488# 0.046053f
C86 plus.n31 a_n2204_n1488# 0.01045f
C87 plus.n32 a_n2204_n1488# 0.148984f
C88 plus.n33 a_n2204_n1488# 0.01045f
C89 plus.n34 a_n2204_n1488# 0.144441f
C90 plus.n35 a_n2204_n1488# 1.17495f
C91 drain_right.t0 a_n2204_n1488# 0.567964f
C92 drain_right.t11 a_n2204_n1488# 0.061038f
C93 drain_right.t13 a_n2204_n1488# 0.061038f
C94 drain_right.n0 a_n2204_n1488# 0.440203f
C95 drain_right.n1 a_n2204_n1488# 0.640695f
C96 drain_right.t3 a_n2204_n1488# 0.061038f
C97 drain_right.t12 a_n2204_n1488# 0.061038f
C98 drain_right.n2 a_n2204_n1488# 0.44368f
C99 drain_right.t2 a_n2204_n1488# 0.061038f
C100 drain_right.t6 a_n2204_n1488# 0.061038f
C101 drain_right.n3 a_n2204_n1488# 0.440203f
C102 drain_right.n4 a_n2204_n1488# 0.634787f
C103 drain_right.n5 a_n2204_n1488# 0.836785f
C104 drain_right.t4 a_n2204_n1488# 0.061038f
C105 drain_right.t1 a_n2204_n1488# 0.061038f
C106 drain_right.n6 a_n2204_n1488# 0.443683f
C107 drain_right.t7 a_n2204_n1488# 0.061038f
C108 drain_right.t5 a_n2204_n1488# 0.061038f
C109 drain_right.n7 a_n2204_n1488# 0.440205f
C110 drain_right.n8 a_n2204_n1488# 0.685146f
C111 drain_right.t8 a_n2204_n1488# 0.061038f
C112 drain_right.t10 a_n2204_n1488# 0.061038f
C113 drain_right.n9 a_n2204_n1488# 0.440205f
C114 drain_right.n10 a_n2204_n1488# 0.339126f
C115 drain_right.t9 a_n2204_n1488# 0.56498f
C116 drain_right.n11 a_n2204_n1488# 0.555889f
C117 source.t9 a_n2204_n1488# 0.614803f
C118 source.n0 a_n2204_n1488# 0.884543f
C119 source.t2 a_n2204_n1488# 0.074039f
C120 source.t0 a_n2204_n1488# 0.074039f
C121 source.n1 a_n2204_n1488# 0.469447f
C122 source.n2 a_n2204_n1488# 0.43342f
C123 source.t10 a_n2204_n1488# 0.074039f
C124 source.t7 a_n2204_n1488# 0.074039f
C125 source.n3 a_n2204_n1488# 0.469447f
C126 source.n4 a_n2204_n1488# 0.43342f
C127 source.t27 a_n2204_n1488# 0.074039f
C128 source.t4 a_n2204_n1488# 0.074039f
C129 source.n5 a_n2204_n1488# 0.469447f
C130 source.n6 a_n2204_n1488# 0.44036f
C131 source.t22 a_n2204_n1488# 0.614803f
C132 source.n7 a_n2204_n1488# 0.496927f
C133 source.t15 a_n2204_n1488# 0.074039f
C134 source.t14 a_n2204_n1488# 0.074039f
C135 source.n8 a_n2204_n1488# 0.469447f
C136 source.n9 a_n2204_n1488# 0.43342f
C137 source.t21 a_n2204_n1488# 0.074039f
C138 source.t13 a_n2204_n1488# 0.074039f
C139 source.n10 a_n2204_n1488# 0.469447f
C140 source.n11 a_n2204_n1488# 0.43342f
C141 source.t24 a_n2204_n1488# 0.074039f
C142 source.t23 a_n2204_n1488# 0.074039f
C143 source.n12 a_n2204_n1488# 0.469447f
C144 source.n13 a_n2204_n1488# 1.2405f
C145 source.t12 a_n2204_n1488# 0.074039f
C146 source.t8 a_n2204_n1488# 0.074039f
C147 source.n14 a_n2204_n1488# 0.469444f
C148 source.n15 a_n2204_n1488# 1.2405f
C149 source.t1 a_n2204_n1488# 0.074039f
C150 source.t3 a_n2204_n1488# 0.074039f
C151 source.n16 a_n2204_n1488# 0.469444f
C152 source.n17 a_n2204_n1488# 0.433423f
C153 source.t6 a_n2204_n1488# 0.074039f
C154 source.t5 a_n2204_n1488# 0.074039f
C155 source.n18 a_n2204_n1488# 0.469444f
C156 source.n19 a_n2204_n1488# 0.433423f
C157 source.t11 a_n2204_n1488# 0.6148f
C158 source.n20 a_n2204_n1488# 0.49693f
C159 source.t18 a_n2204_n1488# 0.074039f
C160 source.t26 a_n2204_n1488# 0.074039f
C161 source.n21 a_n2204_n1488# 0.469444f
C162 source.n22 a_n2204_n1488# 0.440363f
C163 source.t16 a_n2204_n1488# 0.074039f
C164 source.t20 a_n2204_n1488# 0.074039f
C165 source.n23 a_n2204_n1488# 0.469444f
C166 source.n24 a_n2204_n1488# 0.433423f
C167 source.t19 a_n2204_n1488# 0.074039f
C168 source.t17 a_n2204_n1488# 0.074039f
C169 source.n25 a_n2204_n1488# 0.469444f
C170 source.n26 a_n2204_n1488# 0.433423f
C171 source.t25 a_n2204_n1488# 0.6148f
C172 source.n27 a_n2204_n1488# 0.653512f
C173 source.n28 a_n2204_n1488# 0.916938f
C174 minus.n0 a_n2204_n1488# 0.044674f
C175 minus.n1 a_n2204_n1488# 0.010137f
C176 minus.t5 a_n2204_n1488# 0.241131f
C177 minus.n2 a_n2204_n1488# 0.059472f
C178 minus.n3 a_n2204_n1488# 0.010137f
C179 minus.t8 a_n2204_n1488# 0.241131f
C180 minus.t12 a_n2204_n1488# 0.257248f
C181 minus.t9 a_n2204_n1488# 0.241131f
C182 minus.n4 a_n2204_n1488# 0.150059f
C183 minus.n5 a_n2204_n1488# 0.129492f
C184 minus.n6 a_n2204_n1488# 0.182767f
C185 minus.n7 a_n2204_n1488# 0.059612f
C186 minus.n8 a_n2204_n1488# 0.143148f
C187 minus.t6 a_n2204_n1488# 0.241131f
C188 minus.n9 a_n2204_n1488# 0.152734f
C189 minus.t3 a_n2204_n1488# 0.241131f
C190 minus.n10 a_n2204_n1488# 0.143148f
C191 minus.n11 a_n2204_n1488# 0.059612f
C192 minus.n12 a_n2204_n1488# 0.044674f
C193 minus.n13 a_n2204_n1488# 0.044674f
C194 minus.n14 a_n2204_n1488# 0.144525f
C195 minus.n15 a_n2204_n1488# 0.010137f
C196 minus.t4 a_n2204_n1488# 0.241131f
C197 minus.n16 a_n2204_n1488# 0.140118f
C198 minus.n17 a_n2204_n1488# 1.21331f
C199 minus.n18 a_n2204_n1488# 0.044674f
C200 minus.n19 a_n2204_n1488# 0.010137f
C201 minus.n20 a_n2204_n1488# 0.059472f
C202 minus.n21 a_n2204_n1488# 0.010137f
C203 minus.t13 a_n2204_n1488# 0.257248f
C204 minus.t2 a_n2204_n1488# 0.241131f
C205 minus.n22 a_n2204_n1488# 0.150059f
C206 minus.n23 a_n2204_n1488# 0.129492f
C207 minus.n24 a_n2204_n1488# 0.182767f
C208 minus.n25 a_n2204_n1488# 0.059612f
C209 minus.t0 a_n2204_n1488# 0.241131f
C210 minus.n26 a_n2204_n1488# 0.143148f
C211 minus.t11 a_n2204_n1488# 0.241131f
C212 minus.n27 a_n2204_n1488# 0.152734f
C213 minus.t7 a_n2204_n1488# 0.241131f
C214 minus.n28 a_n2204_n1488# 0.143148f
C215 minus.n29 a_n2204_n1488# 0.059612f
C216 minus.n30 a_n2204_n1488# 0.044674f
C217 minus.n31 a_n2204_n1488# 0.044674f
C218 minus.t10 a_n2204_n1488# 0.241131f
C219 minus.n32 a_n2204_n1488# 0.144525f
C220 minus.n33 a_n2204_n1488# 0.010137f
C221 minus.t1 a_n2204_n1488# 0.241131f
C222 minus.n34 a_n2204_n1488# 0.140118f
C223 minus.n35 a_n2204_n1488# 0.299867f
C224 minus.n36 a_n2204_n1488# 1.49117f
.ends

