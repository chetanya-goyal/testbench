* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t9 plus.t0 source.t16 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X1 a_n1496_n1288# a_n1496_n1288# a_n1496_n1288# a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=7.6 ps=39.6 w=2 l=0.15
X2 drain_right.t9 minus.t0 source.t2 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X3 drain_right.t8 minus.t1 source.t4 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X4 source.t14 plus.t1 drain_left.t8 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X5 drain_left.t7 plus.t2 source.t12 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X6 a_n1496_n1288# a_n1496_n1288# a_n1496_n1288# a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X7 a_n1496_n1288# a_n1496_n1288# a_n1496_n1288# a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X8 a_n1496_n1288# a_n1496_n1288# a_n1496_n1288# a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X9 source.t5 minus.t2 drain_right.t7 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X10 source.t0 minus.t3 drain_right.t6 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X11 drain_right.t5 minus.t4 source.t1 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X12 drain_right.t4 minus.t5 source.t6 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X13 drain_right.t3 minus.t6 source.t17 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X14 source.t18 minus.t7 drain_right.t2 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X15 source.t19 minus.t8 drain_right.t1 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X16 source.t13 plus.t3 drain_left.t6 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X17 drain_left.t5 plus.t4 source.t11 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X18 drain_right.t0 minus.t9 source.t3 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X19 source.t8 plus.t5 drain_left.t4 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X20 drain_left.t3 plus.t6 source.t15 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X21 drain_left.t2 plus.t7 source.t10 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X22 source.t9 plus.t8 drain_left.t1 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.15
X23 drain_left.t0 plus.t9 source.t7 a_n1496_n1288# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
R0 plus.n3 plus.t4 574.019
R1 plus.n9 plus.t9 574.019
R2 plus.n14 plus.t6 574.019
R3 plus.n20 plus.t0 574.019
R4 plus.n6 plus.t7 530.201
R5 plus.n2 plus.t8 530.201
R6 plus.n8 plus.t5 530.201
R7 plus.n17 plus.t2 530.201
R8 plus.n13 plus.t3 530.201
R9 plus.n19 plus.t1 530.201
R10 plus.n4 plus.n3 161.489
R11 plus.n15 plus.n14 161.489
R12 plus.n4 plus.n1 161.3
R13 plus.n6 plus.n5 161.3
R14 plus.n7 plus.n0 161.3
R15 plus.n10 plus.n9 161.3
R16 plus.n15 plus.n12 161.3
R17 plus.n17 plus.n16 161.3
R18 plus.n18 plus.n11 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n6 plus.n1 73.0308
R21 plus.n7 plus.n6 73.0308
R22 plus.n18 plus.n17 73.0308
R23 plus.n17 plus.n12 73.0308
R24 plus.n3 plus.n2 51.1217
R25 plus.n9 plus.n8 51.1217
R26 plus.n20 plus.n19 51.1217
R27 plus.n14 plus.n13 51.1217
R28 plus plus.n21 24.8949
R29 plus.n2 plus.n1 21.9096
R30 plus.n8 plus.n7 21.9096
R31 plus.n19 plus.n18 21.9096
R32 plus.n13 plus.n12 21.9096
R33 plus plus.n10 8.36982
R34 plus.n5 plus.n4 0.189894
R35 plus.n5 plus.n0 0.189894
R36 plus.n10 plus.n0 0.189894
R37 plus.n21 plus.n11 0.189894
R38 plus.n16 plus.n11 0.189894
R39 plus.n16 plus.n15 0.189894
R40 source.n0 source.t7 99.1169
R41 source.n5 source.t6 99.1169
R42 source.n19 source.t2 99.1168
R43 source.n14 source.t15 99.1168
R44 source.n2 source.n1 84.1169
R45 source.n4 source.n3 84.1169
R46 source.n7 source.n6 84.1169
R47 source.n9 source.n8 84.1169
R48 source.n18 source.n17 84.1168
R49 source.n16 source.n15 84.1168
R50 source.n13 source.n12 84.1168
R51 source.n11 source.n10 84.1168
R52 source.n17 source.t1 15.0005
R53 source.n17 source.t5 15.0005
R54 source.n15 source.t4 15.0005
R55 source.n15 source.t19 15.0005
R56 source.n12 source.t12 15.0005
R57 source.n12 source.t13 15.0005
R58 source.n10 source.t16 15.0005
R59 source.n10 source.t14 15.0005
R60 source.n1 source.t10 15.0005
R61 source.n1 source.t8 15.0005
R62 source.n3 source.t11 15.0005
R63 source.n3 source.t9 15.0005
R64 source.n6 source.t3 15.0005
R65 source.n6 source.t0 15.0005
R66 source.n8 source.t17 15.0005
R67 source.n8 source.t18 15.0005
R68 source.n11 source.n9 14.8327
R69 source.n20 source.n0 8.72921
R70 source.n20 source.n19 5.5436
R71 source.n5 source.n4 0.7505
R72 source.n16 source.n14 0.7505
R73 source.n9 source.n7 0.560845
R74 source.n7 source.n5 0.560845
R75 source.n4 source.n2 0.560845
R76 source.n2 source.n0 0.560845
R77 source.n13 source.n11 0.560845
R78 source.n14 source.n13 0.560845
R79 source.n18 source.n16 0.560845
R80 source.n19 source.n18 0.560845
R81 source source.n20 0.188
R82 drain_left.n5 drain_left.t5 116.356
R83 drain_left.n1 drain_left.t9 116.356
R84 drain_left.n3 drain_left.n2 101.16
R85 drain_left.n7 drain_left.n6 100.796
R86 drain_left.n5 drain_left.n4 100.796
R87 drain_left.n1 drain_left.n0 100.796
R88 drain_left drain_left.n3 22.1728
R89 drain_left.n2 drain_left.t6 15.0005
R90 drain_left.n2 drain_left.t3 15.0005
R91 drain_left.n0 drain_left.t8 15.0005
R92 drain_left.n0 drain_left.t7 15.0005
R93 drain_left.n6 drain_left.t4 15.0005
R94 drain_left.n6 drain_left.t0 15.0005
R95 drain_left.n4 drain_left.t1 15.0005
R96 drain_left.n4 drain_left.t2 15.0005
R97 drain_left drain_left.n7 6.21356
R98 drain_left.n7 drain_left.n5 0.560845
R99 drain_left.n3 drain_left.n1 0.0852402
R100 minus.n9 minus.t6 574.019
R101 minus.n3 minus.t5 574.019
R102 minus.n20 minus.t0 574.019
R103 minus.n14 minus.t1 574.019
R104 minus.n6 minus.t9 530.201
R105 minus.n8 minus.t7 530.201
R106 minus.n2 minus.t3 530.201
R107 minus.n17 minus.t4 530.201
R108 minus.n19 minus.t2 530.201
R109 minus.n13 minus.t8 530.201
R110 minus.n4 minus.n3 161.489
R111 minus.n15 minus.n14 161.489
R112 minus.n10 minus.n9 161.3
R113 minus.n7 minus.n0 161.3
R114 minus.n6 minus.n5 161.3
R115 minus.n4 minus.n1 161.3
R116 minus.n21 minus.n20 161.3
R117 minus.n18 minus.n11 161.3
R118 minus.n17 minus.n16 161.3
R119 minus.n15 minus.n12 161.3
R120 minus.n7 minus.n6 73.0308
R121 minus.n6 minus.n1 73.0308
R122 minus.n17 minus.n12 73.0308
R123 minus.n18 minus.n17 73.0308
R124 minus.n9 minus.n8 51.1217
R125 minus.n3 minus.n2 51.1217
R126 minus.n14 minus.n13 51.1217
R127 minus.n20 minus.n19 51.1217
R128 minus.n22 minus.n10 27.2259
R129 minus.n8 minus.n7 21.9096
R130 minus.n2 minus.n1 21.9096
R131 minus.n13 minus.n12 21.9096
R132 minus.n19 minus.n18 21.9096
R133 minus.n22 minus.n21 6.51376
R134 minus.n10 minus.n0 0.189894
R135 minus.n5 minus.n0 0.189894
R136 minus.n5 minus.n4 0.189894
R137 minus.n16 minus.n15 0.189894
R138 minus.n16 minus.n11 0.189894
R139 minus.n21 minus.n11 0.189894
R140 minus minus.n22 0.188
R141 drain_right.n1 drain_right.t8 116.356
R142 drain_right.n7 drain_right.t3 115.796
R143 drain_right.n6 drain_right.n4 101.356
R144 drain_right.n3 drain_right.n2 101.16
R145 drain_right.n6 drain_right.n5 100.796
R146 drain_right.n1 drain_right.n0 100.796
R147 drain_right drain_right.n3 21.6196
R148 drain_right.n2 drain_right.t7 15.0005
R149 drain_right.n2 drain_right.t9 15.0005
R150 drain_right.n0 drain_right.t1 15.0005
R151 drain_right.n0 drain_right.t5 15.0005
R152 drain_right.n4 drain_right.t6 15.0005
R153 drain_right.n4 drain_right.t4 15.0005
R154 drain_right.n5 drain_right.t2 15.0005
R155 drain_right.n5 drain_right.t0 15.0005
R156 drain_right drain_right.n7 5.93339
R157 drain_right.n7 drain_right.n6 0.560845
R158 drain_right.n3 drain_right.n1 0.0852402
C0 source minus 0.792553f
C1 drain_right source 5.39492f
C2 plus drain_left 0.880843f
C3 drain_right minus 0.738362f
C4 source plus 0.806624f
C5 plus minus 3.15945f
C6 drain_right plus 0.303657f
C7 source drain_left 5.39769f
C8 minus drain_left 0.176976f
C9 drain_right drain_left 0.732647f
C10 drain_right a_n1496_n1288# 3.48928f
C11 drain_left a_n1496_n1288# 3.70086f
C12 source a_n1496_n1288# 2.496369f
C13 minus a_n1496_n1288# 4.707685f
C14 plus a_n1496_n1288# 5.52328f
C15 drain_right.t8 a_n1496_n1288# 0.316501f
C16 drain_right.t1 a_n1496_n1288# 0.053456f
C17 drain_right.t5 a_n1496_n1288# 0.053456f
C18 drain_right.n0 a_n1496_n1288# 0.257994f
C19 drain_right.n1 a_n1496_n1288# 0.481234f
C20 drain_right.t7 a_n1496_n1288# 0.053456f
C21 drain_right.t9 a_n1496_n1288# 0.053456f
C22 drain_right.n2 a_n1496_n1288# 0.258888f
C23 drain_right.n3 a_n1496_n1288# 0.761596f
C24 drain_right.t6 a_n1496_n1288# 0.053456f
C25 drain_right.t4 a_n1496_n1288# 0.053456f
C26 drain_right.n4 a_n1496_n1288# 0.259435f
C27 drain_right.t2 a_n1496_n1288# 0.053456f
C28 drain_right.t0 a_n1496_n1288# 0.053456f
C29 drain_right.n5 a_n1496_n1288# 0.257995f
C30 drain_right.n6 a_n1496_n1288# 0.510488f
C31 drain_right.t3 a_n1496_n1288# 0.315254f
C32 drain_right.n7 a_n1496_n1288# 0.446299f
C33 minus.n0 a_n1496_n1288# 0.037606f
C34 minus.t6 a_n1496_n1288# 0.035322f
C35 minus.t7 a_n1496_n1288# 0.033198f
C36 minus.t9 a_n1496_n1288# 0.033198f
C37 minus.n1 a_n1496_n1288# 0.015953f
C38 minus.t3 a_n1496_n1288# 0.033198f
C39 minus.n2 a_n1496_n1288# 0.028982f
C40 minus.t5 a_n1496_n1288# 0.035322f
C41 minus.n3 a_n1496_n1288# 0.041703f
C42 minus.n4 a_n1496_n1288# 0.080958f
C43 minus.n5 a_n1496_n1288# 0.037606f
C44 minus.n6 a_n1496_n1288# 0.041457f
C45 minus.n7 a_n1496_n1288# 0.015953f
C46 minus.n8 a_n1496_n1288# 0.028982f
C47 minus.n9 a_n1496_n1288# 0.041652f
C48 minus.n10 a_n1496_n1288# 0.825914f
C49 minus.n11 a_n1496_n1288# 0.037606f
C50 minus.t2 a_n1496_n1288# 0.033198f
C51 minus.t4 a_n1496_n1288# 0.033198f
C52 minus.n12 a_n1496_n1288# 0.015953f
C53 minus.t1 a_n1496_n1288# 0.035322f
C54 minus.t8 a_n1496_n1288# 0.033198f
C55 minus.n13 a_n1496_n1288# 0.028982f
C56 minus.n14 a_n1496_n1288# 0.041703f
C57 minus.n15 a_n1496_n1288# 0.080958f
C58 minus.n16 a_n1496_n1288# 0.037606f
C59 minus.n17 a_n1496_n1288# 0.041457f
C60 minus.n18 a_n1496_n1288# 0.015953f
C61 minus.n19 a_n1496_n1288# 0.028982f
C62 minus.t0 a_n1496_n1288# 0.035322f
C63 minus.n20 a_n1496_n1288# 0.041652f
C64 minus.n21 a_n1496_n1288# 0.247077f
C65 minus.n22 a_n1496_n1288# 1.02014f
C66 drain_left.t9 a_n1496_n1288# 0.311465f
C67 drain_left.t8 a_n1496_n1288# 0.052605f
C68 drain_left.t7 a_n1496_n1288# 0.052605f
C69 drain_left.n0 a_n1496_n1288# 0.253888f
C70 drain_left.n1 a_n1496_n1288# 0.473575f
C71 drain_left.t6 a_n1496_n1288# 0.052605f
C72 drain_left.t3 a_n1496_n1288# 0.052605f
C73 drain_left.n2 a_n1496_n1288# 0.254768f
C74 drain_left.n3 a_n1496_n1288# 0.792664f
C75 drain_left.t5 a_n1496_n1288# 0.311465f
C76 drain_left.t1 a_n1496_n1288# 0.052605f
C77 drain_left.t2 a_n1496_n1288# 0.052605f
C78 drain_left.n4 a_n1496_n1288# 0.253889f
C79 drain_left.n5 a_n1496_n1288# 0.501229f
C80 drain_left.t4 a_n1496_n1288# 0.052605f
C81 drain_left.t0 a_n1496_n1288# 0.052605f
C82 drain_left.n6 a_n1496_n1288# 0.253889f
C83 drain_left.n7 a_n1496_n1288# 0.430921f
C84 source.t7 a_n1496_n1288# 0.337814f
C85 source.n0 a_n1496_n1288# 0.643864f
C86 source.t10 a_n1496_n1288# 0.064341f
C87 source.t8 a_n1496_n1288# 0.064341f
C88 source.n1 a_n1496_n1288# 0.270767f
C89 source.n2 a_n1496_n1288# 0.305917f
C90 source.t11 a_n1496_n1288# 0.064341f
C91 source.t9 a_n1496_n1288# 0.064341f
C92 source.n3 a_n1496_n1288# 0.270767f
C93 source.n4 a_n1496_n1288# 0.322337f
C94 source.t6 a_n1496_n1288# 0.337813f
C95 source.n5 a_n1496_n1288# 0.371104f
C96 source.t3 a_n1496_n1288# 0.064341f
C97 source.t0 a_n1496_n1288# 0.064341f
C98 source.n6 a_n1496_n1288# 0.270767f
C99 source.n7 a_n1496_n1288# 0.305917f
C100 source.t17 a_n1496_n1288# 0.064341f
C101 source.t18 a_n1496_n1288# 0.064341f
C102 source.n8 a_n1496_n1288# 0.270767f
C103 source.n9 a_n1496_n1288# 0.89444f
C104 source.t16 a_n1496_n1288# 0.064341f
C105 source.t14 a_n1496_n1288# 0.064341f
C106 source.n10 a_n1496_n1288# 0.270766f
C107 source.n11 a_n1496_n1288# 0.894441f
C108 source.t12 a_n1496_n1288# 0.064341f
C109 source.t13 a_n1496_n1288# 0.064341f
C110 source.n12 a_n1496_n1288# 0.270766f
C111 source.n13 a_n1496_n1288# 0.305918f
C112 source.t15 a_n1496_n1288# 0.337812f
C113 source.n14 a_n1496_n1288# 0.371105f
C114 source.t4 a_n1496_n1288# 0.064341f
C115 source.t19 a_n1496_n1288# 0.064341f
C116 source.n15 a_n1496_n1288# 0.270766f
C117 source.n16 a_n1496_n1288# 0.322338f
C118 source.t1 a_n1496_n1288# 0.064341f
C119 source.t5 a_n1496_n1288# 0.064341f
C120 source.n17 a_n1496_n1288# 0.270766f
C121 source.n18 a_n1496_n1288# 0.305918f
C122 source.t2 a_n1496_n1288# 0.337812f
C123 source.n19 a_n1496_n1288# 0.499714f
C124 source.n20 a_n1496_n1288# 0.664923f
C125 plus.n0 a_n1496_n1288# 0.038521f
C126 plus.t5 a_n1496_n1288# 0.034006f
C127 plus.t7 a_n1496_n1288# 0.034006f
C128 plus.n1 a_n1496_n1288# 0.016341f
C129 plus.t4 a_n1496_n1288# 0.036181f
C130 plus.t8 a_n1496_n1288# 0.034006f
C131 plus.n2 a_n1496_n1288# 0.029688f
C132 plus.n3 a_n1496_n1288# 0.042718f
C133 plus.n4 a_n1496_n1288# 0.082928f
C134 plus.n5 a_n1496_n1288# 0.038521f
C135 plus.n6 a_n1496_n1288# 0.042467f
C136 plus.n7 a_n1496_n1288# 0.016341f
C137 plus.n8 a_n1496_n1288# 0.029688f
C138 plus.t9 a_n1496_n1288# 0.036181f
C139 plus.n9 a_n1496_n1288# 0.042666f
C140 plus.n10 a_n1496_n1288# 0.276702f
C141 plus.n11 a_n1496_n1288# 0.038521f
C142 plus.t0 a_n1496_n1288# 0.036181f
C143 plus.t1 a_n1496_n1288# 0.034006f
C144 plus.t2 a_n1496_n1288# 0.034006f
C145 plus.n12 a_n1496_n1288# 0.016341f
C146 plus.t3 a_n1496_n1288# 0.034006f
C147 plus.n13 a_n1496_n1288# 0.029688f
C148 plus.t6 a_n1496_n1288# 0.036181f
C149 plus.n14 a_n1496_n1288# 0.042718f
C150 plus.n15 a_n1496_n1288# 0.082928f
C151 plus.n16 a_n1496_n1288# 0.038521f
C152 plus.n17 a_n1496_n1288# 0.042467f
C153 plus.n18 a_n1496_n1288# 0.016341f
C154 plus.n19 a_n1496_n1288# 0.029688f
C155 plus.n20 a_n1496_n1288# 0.042666f
C156 plus.n21 a_n1496_n1288# 0.810776f
.ends

