* NGSPICE file created from diffpair350.ext - technology: sky130A

.subckt diffpair350 minus drain_right drain_left source plus
X0 drain_right.t1 minus.t0 source.t1 a_n968_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=3.51 ps=18.78 w=9 l=0.3
X1 drain_left.t1 plus.t0 source.t0 a_n968_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=3.51 ps=18.78 w=9 l=0.3
X2 drain_right.t0 minus.t1 source.t2 a_n968_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=3.51 ps=18.78 w=9 l=0.3
X3 a_n968_n2692# a_n968_n2692# a_n968_n2692# a_n968_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.3
X4 drain_left.t0 plus.t1 source.t3 a_n968_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=3.51 ps=18.78 w=9 l=0.3
X5 a_n968_n2692# a_n968_n2692# a_n968_n2692# a_n968_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X6 a_n968_n2692# a_n968_n2692# a_n968_n2692# a_n968_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X7 a_n968_n2692# a_n968_n2692# a_n968_n2692# a_n968_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
R0 minus.n0 minus.t0 1043.25
R1 minus.n0 minus.t1 1019.22
R2 minus minus.n0 0.188
R3 source.n1 source.t1 51.0588
R4 source.n3 source.t2 51.0586
R5 source.n2 source.t0 51.0586
R6 source.n0 source.t3 51.0586
R7 source.n2 source.n1 20.1164
R8 source.n4 source.n0 14.0388
R9 source.n4 source.n3 5.53498
R10 source.n1 source.n0 0.741879
R11 source.n3 source.n2 0.741879
R12 source source.n4 0.188
R13 drain_right drain_right.t0 93.0524
R14 drain_right drain_right.t1 73.6616
R15 plus plus.t0 1038.27
R16 plus plus.t1 1023.73
R17 drain_left drain_left.t1 93.6056
R18 drain_left drain_left.t0 73.9332
C0 drain_right source 5.61763f
C1 drain_left plus 1.23732f
C2 drain_right drain_left 0.425172f
C3 minus plus 3.80743f
C4 drain_right minus 1.15154f
C5 drain_right plus 0.243866f
C6 source drain_left 5.62436f
C7 source minus 0.708331f
C8 drain_left minus 0.171671f
C9 source plus 0.722859f
C10 drain_right a_n968_n2692# 5.39335f
C11 drain_left a_n968_n2692# 5.51641f
C12 source a_n968_n2692# 4.677018f
C13 minus a_n968_n2692# 3.470347f
C14 plus a_n968_n2692# 6.35688f
C15 drain_left.t1 a_n968_n2692# 1.70234f
C16 drain_left.t0 a_n968_n2692# 1.51367f
C17 plus.t1 a_n968_n2692# 0.370228f
C18 plus.t0 a_n968_n2692# 0.392328f
C19 drain_right.t0 a_n968_n2692# 1.71061f
C20 drain_right.t1 a_n968_n2692# 1.53302f
C21 source.t3 a_n968_n2692# 1.55962f
C22 source.n0 a_n968_n2692# 0.911074f
C23 source.t1 a_n968_n2692# 1.55963f
C24 source.n1 a_n968_n2692# 1.24606f
C25 source.t0 a_n968_n2692# 1.55962f
C26 source.n2 a_n968_n2692# 1.24606f
C27 source.t2 a_n968_n2692# 1.55962f
C28 source.n3 a_n968_n2692# 0.451661f
C29 source.n4 a_n968_n2692# 1.07203f
C30 minus.t0 a_n968_n2692# 0.39281f
C31 minus.t1 a_n968_n2692# 0.358538f
C32 minus.n0 a_n968_n2692# 3.0203f
.ends

