* NGSPICE file created from diffpair620.ext - technology: sky130A

.subckt diffpair620 minus drain_right drain_left source plus
X0 drain_right.t1 minus.t0 source.t1 a_n1128_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.7
X1 a_n1128_n4892# a_n1128_n4892# a_n1128_n4892# a_n1128_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.7
X2 a_n1128_n4892# a_n1128_n4892# a_n1128_n4892# a_n1128_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X3 drain_left.t1 plus.t0 source.t3 a_n1128_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.7
X4 drain_left.t0 plus.t1 source.t2 a_n1128_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.7
X5 drain_right.t0 minus.t1 source.t0 a_n1128_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.7
X6 a_n1128_n4892# a_n1128_n4892# a_n1128_n4892# a_n1128_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X7 a_n1128_n4892# a_n1128_n4892# a_n1128_n4892# a_n1128_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
R0 minus.n0 minus.t0 945.576
R1 minus.n0 minus.t1 912.606
R2 minus minus.n0 0.188
R3 source.n0 source.t2 44.1297
R4 source.n1 source.t1 44.1296
R5 source.n3 source.t0 44.1295
R6 source.n2 source.t3 44.1295
R7 source.n2 source.n1 29.1393
R8 source.n4 source.n0 22.5445
R9 source.n4 source.n3 5.7074
R10 source.n1 source.n0 0.914293
R11 source.n3 source.n2 0.914293
R12 source source.n4 0.188
R13 drain_right drain_right.t0 94.9739
R14 drain_right drain_right.t1 66.9051
R15 plus plus.t0 936.427
R16 plus plus.t1 921.28
R17 drain_left drain_left.t1 95.5271
R18 drain_left drain_left.t0 67.3491
C0 drain_right plus 0.262193f
C1 source drain_left 8.823791f
C2 source minus 2.30058f
C3 drain_left minus 0.171858f
C4 source plus 2.31545f
C5 drain_right source 8.81087f
C6 drain_left plus 3.27952f
C7 drain_right drain_left 0.464239f
C8 minus plus 6.02366f
C9 drain_right minus 3.17893f
C10 drain_right a_n1128_n4892# 9.00807f
C11 drain_left a_n1128_n4892# 9.17671f
C12 source a_n1128_n4892# 9.519788f
C13 minus a_n1128_n4892# 4.688766f
C14 plus a_n1128_n4892# 11.20306f
C15 drain_left.t1 a_n1128_n4892# 4.34409f
C16 drain_left.t0 a_n1128_n4892# 3.85724f
C17 plus.t1 a_n1128_n4892# 2.433f
C18 plus.t0 a_n1128_n4892# 2.48842f
C19 drain_right.t0 a_n1128_n4892# 4.31611f
C20 drain_right.t1 a_n1128_n4892# 3.84956f
C21 source.t2 a_n1128_n4892# 3.58574f
C22 source.n0 a_n1128_n4892# 1.56273f
C23 source.t1 a_n1128_n4892# 3.58575f
C24 source.n1 a_n1128_n4892# 1.98077f
C25 source.t3 a_n1128_n4892# 3.58573f
C26 source.n2 a_n1128_n4892# 1.98079f
C27 source.t0 a_n1128_n4892# 3.58573f
C28 source.n3 a_n1128_n4892# 0.496962f
C29 source.n4 a_n1128_n4892# 1.80239f
C30 minus.t0 a_n1128_n4892# 2.48621f
C31 minus.t1 a_n1128_n4892# 2.37038f
C32 minus.n0 a_n1128_n4892# 6.60668f
.ends

