* NGSPICE file created from diffpair81.ext - technology: sky130A

.subckt diffpair81 minus drain_right drain_left source plus
X0 drain_right.t3 minus.t0 source.t4 a_n1106_n1292# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X1 drain_right.t2 minus.t1 source.t7 a_n1106_n1292# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X2 source.t1 plus.t0 drain_left.t3 a_n1106_n1292# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X3 a_n1106_n1292# a_n1106_n1292# a_n1106_n1292# a_n1106_n1292# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=7.6 ps=39.6 w=2 l=0.15
X4 source.t2 plus.t1 drain_left.t2 a_n1106_n1292# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X5 drain_left.t1 plus.t2 source.t3 a_n1106_n1292# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X6 drain_left.t0 plus.t3 source.t0 a_n1106_n1292# sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.95 ps=4.95 w=2 l=0.15
X7 a_n1106_n1292# a_n1106_n1292# a_n1106_n1292# a_n1106_n1292# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X8 source.t6 minus.t2 drain_right.t1 a_n1106_n1292# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
X9 a_n1106_n1292# a_n1106_n1292# a_n1106_n1292# a_n1106_n1292# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X10 a_n1106_n1292# a_n1106_n1292# a_n1106_n1292# a_n1106_n1292# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X11 source.t5 minus.t3 drain_right.t0 a_n1106_n1292# sky130_fd_pr__nfet_01v8 ad=0.95 pd=4.95 as=0.5 ps=2.5 w=2 l=0.15
R0 minus.n0 minus.t3 577.67
R1 minus.n0 minus.t0 577.67
R2 minus.n1 minus.t1 577.67
R3 minus.n1 minus.t2 577.67
R4 minus.n2 minus.n0 187.073
R5 minus.n2 minus.n1 167.823
R6 minus minus.n2 0.188
R7 source.n0 source.t0 99.1169
R8 source.n1 source.t2 99.1169
R9 source.n2 source.t4 99.1169
R10 source.n3 source.t5 99.1169
R11 source.n7 source.t7 99.1168
R12 source.n6 source.t6 99.1168
R13 source.n5 source.t3 99.1168
R14 source.n4 source.t1 99.1168
R15 source.n4 source.n3 14.2875
R16 source.n8 source.n0 8.74436
R17 source.n8 source.n7 5.5436
R18 source.n3 source.n2 0.560845
R19 source.n1 source.n0 0.560845
R20 source.n5 source.n4 0.560845
R21 source.n7 source.n6 0.560845
R22 source.n2 source.n1 0.470328
R23 source.n6 source.n5 0.470328
R24 source source.n8 0.188
R25 drain_right drain_right.n0 121.169
R26 drain_right drain_right.n1 107.008
R27 drain_right.n0 drain_right.t1 15.0005
R28 drain_right.n0 drain_right.t2 15.0005
R29 drain_right.n1 drain_right.t0 15.0005
R30 drain_right.n1 drain_right.t3 15.0005
R31 plus.n0 plus.t1 577.67
R32 plus.n0 plus.t3 577.67
R33 plus.n1 plus.t2 577.67
R34 plus.n1 plus.t0 577.67
R35 plus plus.n1 184.743
R36 plus plus.n0 169.679
R37 drain_left drain_left.n0 121.722
R38 drain_left drain_left.n1 107.008
R39 drain_left.n0 drain_left.t3 15.0005
R40 drain_left.n0 drain_left.t1 15.0005
R41 drain_left.n1 drain_left.t2 15.0005
R42 drain_left.n1 drain_left.t0 15.0005
C0 plus drain_right 0.262487f
C1 plus source 0.452448f
C2 plus minus 2.66614f
C3 drain_left drain_right 0.481825f
C4 drain_left source 2.74183f
C5 drain_left minus 0.176915f
C6 source drain_right 2.7405f
C7 minus drain_right 0.477842f
C8 source minus 0.438485f
C9 plus drain_left 0.580155f
C10 drain_right a_n1106_n1292# 3.49622f
C11 drain_left a_n1106_n1292# 3.62299f
C12 source a_n1106_n1292# 2.823476f
C13 minus a_n1106_n1292# 3.253825f
C14 plus a_n1106_n1292# 5.29165f
C15 drain_left.t3 a_n1106_n1292# 0.05152f
C16 drain_left.t1 a_n1106_n1292# 0.05152f
C17 drain_left.n0 a_n1106_n1292# 0.341347f
C18 drain_left.t2 a_n1106_n1292# 0.05152f
C19 drain_left.t0 a_n1106_n1292# 0.05152f
C20 drain_left.n1 a_n1106_n1292# 0.273663f
C21 plus.t1 a_n1106_n1292# 0.04447f
C22 plus.t3 a_n1106_n1292# 0.04447f
C23 plus.n0 a_n1106_n1292# 0.102397f
C24 plus.t0 a_n1106_n1292# 0.04447f
C25 plus.t2 a_n1106_n1292# 0.04447f
C26 plus.n1 a_n1106_n1292# 0.200891f
C27 drain_right.t1 a_n1106_n1292# 0.053178f
C28 drain_right.t2 a_n1106_n1292# 0.053178f
C29 drain_right.n0 a_n1106_n1292# 0.342853f
C30 drain_right.t0 a_n1106_n1292# 0.053178f
C31 drain_right.t3 a_n1106_n1292# 0.053178f
C32 drain_right.n1 a_n1106_n1292# 0.282468f
C33 source.t0 a_n1106_n1292# 0.23569f
C34 source.n0 a_n1106_n1292# 0.449956f
C35 source.t2 a_n1106_n1292# 0.23569f
C36 source.n1 a_n1106_n1292# 0.241992f
C37 source.t4 a_n1106_n1292# 0.23569f
C38 source.n2 a_n1106_n1292# 0.241992f
C39 source.t5 a_n1106_n1292# 0.23569f
C40 source.n3 a_n1106_n1292# 0.625406f
C41 source.t1 a_n1106_n1292# 0.235689f
C42 source.n4 a_n1106_n1292# 0.625407f
C43 source.t3 a_n1106_n1292# 0.235689f
C44 source.n5 a_n1106_n1292# 0.241993f
C45 source.t6 a_n1106_n1292# 0.235689f
C46 source.n6 a_n1106_n1292# 0.241993f
C47 source.t7 a_n1106_n1292# 0.235689f
C48 source.n7 a_n1106_n1292# 0.348646f
C49 source.n8 a_n1106_n1292# 0.465544f
C50 minus.t3 a_n1106_n1292# 0.042956f
C51 minus.t0 a_n1106_n1292# 0.042956f
C52 minus.n0 a_n1106_n1292# 0.207958f
C53 minus.t2 a_n1106_n1292# 0.042956f
C54 minus.t1 a_n1106_n1292# 0.042956f
C55 minus.n1 a_n1106_n1292# 0.094293f
C56 minus.n2 a_n1106_n1292# 2.19607f
.ends

