* NGSPICE file created from diffpair460.ext - technology: sky130A

.subckt diffpair460 minus drain_right drain_left source plus
X0 drain_right minus source a_n1128_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.7
X1 a_n1128_n3292# a_n1128_n3292# a_n1128_n3292# a_n1128_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.7
X2 a_n1128_n3292# a_n1128_n3292# a_n1128_n3292# a_n1128_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X3 drain_left plus source a_n1128_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.7
X4 drain_right minus source a_n1128_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.7
X5 drain_left plus source a_n1128_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.7
X6 a_n1128_n3292# a_n1128_n3292# a_n1128_n3292# a_n1128_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
X7 a_n1128_n3292# a_n1128_n3292# a_n1128_n3292# a_n1128_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.7
.ends

