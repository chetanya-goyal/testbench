* NGSPICE file created from diffpair245.ext - technology: sky130A

.subckt diffpair245 minus drain_right drain_left source plus
X0 source.t21 plus.t0 drain_left.t1 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X1 source.t5 minus.t0 drain_right.t11 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X2 drain_left.t8 plus.t1 source.t20 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X3 drain_left.t7 plus.t2 source.t19 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X4 drain_right.t10 minus.t1 source.t2 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X5 a_n1626_n2088# a_n1626_n2088# a_n1626_n2088# a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=22.8 ps=103.6 w=6 l=0.15
X6 drain_right.t9 minus.t2 source.t9 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X7 a_n1626_n2088# a_n1626_n2088# a_n1626_n2088# a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X8 source.t18 plus.t3 drain_left.t6 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X9 a_n1626_n2088# a_n1626_n2088# a_n1626_n2088# a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X10 source.t8 minus.t3 drain_right.t8 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X11 source.t3 minus.t4 drain_right.t7 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X12 drain_right.t6 minus.t5 source.t4 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X13 drain_right.t5 minus.t6 source.t6 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X14 drain_right.t4 minus.t7 source.t0 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X15 source.t1 minus.t8 drain_right.t3 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X16 a_n1626_n2088# a_n1626_n2088# a_n1626_n2088# a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X17 source.t17 plus.t4 drain_left.t3 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X18 drain_right.t2 minus.t9 source.t7 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X19 source.t22 minus.t10 drain_right.t1 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X20 source.t16 plus.t5 drain_left.t2 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X21 drain_left.t0 plus.t6 source.t15 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X22 source.t23 minus.t11 drain_right.t0 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X23 source.t14 plus.t7 drain_left.t5 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X24 drain_left.t11 plus.t8 source.t13 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X25 drain_left.t10 plus.t9 source.t12 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X26 drain_left.t9 plus.t10 source.t11 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X27 source.t10 plus.t11 drain_left.t4 a_n1626_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
R0 plus.n2 plus.t4 1227.64
R1 plus.n13 plus.t9 1227.64
R2 plus.n17 plus.t1 1227.64
R3 plus.n28 plus.t5 1227.64
R4 plus.n3 plus.t10 1172.87
R5 plus.n4 plus.t7 1172.87
R6 plus.n10 plus.t6 1172.87
R7 plus.n12 plus.t11 1172.87
R8 plus.n19 plus.t3 1172.87
R9 plus.n18 plus.t8 1172.87
R10 plus.n25 plus.t0 1172.87
R11 plus.n27 plus.t2 1172.87
R12 plus.n6 plus.n2 161.489
R13 plus.n21 plus.n17 161.489
R14 plus.n6 plus.n5 161.3
R15 plus.n7 plus.n1 161.3
R16 plus.n9 plus.n8 161.3
R17 plus.n11 plus.n0 161.3
R18 plus.n14 plus.n13 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n22 plus.n16 161.3
R21 plus.n24 plus.n23 161.3
R22 plus.n26 plus.n15 161.3
R23 plus.n29 plus.n28 161.3
R24 plus.n9 plus.n1 73.0308
R25 plus.n24 plus.n16 73.0308
R26 plus.n5 plus.n4 62.0763
R27 plus.n11 plus.n10 62.0763
R28 plus.n26 plus.n25 62.0763
R29 plus.n20 plus.n18 62.0763
R30 plus.n3 plus.n2 40.1672
R31 plus.n13 plus.n12 40.1672
R32 plus.n28 plus.n27 40.1672
R33 plus.n19 plus.n17 40.1672
R34 plus.n5 plus.n3 32.8641
R35 plus.n12 plus.n11 32.8641
R36 plus.n27 plus.n26 32.8641
R37 plus.n20 plus.n19 32.8641
R38 plus plus.n29 26.9308
R39 plus.n4 plus.n1 10.955
R40 plus.n10 plus.n9 10.955
R41 plus.n25 plus.n24 10.955
R42 plus.n18 plus.n16 10.955
R43 plus plus.n14 9.91338
R44 plus.n7 plus.n6 0.189894
R45 plus.n8 plus.n7 0.189894
R46 plus.n8 plus.n0 0.189894
R47 plus.n14 plus.n0 0.189894
R48 plus.n29 plus.n15 0.189894
R49 plus.n23 plus.n15 0.189894
R50 plus.n23 plus.n22 0.189894
R51 plus.n22 plus.n21 0.189894
R52 drain_left.n6 drain_left.n4 67.7512
R53 drain_left.n3 drain_left.n2 67.6957
R54 drain_left.n3 drain_left.n0 67.6957
R55 drain_left.n6 drain_left.n5 67.1908
R56 drain_left.n8 drain_left.n7 67.1907
R57 drain_left.n3 drain_left.n1 67.1907
R58 drain_left drain_left.n3 25.6233
R59 drain_left drain_left.n8 6.21356
R60 drain_left.n1 drain_left.t1 5.0005
R61 drain_left.n1 drain_left.t11 5.0005
R62 drain_left.n2 drain_left.t6 5.0005
R63 drain_left.n2 drain_left.t8 5.0005
R64 drain_left.n0 drain_left.t2 5.0005
R65 drain_left.n0 drain_left.t7 5.0005
R66 drain_left.n7 drain_left.t4 5.0005
R67 drain_left.n7 drain_left.t10 5.0005
R68 drain_left.n5 drain_left.t5 5.0005
R69 drain_left.n5 drain_left.t0 5.0005
R70 drain_left.n4 drain_left.t3 5.0005
R71 drain_left.n4 drain_left.t9 5.0005
R72 drain_left.n8 drain_left.n6 0.560845
R73 source.n5 source.t17 55.512
R74 source.n6 source.t4 55.512
R75 source.n11 source.t23 55.512
R76 source.n0 source.t12 55.5119
R77 source.n23 source.t9 55.5119
R78 source.n18 source.t22 55.5119
R79 source.n17 source.t20 55.5119
R80 source.n12 source.t16 55.5119
R81 source.n2 source.n1 50.512
R82 source.n4 source.n3 50.512
R83 source.n8 source.n7 50.512
R84 source.n10 source.n9 50.512
R85 source.n22 source.n21 50.5119
R86 source.n20 source.n19 50.5119
R87 source.n16 source.n15 50.5119
R88 source.n14 source.n13 50.5119
R89 source.n12 source.n11 17.3026
R90 source.n24 source.n0 11.7595
R91 source.n24 source.n23 5.5436
R92 source.n21 source.t0 5.0005
R93 source.n21 source.t5 5.0005
R94 source.n19 source.t2 5.0005
R95 source.n19 source.t8 5.0005
R96 source.n15 source.t13 5.0005
R97 source.n15 source.t18 5.0005
R98 source.n13 source.t19 5.0005
R99 source.n13 source.t21 5.0005
R100 source.n1 source.t15 5.0005
R101 source.n1 source.t10 5.0005
R102 source.n3 source.t11 5.0005
R103 source.n3 source.t14 5.0005
R104 source.n7 source.t7 5.0005
R105 source.n7 source.t3 5.0005
R106 source.n9 source.t6 5.0005
R107 source.n9 source.t1 5.0005
R108 source.n11 source.n10 0.560845
R109 source.n10 source.n8 0.560845
R110 source.n8 source.n6 0.560845
R111 source.n5 source.n4 0.560845
R112 source.n4 source.n2 0.560845
R113 source.n2 source.n0 0.560845
R114 source.n14 source.n12 0.560845
R115 source.n16 source.n14 0.560845
R116 source.n17 source.n16 0.560845
R117 source.n20 source.n18 0.560845
R118 source.n22 source.n20 0.560845
R119 source.n23 source.n22 0.560845
R120 source.n6 source.n5 0.470328
R121 source.n18 source.n17 0.470328
R122 source source.n24 0.188
R123 minus.n13 minus.t11 1227.64
R124 minus.n2 minus.t5 1227.64
R125 minus.n28 minus.t2 1227.64
R126 minus.n17 minus.t10 1227.64
R127 minus.n12 minus.t6 1172.87
R128 minus.n10 minus.t8 1172.87
R129 minus.n3 minus.t9 1172.87
R130 minus.n4 minus.t4 1172.87
R131 minus.n27 minus.t0 1172.87
R132 minus.n25 minus.t7 1172.87
R133 minus.n19 minus.t3 1172.87
R134 minus.n18 minus.t1 1172.87
R135 minus.n6 minus.n2 161.489
R136 minus.n21 minus.n17 161.489
R137 minus.n14 minus.n13 161.3
R138 minus.n11 minus.n0 161.3
R139 minus.n9 minus.n8 161.3
R140 minus.n7 minus.n1 161.3
R141 minus.n6 minus.n5 161.3
R142 minus.n29 minus.n28 161.3
R143 minus.n26 minus.n15 161.3
R144 minus.n24 minus.n23 161.3
R145 minus.n22 minus.n16 161.3
R146 minus.n21 minus.n20 161.3
R147 minus.n9 minus.n1 73.0308
R148 minus.n24 minus.n16 73.0308
R149 minus.n11 minus.n10 62.0763
R150 minus.n5 minus.n3 62.0763
R151 minus.n20 minus.n19 62.0763
R152 minus.n26 minus.n25 62.0763
R153 minus.n13 minus.n12 40.1672
R154 minus.n4 minus.n2 40.1672
R155 minus.n18 minus.n17 40.1672
R156 minus.n28 minus.n27 40.1672
R157 minus.n12 minus.n11 32.8641
R158 minus.n5 minus.n4 32.8641
R159 minus.n20 minus.n18 32.8641
R160 minus.n27 minus.n26 32.8641
R161 minus.n30 minus.n14 30.777
R162 minus.n10 minus.n9 10.955
R163 minus.n3 minus.n1 10.955
R164 minus.n19 minus.n16 10.955
R165 minus.n25 minus.n24 10.955
R166 minus.n30 minus.n29 6.54217
R167 minus.n14 minus.n0 0.189894
R168 minus.n8 minus.n0 0.189894
R169 minus.n8 minus.n7 0.189894
R170 minus.n7 minus.n6 0.189894
R171 minus.n22 minus.n21 0.189894
R172 minus.n23 minus.n22 0.189894
R173 minus.n23 minus.n15 0.189894
R174 minus.n29 minus.n15 0.189894
R175 minus minus.n30 0.188
R176 drain_right.n6 drain_right.n4 67.751
R177 drain_right.n3 drain_right.n2 67.6957
R178 drain_right.n3 drain_right.n0 67.6957
R179 drain_right.n6 drain_right.n5 67.1908
R180 drain_right.n8 drain_right.n7 67.1908
R181 drain_right.n3 drain_right.n1 67.1907
R182 drain_right drain_right.n3 25.0701
R183 drain_right drain_right.n8 6.21356
R184 drain_right.n1 drain_right.t8 5.0005
R185 drain_right.n1 drain_right.t4 5.0005
R186 drain_right.n2 drain_right.t11 5.0005
R187 drain_right.n2 drain_right.t9 5.0005
R188 drain_right.n0 drain_right.t1 5.0005
R189 drain_right.n0 drain_right.t10 5.0005
R190 drain_right.n4 drain_right.t7 5.0005
R191 drain_right.n4 drain_right.t6 5.0005
R192 drain_right.n5 drain_right.t3 5.0005
R193 drain_right.n5 drain_right.t2 5.0005
R194 drain_right.n7 drain_right.t0 5.0005
R195 drain_right.n7 drain_right.t5 5.0005
R196 drain_right.n8 drain_right.n6 0.560845
C0 plus drain_right 0.309819f
C1 source drain_left 13.1928f
C2 minus plus 4.05263f
C3 source drain_right 13.1927f
C4 source minus 1.46066f
C5 source plus 1.47468f
C6 drain_right drain_left 0.801529f
C7 minus drain_left 0.170585f
C8 plus drain_left 1.80987f
C9 minus drain_right 1.65338f
C10 drain_right a_n1626_n2088# 4.2953f
C11 drain_left a_n1626_n2088# 4.52048f
C12 source a_n1626_n2088# 5.302059f
C13 minus a_n1626_n2088# 5.496103f
C14 plus a_n1626_n2088# 6.37748f
C15 drain_right.t1 a_n1626_n2088# 0.178268f
C16 drain_right.t10 a_n1626_n2088# 0.178268f
C17 drain_right.n0 a_n1626_n2088# 1.1047f
C18 drain_right.t8 a_n1626_n2088# 0.178268f
C19 drain_right.t4 a_n1626_n2088# 0.178268f
C20 drain_right.n1 a_n1626_n2088# 1.10248f
C21 drain_right.t11 a_n1626_n2088# 0.178268f
C22 drain_right.t9 a_n1626_n2088# 0.178268f
C23 drain_right.n2 a_n1626_n2088# 1.1047f
C24 drain_right.n3 a_n1626_n2088# 1.62696f
C25 drain_right.t7 a_n1626_n2088# 0.178268f
C26 drain_right.t6 a_n1626_n2088# 0.178268f
C27 drain_right.n4 a_n1626_n2088# 1.10497f
C28 drain_right.t3 a_n1626_n2088# 0.178268f
C29 drain_right.t2 a_n1626_n2088# 0.178268f
C30 drain_right.n5 a_n1626_n2088# 1.10249f
C31 drain_right.n6 a_n1626_n2088# 0.589532f
C32 drain_right.t0 a_n1626_n2088# 0.178268f
C33 drain_right.t5 a_n1626_n2088# 0.178268f
C34 drain_right.n7 a_n1626_n2088# 1.10249f
C35 drain_right.n8 a_n1626_n2088# 0.498241f
C36 minus.n0 a_n1626_n2088# 0.031496f
C37 minus.t11 a_n1626_n2088# 0.082657f
C38 minus.t6 a_n1626_n2088# 0.080765f
C39 minus.t8 a_n1626_n2088# 0.080765f
C40 minus.n1 a_n1626_n2088# 0.011905f
C41 minus.t5 a_n1626_n2088# 0.082657f
C42 minus.n2 a_n1626_n2088# 0.053927f
C43 minus.t9 a_n1626_n2088# 0.080765f
C44 minus.n3 a_n1626_n2088# 0.041927f
C45 minus.t4 a_n1626_n2088# 0.080765f
C46 minus.n4 a_n1626_n2088# 0.041927f
C47 minus.n5 a_n1626_n2088# 0.013361f
C48 minus.n6 a_n1626_n2088# 0.070714f
C49 minus.n7 a_n1626_n2088# 0.031496f
C50 minus.n8 a_n1626_n2088# 0.031496f
C51 minus.n9 a_n1626_n2088# 0.011905f
C52 minus.n10 a_n1626_n2088# 0.041927f
C53 minus.n11 a_n1626_n2088# 0.013361f
C54 minus.n12 a_n1626_n2088# 0.041927f
C55 minus.n13 a_n1626_n2088# 0.053881f
C56 minus.n14 a_n1626_n2088# 0.856883f
C57 minus.n15 a_n1626_n2088# 0.031496f
C58 minus.t0 a_n1626_n2088# 0.080765f
C59 minus.t7 a_n1626_n2088# 0.080765f
C60 minus.n16 a_n1626_n2088# 0.011905f
C61 minus.t10 a_n1626_n2088# 0.082657f
C62 minus.n17 a_n1626_n2088# 0.053927f
C63 minus.t1 a_n1626_n2088# 0.080765f
C64 minus.n18 a_n1626_n2088# 0.041927f
C65 minus.t3 a_n1626_n2088# 0.080765f
C66 minus.n19 a_n1626_n2088# 0.041927f
C67 minus.n20 a_n1626_n2088# 0.013361f
C68 minus.n21 a_n1626_n2088# 0.070714f
C69 minus.n22 a_n1626_n2088# 0.031496f
C70 minus.n23 a_n1626_n2088# 0.031496f
C71 minus.n24 a_n1626_n2088# 0.011905f
C72 minus.n25 a_n1626_n2088# 0.041927f
C73 minus.n26 a_n1626_n2088# 0.013361f
C74 minus.n27 a_n1626_n2088# 0.041927f
C75 minus.t2 a_n1626_n2088# 0.082657f
C76 minus.n28 a_n1626_n2088# 0.053881f
C77 minus.n29 a_n1626_n2088# 0.209037f
C78 minus.n30 a_n1626_n2088# 1.05415f
C79 source.t12 a_n1626_n2088# 1.08537f
C80 source.n0 a_n1626_n2088# 0.798479f
C81 source.t15 a_n1626_n2088# 0.154527f
C82 source.t10 a_n1626_n2088# 0.154527f
C83 source.n1 a_n1626_n2088# 0.899366f
C84 source.n2 a_n1626_n2088# 0.279312f
C85 source.t11 a_n1626_n2088# 0.154527f
C86 source.t14 a_n1626_n2088# 0.154527f
C87 source.n3 a_n1626_n2088# 0.899366f
C88 source.n4 a_n1626_n2088# 0.279312f
C89 source.t17 a_n1626_n2088# 1.08537f
C90 source.n5 a_n1626_n2088# 0.36518f
C91 source.t4 a_n1626_n2088# 1.08537f
C92 source.n6 a_n1626_n2088# 0.36518f
C93 source.t7 a_n1626_n2088# 0.154527f
C94 source.t3 a_n1626_n2088# 0.154527f
C95 source.n7 a_n1626_n2088# 0.899366f
C96 source.n8 a_n1626_n2088# 0.279312f
C97 source.t6 a_n1626_n2088# 0.154527f
C98 source.t1 a_n1626_n2088# 0.154527f
C99 source.n9 a_n1626_n2088# 0.899366f
C100 source.n10 a_n1626_n2088# 0.279312f
C101 source.t23 a_n1626_n2088# 1.08537f
C102 source.n11 a_n1626_n2088# 1.07573f
C103 source.t16 a_n1626_n2088# 1.08537f
C104 source.n12 a_n1626_n2088# 1.07574f
C105 source.t19 a_n1626_n2088# 0.154527f
C106 source.t21 a_n1626_n2088# 0.154527f
C107 source.n13 a_n1626_n2088# 0.899361f
C108 source.n14 a_n1626_n2088# 0.279317f
C109 source.t13 a_n1626_n2088# 0.154527f
C110 source.t18 a_n1626_n2088# 0.154527f
C111 source.n15 a_n1626_n2088# 0.899361f
C112 source.n16 a_n1626_n2088# 0.279317f
C113 source.t20 a_n1626_n2088# 1.08537f
C114 source.n17 a_n1626_n2088# 0.365185f
C115 source.t22 a_n1626_n2088# 1.08537f
C116 source.n18 a_n1626_n2088# 0.365185f
C117 source.t2 a_n1626_n2088# 0.154527f
C118 source.t8 a_n1626_n2088# 0.154527f
C119 source.n19 a_n1626_n2088# 0.899361f
C120 source.n20 a_n1626_n2088# 0.279317f
C121 source.t0 a_n1626_n2088# 0.154527f
C122 source.t5 a_n1626_n2088# 0.154527f
C123 source.n21 a_n1626_n2088# 0.899361f
C124 source.n22 a_n1626_n2088# 0.279317f
C125 source.t9 a_n1626_n2088# 1.08537f
C126 source.n23 a_n1626_n2088# 0.487564f
C127 source.n24 a_n1626_n2088# 0.880737f
C128 drain_left.t2 a_n1626_n2088# 0.176966f
C129 drain_left.t7 a_n1626_n2088# 0.176966f
C130 drain_left.n0 a_n1626_n2088# 1.09664f
C131 drain_left.t1 a_n1626_n2088# 0.176966f
C132 drain_left.t11 a_n1626_n2088# 0.176966f
C133 drain_left.n1 a_n1626_n2088# 1.09443f
C134 drain_left.t6 a_n1626_n2088# 0.176966f
C135 drain_left.t8 a_n1626_n2088# 0.176966f
C136 drain_left.n2 a_n1626_n2088# 1.09664f
C137 drain_left.n3 a_n1626_n2088# 1.66527f
C138 drain_left.t3 a_n1626_n2088# 0.176966f
C139 drain_left.t9 a_n1626_n2088# 0.176966f
C140 drain_left.n4 a_n1626_n2088# 1.09691f
C141 drain_left.t5 a_n1626_n2088# 0.176966f
C142 drain_left.t0 a_n1626_n2088# 0.176966f
C143 drain_left.n5 a_n1626_n2088# 1.09444f
C144 drain_left.n6 a_n1626_n2088# 0.585224f
C145 drain_left.t4 a_n1626_n2088# 0.176966f
C146 drain_left.t10 a_n1626_n2088# 0.176966f
C147 drain_left.n7 a_n1626_n2088# 1.09443f
C148 drain_left.n8 a_n1626_n2088# 0.494609f
C149 plus.n0 a_n1626_n2088# 0.031993f
C150 plus.t11 a_n1626_n2088# 0.082039f
C151 plus.t6 a_n1626_n2088# 0.082039f
C152 plus.n1 a_n1626_n2088# 0.012093f
C153 plus.t4 a_n1626_n2088# 0.083961f
C154 plus.n2 a_n1626_n2088# 0.054778f
C155 plus.t10 a_n1626_n2088# 0.082039f
C156 plus.n3 a_n1626_n2088# 0.042589f
C157 plus.t7 a_n1626_n2088# 0.082039f
C158 plus.n4 a_n1626_n2088# 0.042589f
C159 plus.n5 a_n1626_n2088# 0.013572f
C160 plus.n6 a_n1626_n2088# 0.07183f
C161 plus.n7 a_n1626_n2088# 0.031993f
C162 plus.n8 a_n1626_n2088# 0.031993f
C163 plus.n9 a_n1626_n2088# 0.012093f
C164 plus.n10 a_n1626_n2088# 0.042589f
C165 plus.n11 a_n1626_n2088# 0.013572f
C166 plus.n12 a_n1626_n2088# 0.042589f
C167 plus.t9 a_n1626_n2088# 0.083961f
C168 plus.n13 a_n1626_n2088# 0.054731f
C169 plus.n14 a_n1626_n2088# 0.277459f
C170 plus.n15 a_n1626_n2088# 0.031993f
C171 plus.t5 a_n1626_n2088# 0.083961f
C172 plus.t2 a_n1626_n2088# 0.082039f
C173 plus.t0 a_n1626_n2088# 0.082039f
C174 plus.n16 a_n1626_n2088# 0.012093f
C175 plus.t1 a_n1626_n2088# 0.083961f
C176 plus.n17 a_n1626_n2088# 0.054778f
C177 plus.t8 a_n1626_n2088# 0.082039f
C178 plus.n18 a_n1626_n2088# 0.042589f
C179 plus.t3 a_n1626_n2088# 0.082039f
C180 plus.n19 a_n1626_n2088# 0.042589f
C181 plus.n20 a_n1626_n2088# 0.013572f
C182 plus.n21 a_n1626_n2088# 0.07183f
C183 plus.n22 a_n1626_n2088# 0.031993f
C184 plus.n23 a_n1626_n2088# 0.031993f
C185 plus.n24 a_n1626_n2088# 0.012093f
C186 plus.n25 a_n1626_n2088# 0.042589f
C187 plus.n26 a_n1626_n2088# 0.013572f
C188 plus.n27 a_n1626_n2088# 0.042589f
C189 plus.n28 a_n1626_n2088# 0.054731f
C190 plus.n29 a_n1626_n2088# 0.786713f
.ends

