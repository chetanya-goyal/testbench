* NGSPICE file created from diffpair295.ext - technology: sky130A

.subckt diffpair295 minus drain_right drain_left source plus
X0 source.t18 plus.t0 drain_left.t0 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X1 a_n2018_n2088# a_n2018_n2088# a_n2018_n2088# a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.6
X2 drain_left.t1 plus.t1 source.t17 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X3 drain_right.t11 minus.t0 source.t0 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X4 source.t2 minus.t1 drain_right.t10 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X5 a_n2018_n2088# a_n2018_n2088# a_n2018_n2088# a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.6
X6 source.t20 minus.t2 drain_right.t9 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X7 drain_left.t2 plus.t2 source.t16 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X8 source.t15 plus.t3 drain_left.t3 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X9 source.t21 minus.t3 drain_right.t8 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X10 drain_right.t7 minus.t4 source.t22 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X11 drain_left.t4 plus.t4 source.t14 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X12 drain_right.t6 minus.t5 source.t23 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X13 source.t13 plus.t5 drain_left.t5 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X14 drain_left.t6 plus.t6 source.t12 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X15 source.t4 minus.t6 drain_right.t5 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X16 source.t11 plus.t7 drain_left.t7 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X17 drain_right.t4 minus.t7 source.t3 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X18 drain_right.t3 minus.t8 source.t6 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.6
X19 a_n2018_n2088# a_n2018_n2088# a_n2018_n2088# a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.6
X20 drain_left.t8 plus.t8 source.t10 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X21 source.t9 plus.t9 drain_left.t9 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X22 drain_left.t10 plus.t10 source.t8 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X23 source.t5 minus.t9 drain_right.t2 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X24 drain_right.t1 minus.t10 source.t19 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
X25 a_n2018_n2088# a_n2018_n2088# a_n2018_n2088# a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.6
X26 source.t7 plus.t11 drain_left.t11 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.6
X27 source.t1 minus.t11 drain_right.t0 a_n2018_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.6
R0 plus.n4 plus.t9 331.531
R1 plus.n16 plus.t4 331.531
R2 plus.n10 plus.t1 306.473
R3 plus.n8 plus.t3 306.473
R4 plus.n7 plus.t6 306.473
R5 plus.n6 plus.t7 306.473
R6 plus.n5 plus.t8 306.473
R7 plus.n22 plus.t11 306.473
R8 plus.n20 plus.t10 306.473
R9 plus.n19 plus.t5 306.473
R10 plus.n18 plus.t2 306.473
R11 plus.n17 plus.t0 306.473
R12 plus.n8 plus.n1 161.3
R13 plus.n9 plus.n0 161.3
R14 plus.n11 plus.n10 161.3
R15 plus.n20 plus.n13 161.3
R16 plus.n21 plus.n12 161.3
R17 plus.n23 plus.n22 161.3
R18 plus.n6 plus.n3 80.6037
R19 plus.n7 plus.n2 80.6037
R20 plus.n18 plus.n15 80.6037
R21 plus.n19 plus.n14 80.6037
R22 plus.n8 plus.n7 48.2005
R23 plus.n7 plus.n6 48.2005
R24 plus.n6 plus.n5 48.2005
R25 plus.n20 plus.n19 48.2005
R26 plus.n19 plus.n18 48.2005
R27 plus.n18 plus.n17 48.2005
R28 plus.n4 plus.n3 45.0744
R29 plus.n16 plus.n15 45.0744
R30 plus.n10 plus.n9 40.1672
R31 plus.n22 plus.n21 40.1672
R32 plus plus.n23 28.4611
R33 plus.n5 plus.n4 16.1124
R34 plus.n17 plus.n16 16.1124
R35 plus plus.n11 9.95883
R36 plus.n9 plus.n8 8.03383
R37 plus.n21 plus.n20 8.03383
R38 plus.n3 plus.n2 0.380177
R39 plus.n15 plus.n14 0.380177
R40 plus.n2 plus.n1 0.285035
R41 plus.n14 plus.n13 0.285035
R42 plus.n1 plus.n0 0.189894
R43 plus.n11 plus.n0 0.189894
R44 plus.n23 plus.n12 0.189894
R45 plus.n13 plus.n12 0.189894
R46 drain_left.n6 drain_left.n4 67.9925
R47 drain_left.n3 drain_left.n2 67.937
R48 drain_left.n3 drain_left.n0 67.937
R49 drain_left.n6 drain_left.n5 67.1908
R50 drain_left.n8 drain_left.n7 67.1907
R51 drain_left.n3 drain_left.n1 67.1907
R52 drain_left drain_left.n3 26.8302
R53 drain_left drain_left.n8 6.45494
R54 drain_left.n1 drain_left.t5 3.3005
R55 drain_left.n1 drain_left.t2 3.3005
R56 drain_left.n2 drain_left.t0 3.3005
R57 drain_left.n2 drain_left.t4 3.3005
R58 drain_left.n0 drain_left.t11 3.3005
R59 drain_left.n0 drain_left.t10 3.3005
R60 drain_left.n7 drain_left.t3 3.3005
R61 drain_left.n7 drain_left.t1 3.3005
R62 drain_left.n5 drain_left.t7 3.3005
R63 drain_left.n5 drain_left.t6 3.3005
R64 drain_left.n4 drain_left.t9 3.3005
R65 drain_left.n4 drain_left.t8 3.3005
R66 drain_left.n8 drain_left.n6 0.802224
R67 source.n266 source.n240 289.615
R68 source.n230 source.n204 289.615
R69 source.n198 source.n172 289.615
R70 source.n162 source.n136 289.615
R71 source.n26 source.n0 289.615
R72 source.n62 source.n36 289.615
R73 source.n94 source.n68 289.615
R74 source.n130 source.n104 289.615
R75 source.n251 source.n250 185
R76 source.n248 source.n247 185
R77 source.n257 source.n256 185
R78 source.n259 source.n258 185
R79 source.n244 source.n243 185
R80 source.n265 source.n264 185
R81 source.n267 source.n266 185
R82 source.n215 source.n214 185
R83 source.n212 source.n211 185
R84 source.n221 source.n220 185
R85 source.n223 source.n222 185
R86 source.n208 source.n207 185
R87 source.n229 source.n228 185
R88 source.n231 source.n230 185
R89 source.n183 source.n182 185
R90 source.n180 source.n179 185
R91 source.n189 source.n188 185
R92 source.n191 source.n190 185
R93 source.n176 source.n175 185
R94 source.n197 source.n196 185
R95 source.n199 source.n198 185
R96 source.n147 source.n146 185
R97 source.n144 source.n143 185
R98 source.n153 source.n152 185
R99 source.n155 source.n154 185
R100 source.n140 source.n139 185
R101 source.n161 source.n160 185
R102 source.n163 source.n162 185
R103 source.n27 source.n26 185
R104 source.n25 source.n24 185
R105 source.n4 source.n3 185
R106 source.n19 source.n18 185
R107 source.n17 source.n16 185
R108 source.n8 source.n7 185
R109 source.n11 source.n10 185
R110 source.n63 source.n62 185
R111 source.n61 source.n60 185
R112 source.n40 source.n39 185
R113 source.n55 source.n54 185
R114 source.n53 source.n52 185
R115 source.n44 source.n43 185
R116 source.n47 source.n46 185
R117 source.n95 source.n94 185
R118 source.n93 source.n92 185
R119 source.n72 source.n71 185
R120 source.n87 source.n86 185
R121 source.n85 source.n84 185
R122 source.n76 source.n75 185
R123 source.n79 source.n78 185
R124 source.n131 source.n130 185
R125 source.n129 source.n128 185
R126 source.n108 source.n107 185
R127 source.n123 source.n122 185
R128 source.n121 source.n120 185
R129 source.n112 source.n111 185
R130 source.n115 source.n114 185
R131 source.t6 source.n249 147.661
R132 source.t2 source.n213 147.661
R133 source.t14 source.n181 147.661
R134 source.t7 source.n145 147.661
R135 source.t17 source.n9 147.661
R136 source.t9 source.n45 147.661
R137 source.t3 source.n77 147.661
R138 source.t20 source.n113 147.661
R139 source.n250 source.n247 104.615
R140 source.n257 source.n247 104.615
R141 source.n258 source.n257 104.615
R142 source.n258 source.n243 104.615
R143 source.n265 source.n243 104.615
R144 source.n266 source.n265 104.615
R145 source.n214 source.n211 104.615
R146 source.n221 source.n211 104.615
R147 source.n222 source.n221 104.615
R148 source.n222 source.n207 104.615
R149 source.n229 source.n207 104.615
R150 source.n230 source.n229 104.615
R151 source.n182 source.n179 104.615
R152 source.n189 source.n179 104.615
R153 source.n190 source.n189 104.615
R154 source.n190 source.n175 104.615
R155 source.n197 source.n175 104.615
R156 source.n198 source.n197 104.615
R157 source.n146 source.n143 104.615
R158 source.n153 source.n143 104.615
R159 source.n154 source.n153 104.615
R160 source.n154 source.n139 104.615
R161 source.n161 source.n139 104.615
R162 source.n162 source.n161 104.615
R163 source.n26 source.n25 104.615
R164 source.n25 source.n3 104.615
R165 source.n18 source.n3 104.615
R166 source.n18 source.n17 104.615
R167 source.n17 source.n7 104.615
R168 source.n10 source.n7 104.615
R169 source.n62 source.n61 104.615
R170 source.n61 source.n39 104.615
R171 source.n54 source.n39 104.615
R172 source.n54 source.n53 104.615
R173 source.n53 source.n43 104.615
R174 source.n46 source.n43 104.615
R175 source.n94 source.n93 104.615
R176 source.n93 source.n71 104.615
R177 source.n86 source.n71 104.615
R178 source.n86 source.n85 104.615
R179 source.n85 source.n75 104.615
R180 source.n78 source.n75 104.615
R181 source.n130 source.n129 104.615
R182 source.n129 source.n107 104.615
R183 source.n122 source.n107 104.615
R184 source.n122 source.n121 104.615
R185 source.n121 source.n111 104.615
R186 source.n114 source.n111 104.615
R187 source.n250 source.t6 52.3082
R188 source.n214 source.t2 52.3082
R189 source.n182 source.t14 52.3082
R190 source.n146 source.t7 52.3082
R191 source.n10 source.t17 52.3082
R192 source.n46 source.t9 52.3082
R193 source.n78 source.t3 52.3082
R194 source.n114 source.t20 52.3082
R195 source.n33 source.n32 50.512
R196 source.n35 source.n34 50.512
R197 source.n101 source.n100 50.512
R198 source.n103 source.n102 50.512
R199 source.n239 source.n238 50.5119
R200 source.n237 source.n236 50.5119
R201 source.n171 source.n170 50.5119
R202 source.n169 source.n168 50.5119
R203 source.n271 source.n270 32.1853
R204 source.n235 source.n234 32.1853
R205 source.n203 source.n202 32.1853
R206 source.n167 source.n166 32.1853
R207 source.n31 source.n30 32.1853
R208 source.n67 source.n66 32.1853
R209 source.n99 source.n98 32.1853
R210 source.n135 source.n134 32.1853
R211 source.n167 source.n135 17.544
R212 source.n251 source.n249 15.6674
R213 source.n215 source.n213 15.6674
R214 source.n183 source.n181 15.6674
R215 source.n147 source.n145 15.6674
R216 source.n11 source.n9 15.6674
R217 source.n47 source.n45 15.6674
R218 source.n79 source.n77 15.6674
R219 source.n115 source.n113 15.6674
R220 source.n252 source.n248 12.8005
R221 source.n216 source.n212 12.8005
R222 source.n184 source.n180 12.8005
R223 source.n148 source.n144 12.8005
R224 source.n12 source.n8 12.8005
R225 source.n48 source.n44 12.8005
R226 source.n80 source.n76 12.8005
R227 source.n116 source.n112 12.8005
R228 source.n256 source.n255 12.0247
R229 source.n220 source.n219 12.0247
R230 source.n188 source.n187 12.0247
R231 source.n152 source.n151 12.0247
R232 source.n16 source.n15 12.0247
R233 source.n52 source.n51 12.0247
R234 source.n84 source.n83 12.0247
R235 source.n120 source.n119 12.0247
R236 source.n272 source.n31 11.8802
R237 source.n259 source.n246 11.249
R238 source.n223 source.n210 11.249
R239 source.n191 source.n178 11.249
R240 source.n155 source.n142 11.249
R241 source.n19 source.n6 11.249
R242 source.n55 source.n42 11.249
R243 source.n87 source.n74 11.249
R244 source.n123 source.n110 11.249
R245 source.n260 source.n244 10.4732
R246 source.n224 source.n208 10.4732
R247 source.n192 source.n176 10.4732
R248 source.n156 source.n140 10.4732
R249 source.n20 source.n4 10.4732
R250 source.n56 source.n40 10.4732
R251 source.n88 source.n72 10.4732
R252 source.n124 source.n108 10.4732
R253 source.n264 source.n263 9.69747
R254 source.n228 source.n227 9.69747
R255 source.n196 source.n195 9.69747
R256 source.n160 source.n159 9.69747
R257 source.n24 source.n23 9.69747
R258 source.n60 source.n59 9.69747
R259 source.n92 source.n91 9.69747
R260 source.n128 source.n127 9.69747
R261 source.n270 source.n269 9.45567
R262 source.n234 source.n233 9.45567
R263 source.n202 source.n201 9.45567
R264 source.n166 source.n165 9.45567
R265 source.n30 source.n29 9.45567
R266 source.n66 source.n65 9.45567
R267 source.n98 source.n97 9.45567
R268 source.n134 source.n133 9.45567
R269 source.n269 source.n268 9.3005
R270 source.n242 source.n241 9.3005
R271 source.n263 source.n262 9.3005
R272 source.n261 source.n260 9.3005
R273 source.n246 source.n245 9.3005
R274 source.n255 source.n254 9.3005
R275 source.n253 source.n252 9.3005
R276 source.n233 source.n232 9.3005
R277 source.n206 source.n205 9.3005
R278 source.n227 source.n226 9.3005
R279 source.n225 source.n224 9.3005
R280 source.n210 source.n209 9.3005
R281 source.n219 source.n218 9.3005
R282 source.n217 source.n216 9.3005
R283 source.n201 source.n200 9.3005
R284 source.n174 source.n173 9.3005
R285 source.n195 source.n194 9.3005
R286 source.n193 source.n192 9.3005
R287 source.n178 source.n177 9.3005
R288 source.n187 source.n186 9.3005
R289 source.n185 source.n184 9.3005
R290 source.n165 source.n164 9.3005
R291 source.n138 source.n137 9.3005
R292 source.n159 source.n158 9.3005
R293 source.n157 source.n156 9.3005
R294 source.n142 source.n141 9.3005
R295 source.n151 source.n150 9.3005
R296 source.n149 source.n148 9.3005
R297 source.n29 source.n28 9.3005
R298 source.n2 source.n1 9.3005
R299 source.n23 source.n22 9.3005
R300 source.n21 source.n20 9.3005
R301 source.n6 source.n5 9.3005
R302 source.n15 source.n14 9.3005
R303 source.n13 source.n12 9.3005
R304 source.n65 source.n64 9.3005
R305 source.n38 source.n37 9.3005
R306 source.n59 source.n58 9.3005
R307 source.n57 source.n56 9.3005
R308 source.n42 source.n41 9.3005
R309 source.n51 source.n50 9.3005
R310 source.n49 source.n48 9.3005
R311 source.n97 source.n96 9.3005
R312 source.n70 source.n69 9.3005
R313 source.n91 source.n90 9.3005
R314 source.n89 source.n88 9.3005
R315 source.n74 source.n73 9.3005
R316 source.n83 source.n82 9.3005
R317 source.n81 source.n80 9.3005
R318 source.n133 source.n132 9.3005
R319 source.n106 source.n105 9.3005
R320 source.n127 source.n126 9.3005
R321 source.n125 source.n124 9.3005
R322 source.n110 source.n109 9.3005
R323 source.n119 source.n118 9.3005
R324 source.n117 source.n116 9.3005
R325 source.n267 source.n242 8.92171
R326 source.n231 source.n206 8.92171
R327 source.n199 source.n174 8.92171
R328 source.n163 source.n138 8.92171
R329 source.n27 source.n2 8.92171
R330 source.n63 source.n38 8.92171
R331 source.n95 source.n70 8.92171
R332 source.n131 source.n106 8.92171
R333 source.n268 source.n240 8.14595
R334 source.n232 source.n204 8.14595
R335 source.n200 source.n172 8.14595
R336 source.n164 source.n136 8.14595
R337 source.n28 source.n0 8.14595
R338 source.n64 source.n36 8.14595
R339 source.n96 source.n68 8.14595
R340 source.n132 source.n104 8.14595
R341 source.n270 source.n240 5.81868
R342 source.n234 source.n204 5.81868
R343 source.n202 source.n172 5.81868
R344 source.n166 source.n136 5.81868
R345 source.n30 source.n0 5.81868
R346 source.n66 source.n36 5.81868
R347 source.n98 source.n68 5.81868
R348 source.n134 source.n104 5.81868
R349 source.n272 source.n271 5.66429
R350 source.n268 source.n267 5.04292
R351 source.n232 source.n231 5.04292
R352 source.n200 source.n199 5.04292
R353 source.n164 source.n163 5.04292
R354 source.n28 source.n27 5.04292
R355 source.n64 source.n63 5.04292
R356 source.n96 source.n95 5.04292
R357 source.n132 source.n131 5.04292
R358 source.n253 source.n249 4.38594
R359 source.n217 source.n213 4.38594
R360 source.n185 source.n181 4.38594
R361 source.n149 source.n145 4.38594
R362 source.n13 source.n9 4.38594
R363 source.n49 source.n45 4.38594
R364 source.n81 source.n77 4.38594
R365 source.n117 source.n113 4.38594
R366 source.n264 source.n242 4.26717
R367 source.n228 source.n206 4.26717
R368 source.n196 source.n174 4.26717
R369 source.n160 source.n138 4.26717
R370 source.n24 source.n2 4.26717
R371 source.n60 source.n38 4.26717
R372 source.n92 source.n70 4.26717
R373 source.n128 source.n106 4.26717
R374 source.n263 source.n244 3.49141
R375 source.n227 source.n208 3.49141
R376 source.n195 source.n176 3.49141
R377 source.n159 source.n140 3.49141
R378 source.n23 source.n4 3.49141
R379 source.n59 source.n40 3.49141
R380 source.n91 source.n72 3.49141
R381 source.n127 source.n108 3.49141
R382 source.n238 source.t22 3.3005
R383 source.n238 source.t5 3.3005
R384 source.n236 source.t19 3.3005
R385 source.n236 source.t1 3.3005
R386 source.n170 source.t16 3.3005
R387 source.n170 source.t18 3.3005
R388 source.n168 source.t8 3.3005
R389 source.n168 source.t13 3.3005
R390 source.n32 source.t12 3.3005
R391 source.n32 source.t15 3.3005
R392 source.n34 source.t10 3.3005
R393 source.n34 source.t11 3.3005
R394 source.n100 source.t23 3.3005
R395 source.n100 source.t4 3.3005
R396 source.n102 source.t0 3.3005
R397 source.n102 source.t21 3.3005
R398 source.n260 source.n259 2.71565
R399 source.n224 source.n223 2.71565
R400 source.n192 source.n191 2.71565
R401 source.n156 source.n155 2.71565
R402 source.n20 source.n19 2.71565
R403 source.n56 source.n55 2.71565
R404 source.n88 source.n87 2.71565
R405 source.n124 source.n123 2.71565
R406 source.n256 source.n246 1.93989
R407 source.n220 source.n210 1.93989
R408 source.n188 source.n178 1.93989
R409 source.n152 source.n142 1.93989
R410 source.n16 source.n6 1.93989
R411 source.n52 source.n42 1.93989
R412 source.n84 source.n74 1.93989
R413 source.n120 source.n110 1.93989
R414 source.n255 source.n248 1.16414
R415 source.n219 source.n212 1.16414
R416 source.n187 source.n180 1.16414
R417 source.n151 source.n144 1.16414
R418 source.n15 source.n8 1.16414
R419 source.n51 source.n44 1.16414
R420 source.n83 source.n76 1.16414
R421 source.n119 source.n112 1.16414
R422 source.n135 source.n103 0.802224
R423 source.n103 source.n101 0.802224
R424 source.n101 source.n99 0.802224
R425 source.n67 source.n35 0.802224
R426 source.n35 source.n33 0.802224
R427 source.n33 source.n31 0.802224
R428 source.n169 source.n167 0.802224
R429 source.n171 source.n169 0.802224
R430 source.n203 source.n171 0.802224
R431 source.n237 source.n235 0.802224
R432 source.n239 source.n237 0.802224
R433 source.n271 source.n239 0.802224
R434 source.n99 source.n67 0.470328
R435 source.n235 source.n203 0.470328
R436 source.n252 source.n251 0.388379
R437 source.n216 source.n215 0.388379
R438 source.n184 source.n183 0.388379
R439 source.n148 source.n147 0.388379
R440 source.n12 source.n11 0.388379
R441 source.n48 source.n47 0.388379
R442 source.n80 source.n79 0.388379
R443 source.n116 source.n115 0.388379
R444 source source.n272 0.188
R445 source.n254 source.n253 0.155672
R446 source.n254 source.n245 0.155672
R447 source.n261 source.n245 0.155672
R448 source.n262 source.n261 0.155672
R449 source.n262 source.n241 0.155672
R450 source.n269 source.n241 0.155672
R451 source.n218 source.n217 0.155672
R452 source.n218 source.n209 0.155672
R453 source.n225 source.n209 0.155672
R454 source.n226 source.n225 0.155672
R455 source.n226 source.n205 0.155672
R456 source.n233 source.n205 0.155672
R457 source.n186 source.n185 0.155672
R458 source.n186 source.n177 0.155672
R459 source.n193 source.n177 0.155672
R460 source.n194 source.n193 0.155672
R461 source.n194 source.n173 0.155672
R462 source.n201 source.n173 0.155672
R463 source.n150 source.n149 0.155672
R464 source.n150 source.n141 0.155672
R465 source.n157 source.n141 0.155672
R466 source.n158 source.n157 0.155672
R467 source.n158 source.n137 0.155672
R468 source.n165 source.n137 0.155672
R469 source.n29 source.n1 0.155672
R470 source.n22 source.n1 0.155672
R471 source.n22 source.n21 0.155672
R472 source.n21 source.n5 0.155672
R473 source.n14 source.n5 0.155672
R474 source.n14 source.n13 0.155672
R475 source.n65 source.n37 0.155672
R476 source.n58 source.n37 0.155672
R477 source.n58 source.n57 0.155672
R478 source.n57 source.n41 0.155672
R479 source.n50 source.n41 0.155672
R480 source.n50 source.n49 0.155672
R481 source.n97 source.n69 0.155672
R482 source.n90 source.n69 0.155672
R483 source.n90 source.n89 0.155672
R484 source.n89 source.n73 0.155672
R485 source.n82 source.n73 0.155672
R486 source.n82 source.n81 0.155672
R487 source.n133 source.n105 0.155672
R488 source.n126 source.n105 0.155672
R489 source.n126 source.n125 0.155672
R490 source.n125 source.n109 0.155672
R491 source.n118 source.n109 0.155672
R492 source.n118 source.n117 0.155672
R493 minus.n2 minus.t7 331.531
R494 minus.n14 minus.t1 331.531
R495 minus.n3 minus.t6 306.473
R496 minus.n4 minus.t5 306.473
R497 minus.n1 minus.t3 306.473
R498 minus.n8 minus.t0 306.473
R499 minus.n10 minus.t2 306.473
R500 minus.n15 minus.t10 306.473
R501 minus.n16 minus.t11 306.473
R502 minus.n13 minus.t4 306.473
R503 minus.n20 minus.t9 306.473
R504 minus.n22 minus.t8 306.473
R505 minus.n11 minus.n10 161.3
R506 minus.n9 minus.n0 161.3
R507 minus.n8 minus.n7 161.3
R508 minus.n23 minus.n22 161.3
R509 minus.n21 minus.n12 161.3
R510 minus.n20 minus.n19 161.3
R511 minus.n6 minus.n1 80.6037
R512 minus.n5 minus.n4 80.6037
R513 minus.n18 minus.n13 80.6037
R514 minus.n17 minus.n16 80.6037
R515 minus.n4 minus.n3 48.2005
R516 minus.n4 minus.n1 48.2005
R517 minus.n8 minus.n1 48.2005
R518 minus.n16 minus.n15 48.2005
R519 minus.n16 minus.n13 48.2005
R520 minus.n20 minus.n13 48.2005
R521 minus.n5 minus.n2 45.0744
R522 minus.n17 minus.n14 45.0744
R523 minus.n10 minus.n9 40.1672
R524 minus.n22 minus.n21 40.1672
R525 minus.n24 minus.n11 32.3073
R526 minus.n3 minus.n2 16.1124
R527 minus.n15 minus.n14 16.1124
R528 minus.n9 minus.n8 8.03383
R529 minus.n21 minus.n20 8.03383
R530 minus.n24 minus.n23 6.58762
R531 minus.n6 minus.n5 0.380177
R532 minus.n18 minus.n17 0.380177
R533 minus.n7 minus.n6 0.285035
R534 minus.n19 minus.n18 0.285035
R535 minus.n11 minus.n0 0.189894
R536 minus.n7 minus.n0 0.189894
R537 minus.n19 minus.n12 0.189894
R538 minus.n23 minus.n12 0.189894
R539 minus minus.n24 0.188
R540 drain_right.n6 drain_right.n4 67.9924
R541 drain_right.n3 drain_right.n2 67.937
R542 drain_right.n3 drain_right.n0 67.937
R543 drain_right.n6 drain_right.n5 67.1908
R544 drain_right.n8 drain_right.n7 67.1908
R545 drain_right.n3 drain_right.n1 67.1907
R546 drain_right drain_right.n3 26.277
R547 drain_right drain_right.n8 6.45494
R548 drain_right.n1 drain_right.t0 3.3005
R549 drain_right.n1 drain_right.t7 3.3005
R550 drain_right.n2 drain_right.t2 3.3005
R551 drain_right.n2 drain_right.t3 3.3005
R552 drain_right.n0 drain_right.t10 3.3005
R553 drain_right.n0 drain_right.t1 3.3005
R554 drain_right.n4 drain_right.t5 3.3005
R555 drain_right.n4 drain_right.t4 3.3005
R556 drain_right.n5 drain_right.t8 3.3005
R557 drain_right.n5 drain_right.t6 3.3005
R558 drain_right.n7 drain_right.t9 3.3005
R559 drain_right.n7 drain_right.t11 3.3005
R560 drain_right.n8 drain_right.n6 0.802224
C0 source drain_left 9.69561f
C1 drain_right minus 3.8498f
C2 drain_right plus 0.352374f
C3 plus minus 4.55291f
C4 source drain_right 9.697121f
C5 source minus 3.99565f
C6 source plus 4.00966f
C7 drain_left drain_right 1.01253f
C8 drain_left minus 0.17204f
C9 drain_left plus 4.04697f
C10 drain_right a_n2018_n2088# 4.93721f
C11 drain_left a_n2018_n2088# 5.23728f
C12 source a_n2018_n2088# 5.4814f
C13 minus a_n2018_n2088# 7.439296f
C14 plus a_n2018_n2088# 8.88491f
C15 drain_right.t10 a_n2018_n2088# 0.130309f
C16 drain_right.t1 a_n2018_n2088# 0.130309f
C17 drain_right.n0 a_n2018_n2088# 1.09086f
C18 drain_right.t0 a_n2018_n2088# 0.130309f
C19 drain_right.t7 a_n2018_n2088# 0.130309f
C20 drain_right.n1 a_n2018_n2088# 1.08678f
C21 drain_right.t2 a_n2018_n2088# 0.130309f
C22 drain_right.t3 a_n2018_n2088# 0.130309f
C23 drain_right.n2 a_n2018_n2088# 1.09086f
C24 drain_right.n3 a_n2018_n2088# 2.03177f
C25 drain_right.t5 a_n2018_n2088# 0.130309f
C26 drain_right.t4 a_n2018_n2088# 0.130309f
C27 drain_right.n4 a_n2018_n2088# 1.09121f
C28 drain_right.t8 a_n2018_n2088# 0.130309f
C29 drain_right.t6 a_n2018_n2088# 0.130309f
C30 drain_right.n5 a_n2018_n2088# 1.08678f
C31 drain_right.n6 a_n2018_n2088# 0.736752f
C32 drain_right.t9 a_n2018_n2088# 0.130309f
C33 drain_right.t11 a_n2018_n2088# 0.130309f
C34 drain_right.n7 a_n2018_n2088# 1.08678f
C35 drain_right.n8 a_n2018_n2088# 0.604709f
C36 minus.n0 a_n2018_n2088# 0.044764f
C37 minus.t3 a_n2018_n2088# 0.467428f
C38 minus.n1 a_n2018_n2088# 0.228313f
C39 minus.t0 a_n2018_n2088# 0.467428f
C40 minus.t7 a_n2018_n2088# 0.483882f
C41 minus.n2 a_n2018_n2088# 0.204634f
C42 minus.t6 a_n2018_n2088# 0.467428f
C43 minus.n3 a_n2018_n2088# 0.226678f
C44 minus.t5 a_n2018_n2088# 0.467428f
C45 minus.n4 a_n2018_n2088# 0.228313f
C46 minus.n5 a_n2018_n2088# 0.229423f
C47 minus.n6 a_n2018_n2088# 0.07456f
C48 minus.n7 a_n2018_n2088# 0.059732f
C49 minus.n8 a_n2018_n2088# 0.219673f
C50 minus.n9 a_n2018_n2088# 0.010158f
C51 minus.t2 a_n2018_n2088# 0.467428f
C52 minus.n10 a_n2018_n2088# 0.216637f
C53 minus.n11 a_n2018_n2088# 1.32191f
C54 minus.n12 a_n2018_n2088# 0.044764f
C55 minus.t4 a_n2018_n2088# 0.467428f
C56 minus.n13 a_n2018_n2088# 0.228313f
C57 minus.t1 a_n2018_n2088# 0.483882f
C58 minus.n14 a_n2018_n2088# 0.204634f
C59 minus.t10 a_n2018_n2088# 0.467428f
C60 minus.n15 a_n2018_n2088# 0.226678f
C61 minus.t11 a_n2018_n2088# 0.467428f
C62 minus.n16 a_n2018_n2088# 0.228313f
C63 minus.n17 a_n2018_n2088# 0.229423f
C64 minus.n18 a_n2018_n2088# 0.07456f
C65 minus.n19 a_n2018_n2088# 0.059732f
C66 minus.t9 a_n2018_n2088# 0.467428f
C67 minus.n20 a_n2018_n2088# 0.219673f
C68 minus.n21 a_n2018_n2088# 0.010158f
C69 minus.t8 a_n2018_n2088# 0.467428f
C70 minus.n22 a_n2018_n2088# 0.216637f
C71 minus.n23 a_n2018_n2088# 0.30186f
C72 minus.n24 a_n2018_n2088# 1.61902f
C73 source.n0 a_n2018_n2088# 0.034026f
C74 source.n1 a_n2018_n2088# 0.024208f
C75 source.n2 a_n2018_n2088# 0.013008f
C76 source.n3 a_n2018_n2088# 0.030747f
C77 source.n4 a_n2018_n2088# 0.013773f
C78 source.n5 a_n2018_n2088# 0.024208f
C79 source.n6 a_n2018_n2088# 0.013008f
C80 source.n7 a_n2018_n2088# 0.030747f
C81 source.n8 a_n2018_n2088# 0.013773f
C82 source.n9 a_n2018_n2088# 0.103592f
C83 source.t17 a_n2018_n2088# 0.050113f
C84 source.n10 a_n2018_n2088# 0.02306f
C85 source.n11 a_n2018_n2088# 0.018162f
C86 source.n12 a_n2018_n2088# 0.013008f
C87 source.n13 a_n2018_n2088# 0.576001f
C88 source.n14 a_n2018_n2088# 0.024208f
C89 source.n15 a_n2018_n2088# 0.013008f
C90 source.n16 a_n2018_n2088# 0.013773f
C91 source.n17 a_n2018_n2088# 0.030747f
C92 source.n18 a_n2018_n2088# 0.030747f
C93 source.n19 a_n2018_n2088# 0.013773f
C94 source.n20 a_n2018_n2088# 0.013008f
C95 source.n21 a_n2018_n2088# 0.024208f
C96 source.n22 a_n2018_n2088# 0.024208f
C97 source.n23 a_n2018_n2088# 0.013008f
C98 source.n24 a_n2018_n2088# 0.013773f
C99 source.n25 a_n2018_n2088# 0.030747f
C100 source.n26 a_n2018_n2088# 0.066561f
C101 source.n27 a_n2018_n2088# 0.013773f
C102 source.n28 a_n2018_n2088# 0.013008f
C103 source.n29 a_n2018_n2088# 0.055955f
C104 source.n30 a_n2018_n2088# 0.037244f
C105 source.n31 a_n2018_n2088# 0.620902f
C106 source.t12 a_n2018_n2088# 0.114778f
C107 source.t15 a_n2018_n2088# 0.114778f
C108 source.n32 a_n2018_n2088# 0.893904f
C109 source.n33 a_n2018_n2088# 0.351999f
C110 source.t10 a_n2018_n2088# 0.114778f
C111 source.t11 a_n2018_n2088# 0.114778f
C112 source.n34 a_n2018_n2088# 0.893904f
C113 source.n35 a_n2018_n2088# 0.351999f
C114 source.n36 a_n2018_n2088# 0.034026f
C115 source.n37 a_n2018_n2088# 0.024208f
C116 source.n38 a_n2018_n2088# 0.013008f
C117 source.n39 a_n2018_n2088# 0.030747f
C118 source.n40 a_n2018_n2088# 0.013773f
C119 source.n41 a_n2018_n2088# 0.024208f
C120 source.n42 a_n2018_n2088# 0.013008f
C121 source.n43 a_n2018_n2088# 0.030747f
C122 source.n44 a_n2018_n2088# 0.013773f
C123 source.n45 a_n2018_n2088# 0.103592f
C124 source.t9 a_n2018_n2088# 0.050113f
C125 source.n46 a_n2018_n2088# 0.02306f
C126 source.n47 a_n2018_n2088# 0.018162f
C127 source.n48 a_n2018_n2088# 0.013008f
C128 source.n49 a_n2018_n2088# 0.576001f
C129 source.n50 a_n2018_n2088# 0.024208f
C130 source.n51 a_n2018_n2088# 0.013008f
C131 source.n52 a_n2018_n2088# 0.013773f
C132 source.n53 a_n2018_n2088# 0.030747f
C133 source.n54 a_n2018_n2088# 0.030747f
C134 source.n55 a_n2018_n2088# 0.013773f
C135 source.n56 a_n2018_n2088# 0.013008f
C136 source.n57 a_n2018_n2088# 0.024208f
C137 source.n58 a_n2018_n2088# 0.024208f
C138 source.n59 a_n2018_n2088# 0.013008f
C139 source.n60 a_n2018_n2088# 0.013773f
C140 source.n61 a_n2018_n2088# 0.030747f
C141 source.n62 a_n2018_n2088# 0.066561f
C142 source.n63 a_n2018_n2088# 0.013773f
C143 source.n64 a_n2018_n2088# 0.013008f
C144 source.n65 a_n2018_n2088# 0.055955f
C145 source.n66 a_n2018_n2088# 0.037244f
C146 source.n67 a_n2018_n2088# 0.11986f
C147 source.n68 a_n2018_n2088# 0.034026f
C148 source.n69 a_n2018_n2088# 0.024208f
C149 source.n70 a_n2018_n2088# 0.013008f
C150 source.n71 a_n2018_n2088# 0.030747f
C151 source.n72 a_n2018_n2088# 0.013773f
C152 source.n73 a_n2018_n2088# 0.024208f
C153 source.n74 a_n2018_n2088# 0.013008f
C154 source.n75 a_n2018_n2088# 0.030747f
C155 source.n76 a_n2018_n2088# 0.013773f
C156 source.n77 a_n2018_n2088# 0.103592f
C157 source.t3 a_n2018_n2088# 0.050113f
C158 source.n78 a_n2018_n2088# 0.02306f
C159 source.n79 a_n2018_n2088# 0.018162f
C160 source.n80 a_n2018_n2088# 0.013008f
C161 source.n81 a_n2018_n2088# 0.576001f
C162 source.n82 a_n2018_n2088# 0.024208f
C163 source.n83 a_n2018_n2088# 0.013008f
C164 source.n84 a_n2018_n2088# 0.013773f
C165 source.n85 a_n2018_n2088# 0.030747f
C166 source.n86 a_n2018_n2088# 0.030747f
C167 source.n87 a_n2018_n2088# 0.013773f
C168 source.n88 a_n2018_n2088# 0.013008f
C169 source.n89 a_n2018_n2088# 0.024208f
C170 source.n90 a_n2018_n2088# 0.024208f
C171 source.n91 a_n2018_n2088# 0.013008f
C172 source.n92 a_n2018_n2088# 0.013773f
C173 source.n93 a_n2018_n2088# 0.030747f
C174 source.n94 a_n2018_n2088# 0.066561f
C175 source.n95 a_n2018_n2088# 0.013773f
C176 source.n96 a_n2018_n2088# 0.013008f
C177 source.n97 a_n2018_n2088# 0.055955f
C178 source.n98 a_n2018_n2088# 0.037244f
C179 source.n99 a_n2018_n2088# 0.11986f
C180 source.t23 a_n2018_n2088# 0.114778f
C181 source.t4 a_n2018_n2088# 0.114778f
C182 source.n100 a_n2018_n2088# 0.893904f
C183 source.n101 a_n2018_n2088# 0.351999f
C184 source.t0 a_n2018_n2088# 0.114778f
C185 source.t21 a_n2018_n2088# 0.114778f
C186 source.n102 a_n2018_n2088# 0.893904f
C187 source.n103 a_n2018_n2088# 0.351999f
C188 source.n104 a_n2018_n2088# 0.034026f
C189 source.n105 a_n2018_n2088# 0.024208f
C190 source.n106 a_n2018_n2088# 0.013008f
C191 source.n107 a_n2018_n2088# 0.030747f
C192 source.n108 a_n2018_n2088# 0.013773f
C193 source.n109 a_n2018_n2088# 0.024208f
C194 source.n110 a_n2018_n2088# 0.013008f
C195 source.n111 a_n2018_n2088# 0.030747f
C196 source.n112 a_n2018_n2088# 0.013773f
C197 source.n113 a_n2018_n2088# 0.103592f
C198 source.t20 a_n2018_n2088# 0.050113f
C199 source.n114 a_n2018_n2088# 0.02306f
C200 source.n115 a_n2018_n2088# 0.018162f
C201 source.n116 a_n2018_n2088# 0.013008f
C202 source.n117 a_n2018_n2088# 0.576001f
C203 source.n118 a_n2018_n2088# 0.024208f
C204 source.n119 a_n2018_n2088# 0.013008f
C205 source.n120 a_n2018_n2088# 0.013773f
C206 source.n121 a_n2018_n2088# 0.030747f
C207 source.n122 a_n2018_n2088# 0.030747f
C208 source.n123 a_n2018_n2088# 0.013773f
C209 source.n124 a_n2018_n2088# 0.013008f
C210 source.n125 a_n2018_n2088# 0.024208f
C211 source.n126 a_n2018_n2088# 0.024208f
C212 source.n127 a_n2018_n2088# 0.013008f
C213 source.n128 a_n2018_n2088# 0.013773f
C214 source.n129 a_n2018_n2088# 0.030747f
C215 source.n130 a_n2018_n2088# 0.066561f
C216 source.n131 a_n2018_n2088# 0.013773f
C217 source.n132 a_n2018_n2088# 0.013008f
C218 source.n133 a_n2018_n2088# 0.055955f
C219 source.n134 a_n2018_n2088# 0.037244f
C220 source.n135 a_n2018_n2088# 0.938358f
C221 source.n136 a_n2018_n2088# 0.034026f
C222 source.n137 a_n2018_n2088# 0.024208f
C223 source.n138 a_n2018_n2088# 0.013008f
C224 source.n139 a_n2018_n2088# 0.030747f
C225 source.n140 a_n2018_n2088# 0.013773f
C226 source.n141 a_n2018_n2088# 0.024208f
C227 source.n142 a_n2018_n2088# 0.013008f
C228 source.n143 a_n2018_n2088# 0.030747f
C229 source.n144 a_n2018_n2088# 0.013773f
C230 source.n145 a_n2018_n2088# 0.103592f
C231 source.t7 a_n2018_n2088# 0.050113f
C232 source.n146 a_n2018_n2088# 0.02306f
C233 source.n147 a_n2018_n2088# 0.018162f
C234 source.n148 a_n2018_n2088# 0.013008f
C235 source.n149 a_n2018_n2088# 0.576001f
C236 source.n150 a_n2018_n2088# 0.024208f
C237 source.n151 a_n2018_n2088# 0.013008f
C238 source.n152 a_n2018_n2088# 0.013773f
C239 source.n153 a_n2018_n2088# 0.030747f
C240 source.n154 a_n2018_n2088# 0.030747f
C241 source.n155 a_n2018_n2088# 0.013773f
C242 source.n156 a_n2018_n2088# 0.013008f
C243 source.n157 a_n2018_n2088# 0.024208f
C244 source.n158 a_n2018_n2088# 0.024208f
C245 source.n159 a_n2018_n2088# 0.013008f
C246 source.n160 a_n2018_n2088# 0.013773f
C247 source.n161 a_n2018_n2088# 0.030747f
C248 source.n162 a_n2018_n2088# 0.066561f
C249 source.n163 a_n2018_n2088# 0.013773f
C250 source.n164 a_n2018_n2088# 0.013008f
C251 source.n165 a_n2018_n2088# 0.055955f
C252 source.n166 a_n2018_n2088# 0.037244f
C253 source.n167 a_n2018_n2088# 0.938358f
C254 source.t8 a_n2018_n2088# 0.114778f
C255 source.t13 a_n2018_n2088# 0.114778f
C256 source.n168 a_n2018_n2088# 0.893898f
C257 source.n169 a_n2018_n2088# 0.352005f
C258 source.t16 a_n2018_n2088# 0.114778f
C259 source.t18 a_n2018_n2088# 0.114778f
C260 source.n170 a_n2018_n2088# 0.893898f
C261 source.n171 a_n2018_n2088# 0.352005f
C262 source.n172 a_n2018_n2088# 0.034026f
C263 source.n173 a_n2018_n2088# 0.024208f
C264 source.n174 a_n2018_n2088# 0.013008f
C265 source.n175 a_n2018_n2088# 0.030747f
C266 source.n176 a_n2018_n2088# 0.013773f
C267 source.n177 a_n2018_n2088# 0.024208f
C268 source.n178 a_n2018_n2088# 0.013008f
C269 source.n179 a_n2018_n2088# 0.030747f
C270 source.n180 a_n2018_n2088# 0.013773f
C271 source.n181 a_n2018_n2088# 0.103592f
C272 source.t14 a_n2018_n2088# 0.050113f
C273 source.n182 a_n2018_n2088# 0.02306f
C274 source.n183 a_n2018_n2088# 0.018162f
C275 source.n184 a_n2018_n2088# 0.013008f
C276 source.n185 a_n2018_n2088# 0.576001f
C277 source.n186 a_n2018_n2088# 0.024208f
C278 source.n187 a_n2018_n2088# 0.013008f
C279 source.n188 a_n2018_n2088# 0.013773f
C280 source.n189 a_n2018_n2088# 0.030747f
C281 source.n190 a_n2018_n2088# 0.030747f
C282 source.n191 a_n2018_n2088# 0.013773f
C283 source.n192 a_n2018_n2088# 0.013008f
C284 source.n193 a_n2018_n2088# 0.024208f
C285 source.n194 a_n2018_n2088# 0.024208f
C286 source.n195 a_n2018_n2088# 0.013008f
C287 source.n196 a_n2018_n2088# 0.013773f
C288 source.n197 a_n2018_n2088# 0.030747f
C289 source.n198 a_n2018_n2088# 0.066561f
C290 source.n199 a_n2018_n2088# 0.013773f
C291 source.n200 a_n2018_n2088# 0.013008f
C292 source.n201 a_n2018_n2088# 0.055955f
C293 source.n202 a_n2018_n2088# 0.037244f
C294 source.n203 a_n2018_n2088# 0.11986f
C295 source.n204 a_n2018_n2088# 0.034026f
C296 source.n205 a_n2018_n2088# 0.024208f
C297 source.n206 a_n2018_n2088# 0.013008f
C298 source.n207 a_n2018_n2088# 0.030747f
C299 source.n208 a_n2018_n2088# 0.013773f
C300 source.n209 a_n2018_n2088# 0.024208f
C301 source.n210 a_n2018_n2088# 0.013008f
C302 source.n211 a_n2018_n2088# 0.030747f
C303 source.n212 a_n2018_n2088# 0.013773f
C304 source.n213 a_n2018_n2088# 0.103592f
C305 source.t2 a_n2018_n2088# 0.050113f
C306 source.n214 a_n2018_n2088# 0.02306f
C307 source.n215 a_n2018_n2088# 0.018162f
C308 source.n216 a_n2018_n2088# 0.013008f
C309 source.n217 a_n2018_n2088# 0.576001f
C310 source.n218 a_n2018_n2088# 0.024208f
C311 source.n219 a_n2018_n2088# 0.013008f
C312 source.n220 a_n2018_n2088# 0.013773f
C313 source.n221 a_n2018_n2088# 0.030747f
C314 source.n222 a_n2018_n2088# 0.030747f
C315 source.n223 a_n2018_n2088# 0.013773f
C316 source.n224 a_n2018_n2088# 0.013008f
C317 source.n225 a_n2018_n2088# 0.024208f
C318 source.n226 a_n2018_n2088# 0.024208f
C319 source.n227 a_n2018_n2088# 0.013008f
C320 source.n228 a_n2018_n2088# 0.013773f
C321 source.n229 a_n2018_n2088# 0.030747f
C322 source.n230 a_n2018_n2088# 0.066561f
C323 source.n231 a_n2018_n2088# 0.013773f
C324 source.n232 a_n2018_n2088# 0.013008f
C325 source.n233 a_n2018_n2088# 0.055955f
C326 source.n234 a_n2018_n2088# 0.037244f
C327 source.n235 a_n2018_n2088# 0.11986f
C328 source.t19 a_n2018_n2088# 0.114778f
C329 source.t1 a_n2018_n2088# 0.114778f
C330 source.n236 a_n2018_n2088# 0.893898f
C331 source.n237 a_n2018_n2088# 0.352005f
C332 source.t22 a_n2018_n2088# 0.114778f
C333 source.t5 a_n2018_n2088# 0.114778f
C334 source.n238 a_n2018_n2088# 0.893898f
C335 source.n239 a_n2018_n2088# 0.352005f
C336 source.n240 a_n2018_n2088# 0.034026f
C337 source.n241 a_n2018_n2088# 0.024208f
C338 source.n242 a_n2018_n2088# 0.013008f
C339 source.n243 a_n2018_n2088# 0.030747f
C340 source.n244 a_n2018_n2088# 0.013773f
C341 source.n245 a_n2018_n2088# 0.024208f
C342 source.n246 a_n2018_n2088# 0.013008f
C343 source.n247 a_n2018_n2088# 0.030747f
C344 source.n248 a_n2018_n2088# 0.013773f
C345 source.n249 a_n2018_n2088# 0.103592f
C346 source.t6 a_n2018_n2088# 0.050113f
C347 source.n250 a_n2018_n2088# 0.02306f
C348 source.n251 a_n2018_n2088# 0.018162f
C349 source.n252 a_n2018_n2088# 0.013008f
C350 source.n253 a_n2018_n2088# 0.576001f
C351 source.n254 a_n2018_n2088# 0.024208f
C352 source.n255 a_n2018_n2088# 0.013008f
C353 source.n256 a_n2018_n2088# 0.013773f
C354 source.n257 a_n2018_n2088# 0.030747f
C355 source.n258 a_n2018_n2088# 0.030747f
C356 source.n259 a_n2018_n2088# 0.013773f
C357 source.n260 a_n2018_n2088# 0.013008f
C358 source.n261 a_n2018_n2088# 0.024208f
C359 source.n262 a_n2018_n2088# 0.024208f
C360 source.n263 a_n2018_n2088# 0.013008f
C361 source.n264 a_n2018_n2088# 0.013773f
C362 source.n265 a_n2018_n2088# 0.030747f
C363 source.n266 a_n2018_n2088# 0.066561f
C364 source.n267 a_n2018_n2088# 0.013773f
C365 source.n268 a_n2018_n2088# 0.013008f
C366 source.n269 a_n2018_n2088# 0.055955f
C367 source.n270 a_n2018_n2088# 0.037244f
C368 source.n271 a_n2018_n2088# 0.272499f
C369 source.n272 a_n2018_n2088# 1.00053f
C370 drain_left.t11 a_n2018_n2088# 0.131195f
C371 drain_left.t10 a_n2018_n2088# 0.131195f
C372 drain_left.n0 a_n2018_n2088# 1.09828f
C373 drain_left.t5 a_n2018_n2088# 0.131195f
C374 drain_left.t2 a_n2018_n2088# 0.131195f
C375 drain_left.n1 a_n2018_n2088# 1.09416f
C376 drain_left.t0 a_n2018_n2088# 0.131195f
C377 drain_left.t4 a_n2018_n2088# 0.131195f
C378 drain_left.n2 a_n2018_n2088# 1.09828f
C379 drain_left.n3 a_n2018_n2088# 2.1016f
C380 drain_left.t9 a_n2018_n2088# 0.131195f
C381 drain_left.t8 a_n2018_n2088# 0.131195f
C382 drain_left.n4 a_n2018_n2088# 1.09863f
C383 drain_left.t7 a_n2018_n2088# 0.131195f
C384 drain_left.t6 a_n2018_n2088# 0.131195f
C385 drain_left.n5 a_n2018_n2088# 1.09417f
C386 drain_left.n6 a_n2018_n2088# 0.741755f
C387 drain_left.t3 a_n2018_n2088# 0.131195f
C388 drain_left.t1 a_n2018_n2088# 0.131195f
C389 drain_left.n7 a_n2018_n2088# 1.09416f
C390 drain_left.n8 a_n2018_n2088# 0.608824f
C391 plus.n0 a_n2018_n2088# 0.045821f
C392 plus.t1 a_n2018_n2088# 0.47846f
C393 plus.t3 a_n2018_n2088# 0.47846f
C394 plus.n1 a_n2018_n2088# 0.061142f
C395 plus.t6 a_n2018_n2088# 0.47846f
C396 plus.n2 a_n2018_n2088# 0.07632f
C397 plus.t7 a_n2018_n2088# 0.47846f
C398 plus.n3 a_n2018_n2088# 0.234838f
C399 plus.t8 a_n2018_n2088# 0.47846f
C400 plus.t9 a_n2018_n2088# 0.495302f
C401 plus.n4 a_n2018_n2088# 0.209464f
C402 plus.n5 a_n2018_n2088# 0.232028f
C403 plus.n6 a_n2018_n2088# 0.233701f
C404 plus.n7 a_n2018_n2088# 0.233701f
C405 plus.n8 a_n2018_n2088# 0.224857f
C406 plus.n9 a_n2018_n2088# 0.010398f
C407 plus.n10 a_n2018_n2088# 0.22175f
C408 plus.n11 a_n2018_n2088# 0.402472f
C409 plus.n12 a_n2018_n2088# 0.045821f
C410 plus.t11 a_n2018_n2088# 0.47846f
C411 plus.n13 a_n2018_n2088# 0.061142f
C412 plus.t10 a_n2018_n2088# 0.47846f
C413 plus.n14 a_n2018_n2088# 0.07632f
C414 plus.t5 a_n2018_n2088# 0.47846f
C415 plus.n15 a_n2018_n2088# 0.234838f
C416 plus.t2 a_n2018_n2088# 0.47846f
C417 plus.t4 a_n2018_n2088# 0.495302f
C418 plus.n16 a_n2018_n2088# 0.209464f
C419 plus.t0 a_n2018_n2088# 0.47846f
C420 plus.n17 a_n2018_n2088# 0.232028f
C421 plus.n18 a_n2018_n2088# 0.233701f
C422 plus.n19 a_n2018_n2088# 0.233701f
C423 plus.n20 a_n2018_n2088# 0.224857f
C424 plus.n21 a_n2018_n2088# 0.010398f
C425 plus.n22 a_n2018_n2088# 0.22175f
C426 plus.n23 a_n2018_n2088# 1.22324f
.ends

