* NGSPICE file created from diffpair371.ext - technology: sky130A

.subckt diffpair371 minus drain_right drain_left source plus
X0 a_n1274_n2688# a_n1274_n2688# a_n1274_n2688# a_n1274_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.6
X1 a_n1274_n2688# a_n1274_n2688# a_n1274_n2688# a_n1274_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X2 a_n1274_n2688# a_n1274_n2688# a_n1274_n2688# a_n1274_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X3 source plus drain_left a_n1274_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X4 source minus drain_right a_n1274_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X5 a_n1274_n2688# a_n1274_n2688# a_n1274_n2688# a_n1274_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X6 source minus drain_right a_n1274_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X7 drain_right minus source a_n1274_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X8 drain_left plus source a_n1274_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X9 source plus drain_left a_n1274_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X10 drain_left plus source a_n1274_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X11 drain_right minus source a_n1274_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
.ends

