* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t32 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X1 a_n2762_n1088# a_n2762_n1088# a_n2762_n1088# a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.6
X2 drain_left.t18 plus.t1 source.t26 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X3 source.t31 plus.t2 drain_left.t17 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X4 drain_left.t16 plus.t3 source.t33 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X5 source.t17 minus.t0 drain_right.t19 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X6 source.t28 plus.t4 drain_left.t15 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X7 source.t22 plus.t5 drain_left.t14 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X8 drain_right.t18 minus.t1 source.t39 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X9 drain_left.t13 plus.t6 source.t19 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X10 source.t18 minus.t2 drain_right.t17 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X11 drain_right.t16 minus.t3 source.t16 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X12 drain_right.t15 minus.t4 source.t14 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X13 drain_right.t14 minus.t5 source.t15 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X14 source.t1 minus.t6 drain_right.t13 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X15 source.t7 minus.t7 drain_right.t12 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X16 source.t23 plus.t7 drain_left.t12 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X17 a_n2762_n1088# a_n2762_n1088# a_n2762_n1088# a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X18 a_n2762_n1088# a_n2762_n1088# a_n2762_n1088# a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X19 source.t11 minus.t8 drain_right.t11 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X20 drain_right.t10 minus.t9 source.t9 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X21 source.t24 plus.t8 drain_left.t11 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X22 source.t38 plus.t9 drain_left.t10 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X23 source.t0 minus.t10 drain_right.t9 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X24 drain_right.t8 minus.t11 source.t6 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X25 drain_left.t9 plus.t10 source.t29 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X26 drain_left.t8 plus.t11 source.t20 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X27 source.t10 minus.t12 drain_right.t7 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X28 drain_left.t7 plus.t12 source.t36 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X29 source.t27 plus.t13 drain_left.t6 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X30 drain_right.t6 minus.t13 source.t8 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X31 drain_right.t5 minus.t14 source.t5 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X32 drain_left.t5 plus.t14 source.t21 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X33 drain_left.t4 plus.t15 source.t30 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X34 source.t37 plus.t16 drain_left.t3 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X35 source.t4 minus.t15 drain_right.t4 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X36 source.t34 plus.t17 drain_left.t2 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X37 source.t3 minus.t16 drain_right.t3 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X38 drain_right.t2 minus.t17 source.t2 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X39 source.t25 plus.t18 drain_left.t1 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X40 drain_right.t1 minus.t18 source.t12 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X41 source.t13 minus.t19 drain_right.t0 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X42 a_n2762_n1088# a_n2762_n1088# a_n2762_n1088# a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X43 drain_left.t0 plus.t19 source.t35 a_n2762_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
R0 plus.n9 plus.n6 161.3
R1 plus.n11 plus.n10 161.3
R2 plus.n12 plus.n5 161.3
R3 plus.n14 plus.n13 161.3
R4 plus.n15 plus.n4 161.3
R5 plus.n17 plus.n16 161.3
R6 plus.n18 plus.n3 161.3
R7 plus.n20 plus.n19 161.3
R8 plus.n21 plus.n2 161.3
R9 plus.n23 plus.n22 161.3
R10 plus.n24 plus.n1 161.3
R11 plus.n27 plus.n26 161.3
R12 plus.n37 plus.n34 161.3
R13 plus.n39 plus.n38 161.3
R14 plus.n40 plus.n33 161.3
R15 plus.n42 plus.n41 161.3
R16 plus.n43 plus.n32 161.3
R17 plus.n45 plus.n44 161.3
R18 plus.n46 plus.n31 161.3
R19 plus.n48 plus.n47 161.3
R20 plus.n49 plus.n30 161.3
R21 plus.n51 plus.n50 161.3
R22 plus.n52 plus.n29 161.3
R23 plus.n55 plus.n54 161.3
R24 plus.n8 plus.t16 132.459
R25 plus.n36 plus.t10 132.459
R26 plus.n26 plus.t0 105.638
R27 plus.n25 plus.t2 105.638
R28 plus.n24 plus.t3 105.638
R29 plus.n2 plus.t5 105.638
R30 plus.n18 plus.t6 105.638
R31 plus.n4 plus.t9 105.638
R32 plus.n12 plus.t11 105.638
R33 plus.n6 plus.t13 105.638
R34 plus.n7 plus.t15 105.638
R35 plus.n54 plus.t7 105.638
R36 plus.n53 plus.t14 105.638
R37 plus.n52 plus.t18 105.638
R38 plus.n30 plus.t1 105.638
R39 plus.n46 plus.t8 105.638
R40 plus.n32 plus.t12 105.638
R41 plus.n40 plus.t17 105.638
R42 plus.n34 plus.t19 105.638
R43 plus.n35 plus.t4 105.638
R44 plus.n25 plus.n0 80.6037
R45 plus.n53 plus.n28 80.6037
R46 plus.n26 plus.n25 48.2005
R47 plus.n25 plus.n24 48.2005
R48 plus.n7 plus.n6 48.2005
R49 plus.n54 plus.n53 48.2005
R50 plus.n53 plus.n52 48.2005
R51 plus.n35 plus.n34 48.2005
R52 plus.n9 plus.n8 45.1367
R53 plus.n37 plus.n36 45.1367
R54 plus.n23 plus.n2 44.549
R55 plus.n12 plus.n11 44.549
R56 plus.n51 plus.n30 44.549
R57 plus.n40 plus.n39 44.549
R58 plus.n19 plus.n18 34.3247
R59 plus.n13 plus.n4 34.3247
R60 plus.n47 plus.n46 34.3247
R61 plus.n41 plus.n32 34.3247
R62 plus plus.n55 29.4271
R63 plus.n17 plus.n4 24.1005
R64 plus.n18 plus.n17 24.1005
R65 plus.n46 plus.n45 24.1005
R66 plus.n45 plus.n32 24.1005
R67 plus.n19 plus.n2 13.8763
R68 plus.n13 plus.n12 13.8763
R69 plus.n47 plus.n30 13.8763
R70 plus.n41 plus.n40 13.8763
R71 plus.n8 plus.n7 13.3799
R72 plus.n36 plus.n35 13.3799
R73 plus plus.n27 8.10656
R74 plus.n24 plus.n23 3.65202
R75 plus.n11 plus.n6 3.65202
R76 plus.n52 plus.n51 3.65202
R77 plus.n39 plus.n34 3.65202
R78 plus.n1 plus.n0 0.285035
R79 plus.n27 plus.n0 0.285035
R80 plus.n55 plus.n28 0.285035
R81 plus.n29 plus.n28 0.285035
R82 plus.n10 plus.n9 0.189894
R83 plus.n10 plus.n5 0.189894
R84 plus.n14 plus.n5 0.189894
R85 plus.n15 plus.n14 0.189894
R86 plus.n16 plus.n15 0.189894
R87 plus.n16 plus.n3 0.189894
R88 plus.n20 plus.n3 0.189894
R89 plus.n21 plus.n20 0.189894
R90 plus.n22 plus.n21 0.189894
R91 plus.n22 plus.n1 0.189894
R92 plus.n50 plus.n29 0.189894
R93 plus.n50 plus.n49 0.189894
R94 plus.n49 plus.n48 0.189894
R95 plus.n48 plus.n31 0.189894
R96 plus.n44 plus.n31 0.189894
R97 plus.n44 plus.n43 0.189894
R98 plus.n43 plus.n42 0.189894
R99 plus.n42 plus.n33 0.189894
R100 plus.n38 plus.n33 0.189894
R101 plus.n38 plus.n37 0.189894
R102 source.n0 source.t32 243.255
R103 source.n9 source.t37 243.255
R104 source.n10 source.t8 243.255
R105 source.n19 source.t17 243.255
R106 source.n39 source.t5 243.254
R107 source.n30 source.t13 243.254
R108 source.n29 source.t29 243.254
R109 source.n20 source.t23 243.254
R110 source.n2 source.n1 223.454
R111 source.n4 source.n3 223.454
R112 source.n6 source.n5 223.454
R113 source.n8 source.n7 223.454
R114 source.n12 source.n11 223.454
R115 source.n14 source.n13 223.454
R116 source.n16 source.n15 223.454
R117 source.n18 source.n17 223.454
R118 source.n38 source.n37 223.453
R119 source.n36 source.n35 223.453
R120 source.n34 source.n33 223.453
R121 source.n32 source.n31 223.453
R122 source.n28 source.n27 223.453
R123 source.n26 source.n25 223.453
R124 source.n24 source.n23 223.453
R125 source.n22 source.n21 223.453
R126 source.n37 source.t15 19.8005
R127 source.n37 source.t3 19.8005
R128 source.n35 source.t2 19.8005
R129 source.n35 source.t11 19.8005
R130 source.n33 source.t12 19.8005
R131 source.n33 source.t4 19.8005
R132 source.n31 source.t9 19.8005
R133 source.n31 source.t7 19.8005
R134 source.n27 source.t35 19.8005
R135 source.n27 source.t28 19.8005
R136 source.n25 source.t36 19.8005
R137 source.n25 source.t34 19.8005
R138 source.n23 source.t26 19.8005
R139 source.n23 source.t24 19.8005
R140 source.n21 source.t21 19.8005
R141 source.n21 source.t25 19.8005
R142 source.n1 source.t33 19.8005
R143 source.n1 source.t31 19.8005
R144 source.n3 source.t19 19.8005
R145 source.n3 source.t22 19.8005
R146 source.n5 source.t20 19.8005
R147 source.n5 source.t38 19.8005
R148 source.n7 source.t30 19.8005
R149 source.n7 source.t27 19.8005
R150 source.n11 source.t6 19.8005
R151 source.n11 source.t10 19.8005
R152 source.n13 source.t16 19.8005
R153 source.n13 source.t0 19.8005
R154 source.n15 source.t14 19.8005
R155 source.n15 source.t1 19.8005
R156 source.n17 source.t39 19.8005
R157 source.n17 source.t18 19.8005
R158 source.n20 source.n19 13.7561
R159 source.n40 source.n0 8.09232
R160 source.n40 source.n39 5.66429
R161 source.n19 source.n18 0.802224
R162 source.n18 source.n16 0.802224
R163 source.n16 source.n14 0.802224
R164 source.n14 source.n12 0.802224
R165 source.n12 source.n10 0.802224
R166 source.n9 source.n8 0.802224
R167 source.n8 source.n6 0.802224
R168 source.n6 source.n4 0.802224
R169 source.n4 source.n2 0.802224
R170 source.n2 source.n0 0.802224
R171 source.n22 source.n20 0.802224
R172 source.n24 source.n22 0.802224
R173 source.n26 source.n24 0.802224
R174 source.n28 source.n26 0.802224
R175 source.n29 source.n28 0.802224
R176 source.n32 source.n30 0.802224
R177 source.n34 source.n32 0.802224
R178 source.n36 source.n34 0.802224
R179 source.n38 source.n36 0.802224
R180 source.n39 source.n38 0.802224
R181 source.n10 source.n9 0.470328
R182 source.n30 source.n29 0.470328
R183 source source.n40 0.188
R184 drain_left.n10 drain_left.n8 240.935
R185 drain_left.n6 drain_left.n4 240.934
R186 drain_left.n2 drain_left.n0 240.934
R187 drain_left.n16 drain_left.n15 240.132
R188 drain_left.n14 drain_left.n13 240.132
R189 drain_left.n12 drain_left.n11 240.132
R190 drain_left.n10 drain_left.n9 240.132
R191 drain_left.n7 drain_left.n3 240.131
R192 drain_left.n6 drain_left.n5 240.131
R193 drain_left.n2 drain_left.n1 240.131
R194 drain_left drain_left.n7 25.4475
R195 drain_left.n3 drain_left.t11 19.8005
R196 drain_left.n3 drain_left.t7 19.8005
R197 drain_left.n4 drain_left.t15 19.8005
R198 drain_left.n4 drain_left.t9 19.8005
R199 drain_left.n5 drain_left.t2 19.8005
R200 drain_left.n5 drain_left.t0 19.8005
R201 drain_left.n1 drain_left.t1 19.8005
R202 drain_left.n1 drain_left.t18 19.8005
R203 drain_left.n0 drain_left.t12 19.8005
R204 drain_left.n0 drain_left.t5 19.8005
R205 drain_left.n15 drain_left.t17 19.8005
R206 drain_left.n15 drain_left.t19 19.8005
R207 drain_left.n13 drain_left.t14 19.8005
R208 drain_left.n13 drain_left.t16 19.8005
R209 drain_left.n11 drain_left.t10 19.8005
R210 drain_left.n11 drain_left.t13 19.8005
R211 drain_left.n9 drain_left.t6 19.8005
R212 drain_left.n9 drain_left.t8 19.8005
R213 drain_left.n8 drain_left.t3 19.8005
R214 drain_left.n8 drain_left.t4 19.8005
R215 drain_left drain_left.n16 6.45494
R216 drain_left.n12 drain_left.n10 0.802224
R217 drain_left.n14 drain_left.n12 0.802224
R218 drain_left.n16 drain_left.n14 0.802224
R219 drain_left.n7 drain_left.n6 0.746878
R220 drain_left.n7 drain_left.n2 0.746878
R221 minus.n27 minus.n26 161.3
R222 minus.n24 minus.n23 161.3
R223 minus.n22 minus.n1 161.3
R224 minus.n21 minus.n20 161.3
R225 minus.n19 minus.n2 161.3
R226 minus.n18 minus.n17 161.3
R227 minus.n16 minus.n3 161.3
R228 minus.n15 minus.n14 161.3
R229 minus.n13 minus.n4 161.3
R230 minus.n12 minus.n11 161.3
R231 minus.n10 minus.n5 161.3
R232 minus.n9 minus.n8 161.3
R233 minus.n55 minus.n54 161.3
R234 minus.n52 minus.n51 161.3
R235 minus.n50 minus.n29 161.3
R236 minus.n49 minus.n48 161.3
R237 minus.n47 minus.n30 161.3
R238 minus.n46 minus.n45 161.3
R239 minus.n44 minus.n31 161.3
R240 minus.n43 minus.n42 161.3
R241 minus.n41 minus.n32 161.3
R242 minus.n40 minus.n39 161.3
R243 minus.n38 minus.n33 161.3
R244 minus.n37 minus.n36 161.3
R245 minus.n6 minus.t13 132.459
R246 minus.n34 minus.t19 132.459
R247 minus.n7 minus.t12 105.638
R248 minus.n8 minus.t11 105.638
R249 minus.n12 minus.t10 105.638
R250 minus.n14 minus.t3 105.638
R251 minus.n18 minus.t6 105.638
R252 minus.n20 minus.t4 105.638
R253 minus.n24 minus.t2 105.638
R254 minus.n25 minus.t1 105.638
R255 minus.n26 minus.t0 105.638
R256 minus.n35 minus.t9 105.638
R257 minus.n36 minus.t7 105.638
R258 minus.n40 minus.t18 105.638
R259 minus.n42 minus.t15 105.638
R260 minus.n46 minus.t17 105.638
R261 minus.n48 minus.t8 105.638
R262 minus.n52 minus.t5 105.638
R263 minus.n53 minus.t16 105.638
R264 minus.n54 minus.t14 105.638
R265 minus.n25 minus.n0 80.6037
R266 minus.n53 minus.n28 80.6037
R267 minus.n8 minus.n7 48.2005
R268 minus.n25 minus.n24 48.2005
R269 minus.n26 minus.n25 48.2005
R270 minus.n36 minus.n35 48.2005
R271 minus.n53 minus.n52 48.2005
R272 minus.n54 minus.n53 48.2005
R273 minus.n9 minus.n6 45.1367
R274 minus.n37 minus.n34 45.1367
R275 minus.n12 minus.n5 44.549
R276 minus.n20 minus.n1 44.549
R277 minus.n40 minus.n33 44.549
R278 minus.n48 minus.n29 44.549
R279 minus.n14 minus.n13 34.3247
R280 minus.n19 minus.n18 34.3247
R281 minus.n42 minus.n41 34.3247
R282 minus.n47 minus.n46 34.3247
R283 minus.n56 minus.n27 31.3793
R284 minus.n18 minus.n3 24.1005
R285 minus.n14 minus.n3 24.1005
R286 minus.n42 minus.n31 24.1005
R287 minus.n46 minus.n31 24.1005
R288 minus.n13 minus.n12 13.8763
R289 minus.n20 minus.n19 13.8763
R290 minus.n41 minus.n40 13.8763
R291 minus.n48 minus.n47 13.8763
R292 minus.n7 minus.n6 13.3799
R293 minus.n35 minus.n34 13.3799
R294 minus.n56 minus.n55 6.62929
R295 minus.n8 minus.n5 3.65202
R296 minus.n24 minus.n1 3.65202
R297 minus.n36 minus.n33 3.65202
R298 minus.n52 minus.n29 3.65202
R299 minus.n27 minus.n0 0.285035
R300 minus.n23 minus.n0 0.285035
R301 minus.n51 minus.n28 0.285035
R302 minus.n55 minus.n28 0.285035
R303 minus.n23 minus.n22 0.189894
R304 minus.n22 minus.n21 0.189894
R305 minus.n21 minus.n2 0.189894
R306 minus.n17 minus.n2 0.189894
R307 minus.n17 minus.n16 0.189894
R308 minus.n16 minus.n15 0.189894
R309 minus.n15 minus.n4 0.189894
R310 minus.n11 minus.n4 0.189894
R311 minus.n11 minus.n10 0.189894
R312 minus.n10 minus.n9 0.189894
R313 minus.n38 minus.n37 0.189894
R314 minus.n39 minus.n38 0.189894
R315 minus.n39 minus.n32 0.189894
R316 minus.n43 minus.n32 0.189894
R317 minus.n44 minus.n43 0.189894
R318 minus.n45 minus.n44 0.189894
R319 minus.n45 minus.n30 0.189894
R320 minus.n49 minus.n30 0.189894
R321 minus.n50 minus.n49 0.189894
R322 minus.n51 minus.n50 0.189894
R323 minus minus.n56 0.188
R324 drain_right.n10 drain_right.n8 240.935
R325 drain_right.n6 drain_right.n4 240.934
R326 drain_right.n2 drain_right.n0 240.934
R327 drain_right.n10 drain_right.n9 240.132
R328 drain_right.n12 drain_right.n11 240.132
R329 drain_right.n14 drain_right.n13 240.132
R330 drain_right.n16 drain_right.n15 240.132
R331 drain_right.n7 drain_right.n3 240.131
R332 drain_right.n6 drain_right.n5 240.131
R333 drain_right.n2 drain_right.n1 240.131
R334 drain_right drain_right.n7 24.8943
R335 drain_right.n3 drain_right.t4 19.8005
R336 drain_right.n3 drain_right.t2 19.8005
R337 drain_right.n4 drain_right.t3 19.8005
R338 drain_right.n4 drain_right.t5 19.8005
R339 drain_right.n5 drain_right.t11 19.8005
R340 drain_right.n5 drain_right.t14 19.8005
R341 drain_right.n1 drain_right.t12 19.8005
R342 drain_right.n1 drain_right.t1 19.8005
R343 drain_right.n0 drain_right.t0 19.8005
R344 drain_right.n0 drain_right.t10 19.8005
R345 drain_right.n8 drain_right.t7 19.8005
R346 drain_right.n8 drain_right.t6 19.8005
R347 drain_right.n9 drain_right.t9 19.8005
R348 drain_right.n9 drain_right.t8 19.8005
R349 drain_right.n11 drain_right.t13 19.8005
R350 drain_right.n11 drain_right.t16 19.8005
R351 drain_right.n13 drain_right.t17 19.8005
R352 drain_right.n13 drain_right.t15 19.8005
R353 drain_right.n15 drain_right.t19 19.8005
R354 drain_right.n15 drain_right.t18 19.8005
R355 drain_right drain_right.n16 6.45494
R356 drain_right.n16 drain_right.n14 0.802224
R357 drain_right.n14 drain_right.n12 0.802224
R358 drain_right.n12 drain_right.n10 0.802224
R359 drain_right.n7 drain_right.n6 0.746878
R360 drain_right.n7 drain_right.n2 0.746878
C0 drain_right plus 0.440483f
C1 drain_right drain_left 1.48725f
C2 drain_right source 5.73711f
C3 plus minus 4.56554f
C4 minus drain_left 0.180909f
C5 minus source 2.29356f
C6 plus drain_left 1.84313f
C7 plus source 2.30743f
C8 source drain_left 5.73529f
C9 drain_right minus 1.56872f
C10 drain_right a_n2762_n1088# 4.58845f
C11 drain_left a_n2762_n1088# 4.93926f
C12 source a_n2762_n1088# 2.855442f
C13 minus a_n2762_n1088# 10.138638f
C14 plus a_n2762_n1088# 11.16678f
C15 drain_right.t0 a_n2762_n1088# 0.016723f
C16 drain_right.t10 a_n2762_n1088# 0.016723f
C17 drain_right.n0 a_n2762_n1088# 0.065864f
C18 drain_right.t12 a_n2762_n1088# 0.016723f
C19 drain_right.t1 a_n2762_n1088# 0.016723f
C20 drain_right.n1 a_n2762_n1088# 0.06498f
C21 drain_right.n2 a_n2762_n1088# 0.519169f
C22 drain_right.t4 a_n2762_n1088# 0.016723f
C23 drain_right.t2 a_n2762_n1088# 0.016723f
C24 drain_right.n3 a_n2762_n1088# 0.06498f
C25 drain_right.t3 a_n2762_n1088# 0.016723f
C26 drain_right.t5 a_n2762_n1088# 0.016723f
C27 drain_right.n4 a_n2762_n1088# 0.065864f
C28 drain_right.t11 a_n2762_n1088# 0.016723f
C29 drain_right.t14 a_n2762_n1088# 0.016723f
C30 drain_right.n5 a_n2762_n1088# 0.06498f
C31 drain_right.n6 a_n2762_n1088# 0.519169f
C32 drain_right.n7 a_n2762_n1088# 0.937496f
C33 drain_right.t7 a_n2762_n1088# 0.016723f
C34 drain_right.t6 a_n2762_n1088# 0.016723f
C35 drain_right.n8 a_n2762_n1088# 0.065864f
C36 drain_right.t9 a_n2762_n1088# 0.016723f
C37 drain_right.t8 a_n2762_n1088# 0.016723f
C38 drain_right.n9 a_n2762_n1088# 0.06498f
C39 drain_right.n10 a_n2762_n1088# 0.522285f
C40 drain_right.t13 a_n2762_n1088# 0.016723f
C41 drain_right.t16 a_n2762_n1088# 0.016723f
C42 drain_right.n11 a_n2762_n1088# 0.06498f
C43 drain_right.n12 a_n2762_n1088# 0.257323f
C44 drain_right.t17 a_n2762_n1088# 0.016723f
C45 drain_right.t15 a_n2762_n1088# 0.016723f
C46 drain_right.n13 a_n2762_n1088# 0.06498f
C47 drain_right.n14 a_n2762_n1088# 0.257323f
C48 drain_right.t19 a_n2762_n1088# 0.016723f
C49 drain_right.t18 a_n2762_n1088# 0.016723f
C50 drain_right.n15 a_n2762_n1088# 0.06498f
C51 drain_right.n16 a_n2762_n1088# 0.441853f
C52 minus.n0 a_n2762_n1088# 0.048734f
C53 minus.n1 a_n2762_n1088# 0.008307f
C54 minus.t2 a_n2762_n1088# 0.074481f
C55 minus.n2 a_n2762_n1088# 0.036607f
C56 minus.n3 a_n2762_n1088# 0.008307f
C57 minus.t6 a_n2762_n1088# 0.074481f
C58 minus.n4 a_n2762_n1088# 0.036607f
C59 minus.n5 a_n2762_n1088# 0.008307f
C60 minus.t10 a_n2762_n1088# 0.074481f
C61 minus.t13 a_n2762_n1088# 0.089853f
C62 minus.n6 a_n2762_n1088# 0.061226f
C63 minus.t12 a_n2762_n1088# 0.074481f
C64 minus.n7 a_n2762_n1088# 0.084119f
C65 minus.t11 a_n2762_n1088# 0.074481f
C66 minus.n8 a_n2762_n1088# 0.076376f
C67 minus.n9 a_n2762_n1088# 0.156251f
C68 minus.n10 a_n2762_n1088# 0.036607f
C69 minus.n11 a_n2762_n1088# 0.036607f
C70 minus.n12 a_n2762_n1088# 0.077392f
C71 minus.n13 a_n2762_n1088# 0.008307f
C72 minus.t3 a_n2762_n1088# 0.074481f
C73 minus.n14 a_n2762_n1088# 0.077392f
C74 minus.n15 a_n2762_n1088# 0.036607f
C75 minus.n16 a_n2762_n1088# 0.036607f
C76 minus.n17 a_n2762_n1088# 0.036607f
C77 minus.n18 a_n2762_n1088# 0.077392f
C78 minus.n19 a_n2762_n1088# 0.008307f
C79 minus.t4 a_n2762_n1088# 0.074481f
C80 minus.n20 a_n2762_n1088# 0.077392f
C81 minus.n21 a_n2762_n1088# 0.036607f
C82 minus.n22 a_n2762_n1088# 0.036607f
C83 minus.n23 a_n2762_n1088# 0.048848f
C84 minus.n24 a_n2762_n1088# 0.076376f
C85 minus.t1 a_n2762_n1088# 0.074481f
C86 minus.n25 a_n2762_n1088# 0.084119f
C87 minus.t0 a_n2762_n1088# 0.074481f
C88 minus.n26 a_n2762_n1088# 0.075812f
C89 minus.n27 a_n2762_n1088# 1.04385f
C90 minus.n28 a_n2762_n1088# 0.048734f
C91 minus.n29 a_n2762_n1088# 0.008307f
C92 minus.n30 a_n2762_n1088# 0.036607f
C93 minus.n31 a_n2762_n1088# 0.008307f
C94 minus.n32 a_n2762_n1088# 0.036607f
C95 minus.n33 a_n2762_n1088# 0.008307f
C96 minus.t19 a_n2762_n1088# 0.089853f
C97 minus.n34 a_n2762_n1088# 0.061226f
C98 minus.t9 a_n2762_n1088# 0.074481f
C99 minus.n35 a_n2762_n1088# 0.084119f
C100 minus.t7 a_n2762_n1088# 0.074481f
C101 minus.n36 a_n2762_n1088# 0.076376f
C102 minus.n37 a_n2762_n1088# 0.156251f
C103 minus.n38 a_n2762_n1088# 0.036607f
C104 minus.n39 a_n2762_n1088# 0.036607f
C105 minus.t18 a_n2762_n1088# 0.074481f
C106 minus.n40 a_n2762_n1088# 0.077392f
C107 minus.n41 a_n2762_n1088# 0.008307f
C108 minus.t15 a_n2762_n1088# 0.074481f
C109 minus.n42 a_n2762_n1088# 0.077392f
C110 minus.n43 a_n2762_n1088# 0.036607f
C111 minus.n44 a_n2762_n1088# 0.036607f
C112 minus.n45 a_n2762_n1088# 0.036607f
C113 minus.t17 a_n2762_n1088# 0.074481f
C114 minus.n46 a_n2762_n1088# 0.077392f
C115 minus.n47 a_n2762_n1088# 0.008307f
C116 minus.t8 a_n2762_n1088# 0.074481f
C117 minus.n48 a_n2762_n1088# 0.077392f
C118 minus.n49 a_n2762_n1088# 0.036607f
C119 minus.n50 a_n2762_n1088# 0.036607f
C120 minus.n51 a_n2762_n1088# 0.048848f
C121 minus.t5 a_n2762_n1088# 0.074481f
C122 minus.n52 a_n2762_n1088# 0.076376f
C123 minus.t16 a_n2762_n1088# 0.074481f
C124 minus.n53 a_n2762_n1088# 0.084119f
C125 minus.t14 a_n2762_n1088# 0.074481f
C126 minus.n54 a_n2762_n1088# 0.075812f
C127 minus.n55 a_n2762_n1088# 0.262653f
C128 minus.n56 a_n2762_n1088# 1.26424f
C129 drain_left.t12 a_n2762_n1088# 0.016483f
C130 drain_left.t5 a_n2762_n1088# 0.016483f
C131 drain_left.n0 a_n2762_n1088# 0.064921f
C132 drain_left.t1 a_n2762_n1088# 0.016483f
C133 drain_left.t18 a_n2762_n1088# 0.016483f
C134 drain_left.n1 a_n2762_n1088# 0.064049f
C135 drain_left.n2 a_n2762_n1088# 0.511737f
C136 drain_left.t11 a_n2762_n1088# 0.016483f
C137 drain_left.t7 a_n2762_n1088# 0.016483f
C138 drain_left.n3 a_n2762_n1088# 0.064049f
C139 drain_left.t15 a_n2762_n1088# 0.016483f
C140 drain_left.t9 a_n2762_n1088# 0.016483f
C141 drain_left.n4 a_n2762_n1088# 0.064921f
C142 drain_left.t2 a_n2762_n1088# 0.016483f
C143 drain_left.t0 a_n2762_n1088# 0.016483f
C144 drain_left.n5 a_n2762_n1088# 0.064049f
C145 drain_left.n6 a_n2762_n1088# 0.511737f
C146 drain_left.n7 a_n2762_n1088# 0.964137f
C147 drain_left.t3 a_n2762_n1088# 0.016483f
C148 drain_left.t4 a_n2762_n1088# 0.016483f
C149 drain_left.n8 a_n2762_n1088# 0.064921f
C150 drain_left.t6 a_n2762_n1088# 0.016483f
C151 drain_left.t8 a_n2762_n1088# 0.016483f
C152 drain_left.n9 a_n2762_n1088# 0.064049f
C153 drain_left.n10 a_n2762_n1088# 0.514809f
C154 drain_left.t10 a_n2762_n1088# 0.016483f
C155 drain_left.t13 a_n2762_n1088# 0.016483f
C156 drain_left.n11 a_n2762_n1088# 0.064049f
C157 drain_left.n12 a_n2762_n1088# 0.25364f
C158 drain_left.t14 a_n2762_n1088# 0.016483f
C159 drain_left.t16 a_n2762_n1088# 0.016483f
C160 drain_left.n13 a_n2762_n1088# 0.064049f
C161 drain_left.n14 a_n2762_n1088# 0.25364f
C162 drain_left.t17 a_n2762_n1088# 0.016483f
C163 drain_left.t19 a_n2762_n1088# 0.016483f
C164 drain_left.n15 a_n2762_n1088# 0.064049f
C165 drain_left.n16 a_n2762_n1088# 0.435528f
C166 source.t32 a_n2762_n1088# 0.159466f
C167 source.n0 a_n2762_n1088# 0.738724f
C168 source.t33 a_n2762_n1088# 0.028651f
C169 source.t31 a_n2762_n1088# 0.028651f
C170 source.n1 a_n2762_n1088# 0.092919f
C171 source.n2 a_n2762_n1088# 0.409998f
C172 source.t19 a_n2762_n1088# 0.028651f
C173 source.t22 a_n2762_n1088# 0.028651f
C174 source.n3 a_n2762_n1088# 0.092919f
C175 source.n4 a_n2762_n1088# 0.409998f
C176 source.t20 a_n2762_n1088# 0.028651f
C177 source.t38 a_n2762_n1088# 0.028651f
C178 source.n5 a_n2762_n1088# 0.092919f
C179 source.n6 a_n2762_n1088# 0.409998f
C180 source.t30 a_n2762_n1088# 0.028651f
C181 source.t27 a_n2762_n1088# 0.028651f
C182 source.n7 a_n2762_n1088# 0.092919f
C183 source.n8 a_n2762_n1088# 0.409998f
C184 source.t37 a_n2762_n1088# 0.159466f
C185 source.n9 a_n2762_n1088# 0.382815f
C186 source.t8 a_n2762_n1088# 0.159466f
C187 source.n10 a_n2762_n1088# 0.382815f
C188 source.t6 a_n2762_n1088# 0.028651f
C189 source.t10 a_n2762_n1088# 0.028651f
C190 source.n11 a_n2762_n1088# 0.092919f
C191 source.n12 a_n2762_n1088# 0.409998f
C192 source.t16 a_n2762_n1088# 0.028651f
C193 source.t0 a_n2762_n1088# 0.028651f
C194 source.n13 a_n2762_n1088# 0.092919f
C195 source.n14 a_n2762_n1088# 0.409998f
C196 source.t14 a_n2762_n1088# 0.028651f
C197 source.t1 a_n2762_n1088# 0.028651f
C198 source.n15 a_n2762_n1088# 0.092919f
C199 source.n16 a_n2762_n1088# 0.409998f
C200 source.t39 a_n2762_n1088# 0.028651f
C201 source.t18 a_n2762_n1088# 0.028651f
C202 source.n17 a_n2762_n1088# 0.092919f
C203 source.n18 a_n2762_n1088# 0.409998f
C204 source.t17 a_n2762_n1088# 0.159466f
C205 source.n19 a_n2762_n1088# 1.03567f
C206 source.t23 a_n2762_n1088# 0.159466f
C207 source.n20 a_n2762_n1088# 1.03567f
C208 source.t21 a_n2762_n1088# 0.028651f
C209 source.t25 a_n2762_n1088# 0.028651f
C210 source.n21 a_n2762_n1088# 0.092919f
C211 source.n22 a_n2762_n1088# 0.409998f
C212 source.t26 a_n2762_n1088# 0.028651f
C213 source.t24 a_n2762_n1088# 0.028651f
C214 source.n23 a_n2762_n1088# 0.092919f
C215 source.n24 a_n2762_n1088# 0.409998f
C216 source.t36 a_n2762_n1088# 0.028651f
C217 source.t34 a_n2762_n1088# 0.028651f
C218 source.n25 a_n2762_n1088# 0.092919f
C219 source.n26 a_n2762_n1088# 0.409998f
C220 source.t35 a_n2762_n1088# 0.028651f
C221 source.t28 a_n2762_n1088# 0.028651f
C222 source.n27 a_n2762_n1088# 0.092919f
C223 source.n28 a_n2762_n1088# 0.409998f
C224 source.t29 a_n2762_n1088# 0.159466f
C225 source.n29 a_n2762_n1088# 0.382816f
C226 source.t13 a_n2762_n1088# 0.159466f
C227 source.n30 a_n2762_n1088# 0.382816f
C228 source.t9 a_n2762_n1088# 0.028651f
C229 source.t7 a_n2762_n1088# 0.028651f
C230 source.n31 a_n2762_n1088# 0.092919f
C231 source.n32 a_n2762_n1088# 0.409998f
C232 source.t12 a_n2762_n1088# 0.028651f
C233 source.t4 a_n2762_n1088# 0.028651f
C234 source.n33 a_n2762_n1088# 0.092919f
C235 source.n34 a_n2762_n1088# 0.409998f
C236 source.t2 a_n2762_n1088# 0.028651f
C237 source.t11 a_n2762_n1088# 0.028651f
C238 source.n35 a_n2762_n1088# 0.092919f
C239 source.n36 a_n2762_n1088# 0.409998f
C240 source.t15 a_n2762_n1088# 0.028651f
C241 source.t3 a_n2762_n1088# 0.028651f
C242 source.n37 a_n2762_n1088# 0.092919f
C243 source.n38 a_n2762_n1088# 0.409998f
C244 source.t5 a_n2762_n1088# 0.159466f
C245 source.n39 a_n2762_n1088# 0.611425f
C246 source.n40 a_n2762_n1088# 0.746984f
C247 plus.n0 a_n2762_n1088# 0.049262f
C248 plus.t0 a_n2762_n1088# 0.075289f
C249 plus.t2 a_n2762_n1088# 0.075289f
C250 plus.t3 a_n2762_n1088# 0.075289f
C251 plus.n1 a_n2762_n1088# 0.049378f
C252 plus.t5 a_n2762_n1088# 0.075289f
C253 plus.n2 a_n2762_n1088# 0.078231f
C254 plus.n3 a_n2762_n1088# 0.037004f
C255 plus.t6 a_n2762_n1088# 0.075289f
C256 plus.t9 a_n2762_n1088# 0.075289f
C257 plus.n4 a_n2762_n1088# 0.078231f
C258 plus.n5 a_n2762_n1088# 0.037004f
C259 plus.t11 a_n2762_n1088# 0.075289f
C260 plus.t13 a_n2762_n1088# 0.075289f
C261 plus.n6 a_n2762_n1088# 0.077204f
C262 plus.t15 a_n2762_n1088# 0.075289f
C263 plus.n7 a_n2762_n1088# 0.085031f
C264 plus.t16 a_n2762_n1088# 0.090827f
C265 plus.n8 a_n2762_n1088# 0.06189f
C266 plus.n9 a_n2762_n1088# 0.157946f
C267 plus.n10 a_n2762_n1088# 0.037004f
C268 plus.n11 a_n2762_n1088# 0.008397f
C269 plus.n12 a_n2762_n1088# 0.078231f
C270 plus.n13 a_n2762_n1088# 0.008397f
C271 plus.n14 a_n2762_n1088# 0.037004f
C272 plus.n15 a_n2762_n1088# 0.037004f
C273 plus.n16 a_n2762_n1088# 0.037004f
C274 plus.n17 a_n2762_n1088# 0.008397f
C275 plus.n18 a_n2762_n1088# 0.078231f
C276 plus.n19 a_n2762_n1088# 0.008397f
C277 plus.n20 a_n2762_n1088# 0.037004f
C278 plus.n21 a_n2762_n1088# 0.037004f
C279 plus.n22 a_n2762_n1088# 0.037004f
C280 plus.n23 a_n2762_n1088# 0.008397f
C281 plus.n24 a_n2762_n1088# 0.077204f
C282 plus.n25 a_n2762_n1088# 0.085031f
C283 plus.n26 a_n2762_n1088# 0.076634f
C284 plus.n27 a_n2762_n1088# 0.277887f
C285 plus.n28 a_n2762_n1088# 0.049262f
C286 plus.t7 a_n2762_n1088# 0.075289f
C287 plus.t14 a_n2762_n1088# 0.075289f
C288 plus.n29 a_n2762_n1088# 0.049378f
C289 plus.t18 a_n2762_n1088# 0.075289f
C290 plus.t1 a_n2762_n1088# 0.075289f
C291 plus.n30 a_n2762_n1088# 0.078231f
C292 plus.n31 a_n2762_n1088# 0.037004f
C293 plus.t8 a_n2762_n1088# 0.075289f
C294 plus.t12 a_n2762_n1088# 0.075289f
C295 plus.n32 a_n2762_n1088# 0.078231f
C296 plus.n33 a_n2762_n1088# 0.037004f
C297 plus.t17 a_n2762_n1088# 0.075289f
C298 plus.t19 a_n2762_n1088# 0.075289f
C299 plus.n34 a_n2762_n1088# 0.077204f
C300 plus.t4 a_n2762_n1088# 0.075289f
C301 plus.n35 a_n2762_n1088# 0.085031f
C302 plus.t10 a_n2762_n1088# 0.090827f
C303 plus.n36 a_n2762_n1088# 0.06189f
C304 plus.n37 a_n2762_n1088# 0.157946f
C305 plus.n38 a_n2762_n1088# 0.037004f
C306 plus.n39 a_n2762_n1088# 0.008397f
C307 plus.n40 a_n2762_n1088# 0.078231f
C308 plus.n41 a_n2762_n1088# 0.008397f
C309 plus.n42 a_n2762_n1088# 0.037004f
C310 plus.n43 a_n2762_n1088# 0.037004f
C311 plus.n44 a_n2762_n1088# 0.037004f
C312 plus.n45 a_n2762_n1088# 0.008397f
C313 plus.n46 a_n2762_n1088# 0.078231f
C314 plus.n47 a_n2762_n1088# 0.008397f
C315 plus.n48 a_n2762_n1088# 0.037004f
C316 plus.n49 a_n2762_n1088# 0.037004f
C317 plus.n50 a_n2762_n1088# 0.037004f
C318 plus.n51 a_n2762_n1088# 0.008397f
C319 plus.n52 a_n2762_n1088# 0.077204f
C320 plus.n53 a_n2762_n1088# 0.085031f
C321 plus.n54 a_n2762_n1088# 0.076634f
C322 plus.n55 a_n2762_n1088# 1.01742f
.ends

