* NGSPICE file created from diffpair215.ext - technology: sky130A

.subckt diffpair215 minus drain_right drain_left source plus
X0 source.t18 minus.t0 drain_right.t1 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X1 drain_left.t11 plus.t0 source.t0 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X2 drain_right.t4 minus.t1 source.t17 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X3 source.t2 plus.t1 drain_left.t10 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X4 a_n2018_n1488# a_n2018_n1488# a_n2018_n1488# a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.6
X5 drain_right.t9 minus.t2 source.t16 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X6 source.t15 minus.t3 drain_right.t7 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X7 drain_left.t9 plus.t2 source.t20 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X8 drain_left.t8 plus.t3 source.t21 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X9 source.t22 plus.t4 drain_left.t7 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X10 source.t14 minus.t4 drain_right.t8 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X11 source.t13 minus.t5 drain_right.t2 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X12 drain_right.t0 minus.t6 source.t12 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X13 source.t23 plus.t5 drain_left.t6 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X14 drain_left.t5 plus.t6 source.t4 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X15 source.t11 minus.t7 drain_right.t3 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X16 a_n2018_n1488# a_n2018_n1488# a_n2018_n1488# a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X17 drain_right.t11 minus.t8 source.t10 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X18 drain_right.t10 minus.t9 source.t9 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X19 source.t3 plus.t7 drain_left.t4 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X20 drain_right.t5 minus.t10 source.t8 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X21 source.t7 minus.t11 drain_right.t6 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X22 a_n2018_n1488# a_n2018_n1488# a_n2018_n1488# a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X23 drain_left.t3 plus.t8 source.t6 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X24 source.t5 plus.t9 drain_left.t2 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X25 drain_left.t1 plus.t10 source.t19 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X26 a_n2018_n1488# a_n2018_n1488# a_n2018_n1488# a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X27 source.t1 plus.t11 drain_left.t0 a_n2018_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
R0 minus.n2 minus.t10 211.031
R1 minus.n14 minus.t11 211.031
R2 minus.n3 minus.t7 185.972
R3 minus.n4 minus.t6 185.972
R4 minus.n1 minus.t4 185.972
R5 minus.n8 minus.t2 185.972
R6 minus.n10 minus.t3 185.972
R7 minus.n15 minus.t1 185.972
R8 minus.n16 minus.t0 185.972
R9 minus.n13 minus.t9 185.972
R10 minus.n20 minus.t5 185.972
R11 minus.n22 minus.t8 185.972
R12 minus.n11 minus.n10 161.3
R13 minus.n9 minus.n0 161.3
R14 minus.n8 minus.n7 161.3
R15 minus.n23 minus.n22 161.3
R16 minus.n21 minus.n12 161.3
R17 minus.n20 minus.n19 161.3
R18 minus.n6 minus.n1 80.6037
R19 minus.n5 minus.n4 80.6037
R20 minus.n18 minus.n13 80.6037
R21 minus.n17 minus.n16 80.6037
R22 minus.n4 minus.n3 48.2005
R23 minus.n4 minus.n1 48.2005
R24 minus.n8 minus.n1 48.2005
R25 minus.n16 minus.n15 48.2005
R26 minus.n16 minus.n13 48.2005
R27 minus.n20 minus.n13 48.2005
R28 minus.n5 minus.n2 45.0744
R29 minus.n17 minus.n14 45.0744
R30 minus.n10 minus.n9 40.1672
R31 minus.n22 minus.n21 40.1672
R32 minus.n24 minus.n11 30.0346
R33 minus.n3 minus.n2 16.1124
R34 minus.n15 minus.n14 16.1124
R35 minus.n9 minus.n8 8.03383
R36 minus.n21 minus.n20 8.03383
R37 minus.n24 minus.n23 6.58762
R38 minus.n6 minus.n5 0.380177
R39 minus.n18 minus.n17 0.380177
R40 minus.n7 minus.n6 0.285035
R41 minus.n19 minus.n18 0.285035
R42 minus.n11 minus.n0 0.189894
R43 minus.n7 minus.n0 0.189894
R44 minus.n19 minus.n12 0.189894
R45 minus.n23 minus.n12 0.189894
R46 minus minus.n24 0.188
R47 drain_right.n6 drain_right.n4 80.5748
R48 drain_right.n3 drain_right.n2 80.5194
R49 drain_right.n3 drain_right.n0 80.5194
R50 drain_right.n6 drain_right.n5 79.7731
R51 drain_right.n8 drain_right.n7 79.7731
R52 drain_right.n3 drain_right.n1 79.773
R53 drain_right drain_right.n3 24.0043
R54 drain_right.n1 drain_right.t1 6.6005
R55 drain_right.n1 drain_right.t10 6.6005
R56 drain_right.n2 drain_right.t2 6.6005
R57 drain_right.n2 drain_right.t11 6.6005
R58 drain_right.n0 drain_right.t6 6.6005
R59 drain_right.n0 drain_right.t4 6.6005
R60 drain_right.n4 drain_right.t3 6.6005
R61 drain_right.n4 drain_right.t5 6.6005
R62 drain_right.n5 drain_right.t8 6.6005
R63 drain_right.n5 drain_right.t0 6.6005
R64 drain_right.n7 drain_right.t7 6.6005
R65 drain_right.n7 drain_right.t9 6.6005
R66 drain_right drain_right.n8 6.45494
R67 drain_right.n8 drain_right.n6 0.802224
R68 source.n0 source.t0 69.6943
R69 source.n5 source.t5 69.6943
R70 source.n6 source.t8 69.6943
R71 source.n11 source.t15 69.6943
R72 source.n23 source.t10 69.6942
R73 source.n18 source.t7 69.6942
R74 source.n17 source.t20 69.6942
R75 source.n12 source.t2 69.6942
R76 source.n2 source.n1 63.0943
R77 source.n4 source.n3 63.0943
R78 source.n8 source.n7 63.0943
R79 source.n10 source.n9 63.0943
R80 source.n22 source.n21 63.0942
R81 source.n20 source.n19 63.0942
R82 source.n16 source.n15 63.0942
R83 source.n14 source.n13 63.0942
R84 source.n12 source.n11 15.2713
R85 source.n24 source.n0 9.60747
R86 source.n21 source.t9 6.6005
R87 source.n21 source.t13 6.6005
R88 source.n19 source.t17 6.6005
R89 source.n19 source.t18 6.6005
R90 source.n15 source.t19 6.6005
R91 source.n15 source.t1 6.6005
R92 source.n13 source.t21 6.6005
R93 source.n13 source.t23 6.6005
R94 source.n1 source.t4 6.6005
R95 source.n1 source.t22 6.6005
R96 source.n3 source.t6 6.6005
R97 source.n3 source.t3 6.6005
R98 source.n7 source.t12 6.6005
R99 source.n7 source.t11 6.6005
R100 source.n9 source.t16 6.6005
R101 source.n9 source.t14 6.6005
R102 source.n24 source.n23 5.66429
R103 source.n11 source.n10 0.802224
R104 source.n10 source.n8 0.802224
R105 source.n8 source.n6 0.802224
R106 source.n5 source.n4 0.802224
R107 source.n4 source.n2 0.802224
R108 source.n2 source.n0 0.802224
R109 source.n14 source.n12 0.802224
R110 source.n16 source.n14 0.802224
R111 source.n17 source.n16 0.802224
R112 source.n20 source.n18 0.802224
R113 source.n22 source.n20 0.802224
R114 source.n23 source.n22 0.802224
R115 source.n6 source.n5 0.470328
R116 source.n18 source.n17 0.470328
R117 source source.n24 0.188
R118 plus.n4 plus.t9 211.031
R119 plus.n16 plus.t2 211.031
R120 plus.n10 plus.t0 185.972
R121 plus.n8 plus.t4 185.972
R122 plus.n7 plus.t6 185.972
R123 plus.n6 plus.t7 185.972
R124 plus.n5 plus.t8 185.972
R125 plus.n22 plus.t1 185.972
R126 plus.n20 plus.t3 185.972
R127 plus.n19 plus.t5 185.972
R128 plus.n18 plus.t10 185.972
R129 plus.n17 plus.t11 185.972
R130 plus.n8 plus.n1 161.3
R131 plus.n9 plus.n0 161.3
R132 plus.n11 plus.n10 161.3
R133 plus.n20 plus.n13 161.3
R134 plus.n21 plus.n12 161.3
R135 plus.n23 plus.n22 161.3
R136 plus.n6 plus.n3 80.6037
R137 plus.n7 plus.n2 80.6037
R138 plus.n18 plus.n15 80.6037
R139 plus.n19 plus.n14 80.6037
R140 plus.n8 plus.n7 48.2005
R141 plus.n7 plus.n6 48.2005
R142 plus.n6 plus.n5 48.2005
R143 plus.n20 plus.n19 48.2005
R144 plus.n19 plus.n18 48.2005
R145 plus.n18 plus.n17 48.2005
R146 plus.n4 plus.n3 45.0744
R147 plus.n16 plus.n15 45.0744
R148 plus.n10 plus.n9 40.1672
R149 plus.n22 plus.n21 40.1672
R150 plus plus.n23 27.3248
R151 plus.n5 plus.n4 16.1124
R152 plus.n17 plus.n16 16.1124
R153 plus plus.n11 8.82247
R154 plus.n9 plus.n8 8.03383
R155 plus.n21 plus.n20 8.03383
R156 plus.n3 plus.n2 0.380177
R157 plus.n15 plus.n14 0.380177
R158 plus.n2 plus.n1 0.285035
R159 plus.n14 plus.n13 0.285035
R160 plus.n1 plus.n0 0.189894
R161 plus.n11 plus.n0 0.189894
R162 plus.n23 plus.n12 0.189894
R163 plus.n13 plus.n12 0.189894
R164 drain_left.n6 drain_left.n4 80.5748
R165 drain_left.n3 drain_left.n2 80.5194
R166 drain_left.n3 drain_left.n0 80.5194
R167 drain_left.n8 drain_left.n7 79.7731
R168 drain_left.n6 drain_left.n5 79.7731
R169 drain_left.n3 drain_left.n1 79.773
R170 drain_left drain_left.n3 24.5575
R171 drain_left.n1 drain_left.t6 6.6005
R172 drain_left.n1 drain_left.t1 6.6005
R173 drain_left.n2 drain_left.t0 6.6005
R174 drain_left.n2 drain_left.t9 6.6005
R175 drain_left.n0 drain_left.t10 6.6005
R176 drain_left.n0 drain_left.t8 6.6005
R177 drain_left.n7 drain_left.t7 6.6005
R178 drain_left.n7 drain_left.t11 6.6005
R179 drain_left.n5 drain_left.t4 6.6005
R180 drain_left.n5 drain_left.t5 6.6005
R181 drain_left.n4 drain_left.t2 6.6005
R182 drain_left.n4 drain_left.t3 6.6005
R183 drain_left drain_left.n8 6.45494
R184 drain_left.n8 drain_left.n6 0.802224
C0 minus drain_right 2.1622f
C1 source drain_left 6.18609f
C2 plus drain_right 0.357897f
C3 drain_left drain_right 1.01255f
C4 source drain_right 6.1876f
C5 minus plus 4.00395f
C6 minus drain_left 0.177012f
C7 minus source 2.45573f
C8 plus drain_left 2.35931f
C9 source plus 2.46972f
C10 drain_right a_n2018_n1488# 4.31909f
C11 drain_left a_n2018_n1488# 4.62492f
C12 source a_n2018_n1488# 3.764227f
C13 minus a_n2018_n1488# 7.205065f
C14 plus a_n2018_n1488# 8.50001f
C15 drain_left.t10 a_n2018_n1488# 0.065271f
C16 drain_left.t8 a_n2018_n1488# 0.065271f
C17 drain_left.n0 a_n2018_n1488# 0.474151f
C18 drain_left.t6 a_n2018_n1488# 0.065271f
C19 drain_left.t1 a_n2018_n1488# 0.065271f
C20 drain_left.n1 a_n2018_n1488# 0.470725f
C21 drain_left.t0 a_n2018_n1488# 0.065271f
C22 drain_left.t9 a_n2018_n1488# 0.065271f
C23 drain_left.n2 a_n2018_n1488# 0.474151f
C24 drain_left.n3 a_n2018_n1488# 1.92592f
C25 drain_left.t2 a_n2018_n1488# 0.065271f
C26 drain_left.t3 a_n2018_n1488# 0.065271f
C27 drain_left.n4 a_n2018_n1488# 0.474446f
C28 drain_left.t4 a_n2018_n1488# 0.065271f
C29 drain_left.t5 a_n2018_n1488# 0.065271f
C30 drain_left.n5 a_n2018_n1488# 0.470727f
C31 drain_left.n6 a_n2018_n1488# 0.73265f
C32 drain_left.t7 a_n2018_n1488# 0.065271f
C33 drain_left.t11 a_n2018_n1488# 0.065271f
C34 drain_left.n7 a_n2018_n1488# 0.470727f
C35 drain_left.n8 a_n2018_n1488# 0.602719f
C36 plus.n0 a_n2018_n1488# 0.047625f
C37 plus.t0 a_n2018_n1488# 0.257061f
C38 plus.t4 a_n2018_n1488# 0.257061f
C39 plus.n1 a_n2018_n1488# 0.06355f
C40 plus.t6 a_n2018_n1488# 0.257061f
C41 plus.n2 a_n2018_n1488# 0.079326f
C42 plus.t7 a_n2018_n1488# 0.257061f
C43 plus.n3 a_n2018_n1488# 0.244087f
C44 plus.t8 a_n2018_n1488# 0.257061f
C45 plus.t9 a_n2018_n1488# 0.275052f
C46 plus.n4 a_n2018_n1488# 0.137146f
C47 plus.n5 a_n2018_n1488# 0.161085f
C48 plus.n6 a_n2018_n1488# 0.162824f
C49 plus.n7 a_n2018_n1488# 0.162824f
C50 plus.n8 a_n2018_n1488# 0.153632f
C51 plus.n9 a_n2018_n1488# 0.010807f
C52 plus.n10 a_n2018_n1488# 0.150402f
C53 plus.n11 a_n2018_n1488# 0.366068f
C54 plus.n12 a_n2018_n1488# 0.047625f
C55 plus.t1 a_n2018_n1488# 0.257061f
C56 plus.n13 a_n2018_n1488# 0.06355f
C57 plus.t3 a_n2018_n1488# 0.257061f
C58 plus.n14 a_n2018_n1488# 0.079326f
C59 plus.t5 a_n2018_n1488# 0.257061f
C60 plus.n15 a_n2018_n1488# 0.244087f
C61 plus.t10 a_n2018_n1488# 0.257061f
C62 plus.t2 a_n2018_n1488# 0.275052f
C63 plus.n16 a_n2018_n1488# 0.137146f
C64 plus.t11 a_n2018_n1488# 0.257061f
C65 plus.n17 a_n2018_n1488# 0.161085f
C66 plus.n18 a_n2018_n1488# 0.162824f
C67 plus.n19 a_n2018_n1488# 0.162824f
C68 plus.n20 a_n2018_n1488# 0.153632f
C69 plus.n21 a_n2018_n1488# 0.010807f
C70 plus.n22 a_n2018_n1488# 0.150402f
C71 plus.n23 a_n2018_n1488# 1.17073f
C72 source.t0 a_n2018_n1488# 0.532412f
C73 source.n0 a_n2018_n1488# 0.766003f
C74 source.t4 a_n2018_n1488# 0.064117f
C75 source.t22 a_n2018_n1488# 0.064117f
C76 source.n1 a_n2018_n1488# 0.406535f
C77 source.n2 a_n2018_n1488# 0.375336f
C78 source.t6 a_n2018_n1488# 0.064117f
C79 source.t3 a_n2018_n1488# 0.064117f
C80 source.n3 a_n2018_n1488# 0.406535f
C81 source.n4 a_n2018_n1488# 0.375336f
C82 source.t5 a_n2018_n1488# 0.532412f
C83 source.n5 a_n2018_n1488# 0.395399f
C84 source.t8 a_n2018_n1488# 0.532412f
C85 source.n6 a_n2018_n1488# 0.395399f
C86 source.t12 a_n2018_n1488# 0.064117f
C87 source.t11 a_n2018_n1488# 0.064117f
C88 source.n7 a_n2018_n1488# 0.406535f
C89 source.n8 a_n2018_n1488# 0.375336f
C90 source.t16 a_n2018_n1488# 0.064117f
C91 source.t14 a_n2018_n1488# 0.064117f
C92 source.n9 a_n2018_n1488# 0.406535f
C93 source.n10 a_n2018_n1488# 0.375336f
C94 source.t15 a_n2018_n1488# 0.532412f
C95 source.n11 a_n2018_n1488# 1.05338f
C96 source.t2 a_n2018_n1488# 0.532409f
C97 source.n12 a_n2018_n1488# 1.05338f
C98 source.t21 a_n2018_n1488# 0.064117f
C99 source.t23 a_n2018_n1488# 0.064117f
C100 source.n13 a_n2018_n1488# 0.406532f
C101 source.n14 a_n2018_n1488# 0.375339f
C102 source.t19 a_n2018_n1488# 0.064117f
C103 source.t1 a_n2018_n1488# 0.064117f
C104 source.n15 a_n2018_n1488# 0.406532f
C105 source.n16 a_n2018_n1488# 0.375339f
C106 source.t20 a_n2018_n1488# 0.532409f
C107 source.n17 a_n2018_n1488# 0.395402f
C108 source.t7 a_n2018_n1488# 0.532409f
C109 source.n18 a_n2018_n1488# 0.395402f
C110 source.t17 a_n2018_n1488# 0.064117f
C111 source.t18 a_n2018_n1488# 0.064117f
C112 source.n19 a_n2018_n1488# 0.406532f
C113 source.n20 a_n2018_n1488# 0.375339f
C114 source.t9 a_n2018_n1488# 0.064117f
C115 source.t13 a_n2018_n1488# 0.064117f
C116 source.n21 a_n2018_n1488# 0.406532f
C117 source.n22 a_n2018_n1488# 0.375339f
C118 source.t10 a_n2018_n1488# 0.532409f
C119 source.n23 a_n2018_n1488# 0.565934f
C120 source.n24 a_n2018_n1488# 0.794057f
C121 drain_right.t6 a_n2018_n1488# 0.064561f
C122 drain_right.t4 a_n2018_n1488# 0.064561f
C123 drain_right.n0 a_n2018_n1488# 0.468998f
C124 drain_right.t1 a_n2018_n1488# 0.064561f
C125 drain_right.t10 a_n2018_n1488# 0.064561f
C126 drain_right.n1 a_n2018_n1488# 0.465609f
C127 drain_right.t2 a_n2018_n1488# 0.064561f
C128 drain_right.t11 a_n2018_n1488# 0.064561f
C129 drain_right.n2 a_n2018_n1488# 0.468998f
C130 drain_right.n3 a_n2018_n1488# 1.85114f
C131 drain_right.t3 a_n2018_n1488# 0.064561f
C132 drain_right.t5 a_n2018_n1488# 0.064561f
C133 drain_right.n4 a_n2018_n1488# 0.469289f
C134 drain_right.t8 a_n2018_n1488# 0.064561f
C135 drain_right.t0 a_n2018_n1488# 0.064561f
C136 drain_right.n5 a_n2018_n1488# 0.465611f
C137 drain_right.n6 a_n2018_n1488# 0.724688f
C138 drain_right.t7 a_n2018_n1488# 0.064561f
C139 drain_right.t9 a_n2018_n1488# 0.064561f
C140 drain_right.n7 a_n2018_n1488# 0.465611f
C141 drain_right.n8 a_n2018_n1488# 0.596169f
C142 minus.n0 a_n2018_n1488# 0.046057f
C143 minus.t4 a_n2018_n1488# 0.248594f
C144 minus.n1 a_n2018_n1488# 0.157461f
C145 minus.t2 a_n2018_n1488# 0.248594f
C146 minus.t10 a_n2018_n1488# 0.265993f
C147 minus.n2 a_n2018_n1488# 0.132629f
C148 minus.t7 a_n2018_n1488# 0.248594f
C149 minus.n3 a_n2018_n1488# 0.15578f
C150 minus.t6 a_n2018_n1488# 0.248594f
C151 minus.n4 a_n2018_n1488# 0.157461f
C152 minus.n5 a_n2018_n1488# 0.236047f
C153 minus.n6 a_n2018_n1488# 0.076713f
C154 minus.n7 a_n2018_n1488# 0.061457f
C155 minus.n8 a_n2018_n1488# 0.148572f
C156 minus.n9 a_n2018_n1488# 0.010451f
C157 minus.t3 a_n2018_n1488# 0.248594f
C158 minus.n10 a_n2018_n1488# 0.145448f
C159 minus.n11 a_n2018_n1488# 1.20424f
C160 minus.n12 a_n2018_n1488# 0.046057f
C161 minus.t9 a_n2018_n1488# 0.248594f
C162 minus.n13 a_n2018_n1488# 0.157461f
C163 minus.t11 a_n2018_n1488# 0.265993f
C164 minus.n14 a_n2018_n1488# 0.132629f
C165 minus.t1 a_n2018_n1488# 0.248594f
C166 minus.n15 a_n2018_n1488# 0.15578f
C167 minus.t0 a_n2018_n1488# 0.248594f
C168 minus.n16 a_n2018_n1488# 0.157461f
C169 minus.n17 a_n2018_n1488# 0.236047f
C170 minus.n18 a_n2018_n1488# 0.076713f
C171 minus.n19 a_n2018_n1488# 0.061457f
C172 minus.t5 a_n2018_n1488# 0.248594f
C173 minus.n20 a_n2018_n1488# 0.148572f
C174 minus.n21 a_n2018_n1488# 0.010451f
C175 minus.t8 a_n2018_n1488# 0.248594f
C176 minus.n22 a_n2018_n1488# 0.145448f
C177 minus.n23 a_n2018_n1488# 0.310576f
C178 minus.n24 a_n2018_n1488# 1.48086f
.ends

