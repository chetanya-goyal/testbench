* NGSPICE file created from diffpair361.ext - technology: sky130A

.subckt diffpair361 minus drain_right drain_left source plus
X0 a_n1214_n2688# a_n1214_n2688# a_n1214_n2688# a_n1214_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.5
X1 source.t7 minus.t0 drain_right.t2 a_n1214_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X2 source.t0 plus.t0 drain_left.t3 a_n1214_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X3 a_n1214_n2688# a_n1214_n2688# a_n1214_n2688# a_n1214_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X4 a_n1214_n2688# a_n1214_n2688# a_n1214_n2688# a_n1214_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X5 drain_right.t3 minus.t1 source.t6 a_n1214_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X6 drain_left.t2 plus.t1 source.t2 a_n1214_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X7 drain_left.t1 plus.t2 source.t1 a_n1214_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X8 source.t3 plus.t3 drain_left.t0 a_n1214_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X9 a_n1214_n2688# a_n1214_n2688# a_n1214_n2688# a_n1214_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X10 drain_right.t0 minus.t2 source.t5 a_n1214_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X11 source.t4 minus.t3 drain_right.t1 a_n1214_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
R0 minus.n0 minus.t1 533.348
R1 minus.n1 minus.t3 533.348
R2 minus.n0 minus.t0 533.323
R3 minus.n1 minus.t2 533.323
R4 minus.n2 minus.n0 101.725
R5 minus.n2 minus.n1 76.7783
R6 minus minus.n2 0.188
R7 drain_right drain_right.n0 91.509
R8 drain_right drain_right.n1 71.9057
R9 drain_right.n0 drain_right.t1 2.2005
R10 drain_right.n0 drain_right.t0 2.2005
R11 drain_right.n1 drain_right.t2 2.2005
R12 drain_right.n1 drain_right.t3 2.2005
R13 source.n1 source.t0 51.0588
R14 source.n2 source.t6 51.0588
R15 source.n3 source.t7 51.0588
R16 source.n7 source.t5 51.0586
R17 source.n6 source.t4 51.0586
R18 source.n5 source.t1 51.0586
R19 source.n4 source.t3 51.0586
R20 source.n0 source.t2 51.0586
R21 source.n4 source.n3 19.7305
R22 source.n8 source.n0 14.1098
R23 source.n8 source.n7 5.62119
R24 source.n3 source.n2 0.716017
R25 source.n1 source.n0 0.716017
R26 source.n5 source.n4 0.716017
R27 source.n7 source.n6 0.716017
R28 source.n2 source.n1 0.470328
R29 source.n6 source.n5 0.470328
R30 source source.n8 0.188
R31 plus.n0 plus.t0 533.348
R32 plus.n1 plus.t2 533.348
R33 plus.n0 plus.t1 533.323
R34 plus.n1 plus.t3 533.323
R35 plus plus.n1 96.7427
R36 plus plus.n0 81.2859
R37 drain_left drain_left.n0 92.0622
R38 drain_left drain_left.n1 71.9057
R39 drain_left.n0 drain_left.t0 2.2005
R40 drain_left.n0 drain_left.t1 2.2005
R41 drain_left.n1 drain_left.t3 2.2005
R42 drain_left.n1 drain_left.t2 2.2005
C0 plus source 1.78542f
C1 plus minus 4.10281f
C2 drain_left drain_right 0.522435f
C3 drain_left source 6.24636f
C4 drain_left minus 0.170454f
C5 source drain_right 6.24611f
C6 minus drain_right 2.09591f
C7 source minus 1.77138f
C8 plus drain_left 2.20936f
C9 plus drain_right 0.266739f
C10 drain_right a_n1214_n2688# 5.85051f
C11 drain_left a_n1214_n2688# 6.0555f
C12 source a_n1214_n2688# 6.984302f
C13 minus a_n1214_n2688# 4.373488f
C14 plus a_n1214_n2688# 6.92813f
C15 drain_left.t0 a_n1214_n2688# 0.203894f
C16 drain_left.t1 a_n1214_n2688# 0.203894f
C17 drain_left.n0 a_n1214_n2688# 2.10268f
C18 drain_left.t3 a_n1214_n2688# 0.203894f
C19 drain_left.t2 a_n1214_n2688# 0.203894f
C20 drain_left.n1 a_n1214_n2688# 1.83827f
C21 plus.t1 a_n1214_n2688# 0.57231f
C22 plus.t0 a_n1214_n2688# 0.572323f
C23 plus.n0 a_n1214_n2688# 0.527426f
C24 plus.t3 a_n1214_n2688# 0.57231f
C25 plus.t2 a_n1214_n2688# 0.572323f
C26 plus.n1 a_n1214_n2688# 0.770544f
C27 source.t2 a_n1214_n2688# 1.03222f
C28 source.n0 a_n1214_n2688# 0.606208f
C29 source.t0 a_n1214_n2688# 1.03223f
C30 source.n1 a_n1214_n2688# 0.220959f
C31 source.t6 a_n1214_n2688# 1.03223f
C32 source.n2 a_n1214_n2688# 0.220959f
C33 source.t7 a_n1214_n2688# 1.03223f
C34 source.n3 a_n1214_n2688# 0.80644f
C35 source.t3 a_n1214_n2688# 1.03222f
C36 source.n4 a_n1214_n2688# 0.806443f
C37 source.t1 a_n1214_n2688# 1.03222f
C38 source.n5 a_n1214_n2688# 0.220962f
C39 source.t4 a_n1214_n2688# 1.03222f
C40 source.n6 a_n1214_n2688# 0.220962f
C41 source.t5 a_n1214_n2688# 1.03222f
C42 source.n7 a_n1214_n2688# 0.303803f
C43 source.n8 a_n1214_n2688# 0.712555f
C44 drain_right.t1 a_n1214_n2688# 0.204193f
C45 drain_right.t0 a_n1214_n2688# 0.204193f
C46 drain_right.n0 a_n1214_n2688# 2.084f
C47 drain_right.t2 a_n1214_n2688# 0.204193f
C48 drain_right.t3 a_n1214_n2688# 0.204193f
C49 drain_right.n1 a_n1214_n2688# 1.84097f
C50 minus.t1 a_n1214_n2688# 0.555461f
C51 minus.t0 a_n1214_n2688# 0.555449f
C52 minus.n0 a_n1214_n2688# 0.834546f
C53 minus.t3 a_n1214_n2688# 0.555461f
C54 minus.t2 a_n1214_n2688# 0.555449f
C55 minus.n1 a_n1214_n2688# 0.475975f
C56 minus.n2 a_n1214_n2688# 2.63986f
.ends

