* NGSPICE file created from diffpair405.ext - technology: sky130A

.subckt diffpair405 minus drain_right drain_left source plus
X0 a_n1626_n3288# a_n1626_n3288# a_n1626_n3288# a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=45.6 ps=199.6 w=12 l=0.15
X1 source.t23 minus.t0 drain_right.t5 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X2 source.t3 plus.t0 drain_left.t11 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X3 drain_left.t10 plus.t1 source.t7 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X4 a_n1626_n3288# a_n1626_n3288# a_n1626_n3288# a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X5 a_n1626_n3288# a_n1626_n3288# a_n1626_n3288# a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X6 source.t4 plus.t2 drain_left.t9 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X7 source.t22 minus.t1 drain_right.t11 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X8 drain_left.t8 plus.t3 source.t6 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X9 source.t21 minus.t2 drain_right.t4 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X10 drain_left.t7 plus.t4 source.t8 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X11 drain_right.t9 minus.t3 source.t20 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X12 drain_right.t1 minus.t4 source.t19 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X13 drain_right.t7 minus.t5 source.t18 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X14 source.t17 minus.t6 drain_right.t10 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X15 drain_right.t8 minus.t7 source.t16 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X16 source.t0 plus.t5 drain_left.t6 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X17 source.t10 plus.t6 drain_left.t5 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X18 drain_right.t6 minus.t8 source.t15 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X19 a_n1626_n3288# a_n1626_n3288# a_n1626_n3288# a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=0 ps=0 w=12 l=0.15
X20 drain_left.t4 plus.t7 source.t1 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X21 source.t14 minus.t9 drain_right.t3 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=5.7 pd=24.95 as=3 ps=12.5 w=12 l=0.15
X22 source.t13 minus.t10 drain_right.t2 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X23 source.t5 plus.t8 drain_left.t3 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X24 drain_left.t2 plus.t9 source.t2 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=5.7 ps=24.95 w=12 l=0.15
X25 drain_left.t1 plus.t10 source.t9 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X26 source.t11 plus.t11 drain_left.t0 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
X27 drain_right.t0 minus.t11 source.t12 a_n1626_n3288# sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=3 ps=12.5 w=12 l=0.15
R0 minus.n13 minus.t9 2191.64
R1 minus.n2 minus.t3 2191.64
R2 minus.n28 minus.t7 2191.64
R3 minus.n17 minus.t0 2191.64
R4 minus.n12 minus.t4 2136.87
R5 minus.n10 minus.t6 2136.87
R6 minus.n3 minus.t8 2136.87
R7 minus.n4 minus.t2 2136.87
R8 minus.n27 minus.t1 2136.87
R9 minus.n25 minus.t11 2136.87
R10 minus.n19 minus.t10 2136.87
R11 minus.n18 minus.t5 2136.87
R12 minus.n6 minus.n2 161.489
R13 minus.n21 minus.n17 161.489
R14 minus.n14 minus.n13 161.3
R15 minus.n11 minus.n0 161.3
R16 minus.n9 minus.n8 161.3
R17 minus.n7 minus.n1 161.3
R18 minus.n6 minus.n5 161.3
R19 minus.n29 minus.n28 161.3
R20 minus.n26 minus.n15 161.3
R21 minus.n24 minus.n23 161.3
R22 minus.n22 minus.n16 161.3
R23 minus.n21 minus.n20 161.3
R24 minus.n9 minus.n1 73.0308
R25 minus.n24 minus.n16 73.0308
R26 minus.n11 minus.n10 62.0763
R27 minus.n5 minus.n3 62.0763
R28 minus.n20 minus.n19 62.0763
R29 minus.n26 minus.n25 62.0763
R30 minus.n13 minus.n12 40.1672
R31 minus.n4 minus.n2 40.1672
R32 minus.n18 minus.n17 40.1672
R33 minus.n28 minus.n27 40.1672
R34 minus.n30 minus.n14 35.3225
R35 minus.n12 minus.n11 32.8641
R36 minus.n5 minus.n4 32.8641
R37 minus.n20 minus.n18 32.8641
R38 minus.n27 minus.n26 32.8641
R39 minus.n10 minus.n9 10.955
R40 minus.n3 minus.n1 10.955
R41 minus.n19 minus.n16 10.955
R42 minus.n25 minus.n24 10.955
R43 minus.n30 minus.n29 6.54217
R44 minus.n14 minus.n0 0.189894
R45 minus.n8 minus.n0 0.189894
R46 minus.n8 minus.n7 0.189894
R47 minus.n7 minus.n6 0.189894
R48 minus.n22 minus.n21 0.189894
R49 minus.n23 minus.n22 0.189894
R50 minus.n23 minus.n15 0.189894
R51 minus.n29 minus.n15 0.189894
R52 minus minus.n30 0.188
R53 drain_right.n6 drain_right.n4 60.1128
R54 drain_right.n3 drain_right.n2 60.0575
R55 drain_right.n3 drain_right.n0 60.0575
R56 drain_right.n6 drain_right.n5 59.5527
R57 drain_right.n8 drain_right.n7 59.5527
R58 drain_right.n3 drain_right.n1 59.5525
R59 drain_right drain_right.n3 29.6156
R60 drain_right drain_right.n8 6.21356
R61 drain_right.n1 drain_right.t2 2.5005
R62 drain_right.n1 drain_right.t0 2.5005
R63 drain_right.n2 drain_right.t11 2.5005
R64 drain_right.n2 drain_right.t8 2.5005
R65 drain_right.n0 drain_right.t5 2.5005
R66 drain_right.n0 drain_right.t7 2.5005
R67 drain_right.n4 drain_right.t4 2.5005
R68 drain_right.n4 drain_right.t9 2.5005
R69 drain_right.n5 drain_right.t10 2.5005
R70 drain_right.n5 drain_right.t6 2.5005
R71 drain_right.n7 drain_right.t3 2.5005
R72 drain_right.n7 drain_right.t1 2.5005
R73 drain_right.n8 drain_right.n6 0.560845
R74 source.n5 source.t10 45.3739
R75 source.n6 source.t20 45.3739
R76 source.n11 source.t14 45.3739
R77 source.n23 source.t16 45.3737
R78 source.n18 source.t23 45.3737
R79 source.n17 source.t6 45.3737
R80 source.n12 source.t3 45.3737
R81 source.n0 source.t2 45.3737
R82 source.n2 source.n1 42.8739
R83 source.n4 source.n3 42.8739
R84 source.n8 source.n7 42.8739
R85 source.n10 source.n9 42.8739
R86 source.n22 source.n21 42.8737
R87 source.n20 source.n19 42.8737
R88 source.n16 source.n15 42.8737
R89 source.n14 source.n13 42.8737
R90 source.n12 source.n11 21.8481
R91 source.n24 source.n0 16.305
R92 source.n24 source.n23 5.5436
R93 source.n21 source.t12 2.5005
R94 source.n21 source.t22 2.5005
R95 source.n19 source.t18 2.5005
R96 source.n19 source.t13 2.5005
R97 source.n15 source.t7 2.5005
R98 source.n15 source.t0 2.5005
R99 source.n13 source.t8 2.5005
R100 source.n13 source.t4 2.5005
R101 source.n1 source.t1 2.5005
R102 source.n1 source.t11 2.5005
R103 source.n3 source.t9 2.5005
R104 source.n3 source.t5 2.5005
R105 source.n7 source.t15 2.5005
R106 source.n7 source.t21 2.5005
R107 source.n9 source.t19 2.5005
R108 source.n9 source.t17 2.5005
R109 source.n11 source.n10 0.560845
R110 source.n10 source.n8 0.560845
R111 source.n8 source.n6 0.560845
R112 source.n5 source.n4 0.560845
R113 source.n4 source.n2 0.560845
R114 source.n2 source.n0 0.560845
R115 source.n14 source.n12 0.560845
R116 source.n16 source.n14 0.560845
R117 source.n17 source.n16 0.560845
R118 source.n20 source.n18 0.560845
R119 source.n22 source.n20 0.560845
R120 source.n23 source.n22 0.560845
R121 source.n6 source.n5 0.470328
R122 source.n18 source.n17 0.470328
R123 source source.n24 0.188
R124 plus.n2 plus.t6 2191.64
R125 plus.n13 plus.t9 2191.64
R126 plus.n17 plus.t3 2191.64
R127 plus.n28 plus.t0 2191.64
R128 plus.n3 plus.t10 2136.87
R129 plus.n4 plus.t8 2136.87
R130 plus.n10 plus.t7 2136.87
R131 plus.n12 plus.t11 2136.87
R132 plus.n19 plus.t5 2136.87
R133 plus.n18 plus.t1 2136.87
R134 plus.n25 plus.t2 2136.87
R135 plus.n27 plus.t4 2136.87
R136 plus.n6 plus.n2 161.489
R137 plus.n21 plus.n17 161.489
R138 plus.n6 plus.n5 161.3
R139 plus.n7 plus.n1 161.3
R140 plus.n9 plus.n8 161.3
R141 plus.n11 plus.n0 161.3
R142 plus.n14 plus.n13 161.3
R143 plus.n21 plus.n20 161.3
R144 plus.n22 plus.n16 161.3
R145 plus.n24 plus.n23 161.3
R146 plus.n26 plus.n15 161.3
R147 plus.n29 plus.n28 161.3
R148 plus.n9 plus.n1 73.0308
R149 plus.n24 plus.n16 73.0308
R150 plus.n5 plus.n4 62.0763
R151 plus.n11 plus.n10 62.0763
R152 plus.n26 plus.n25 62.0763
R153 plus.n20 plus.n18 62.0763
R154 plus.n3 plus.n2 40.1672
R155 plus.n13 plus.n12 40.1672
R156 plus.n28 plus.n27 40.1672
R157 plus.n19 plus.n17 40.1672
R158 plus.n5 plus.n3 32.8641
R159 plus.n12 plus.n11 32.8641
R160 plus.n27 plus.n26 32.8641
R161 plus.n20 plus.n19 32.8641
R162 plus plus.n29 29.2036
R163 plus plus.n14 12.1861
R164 plus.n4 plus.n1 10.955
R165 plus.n10 plus.n9 10.955
R166 plus.n25 plus.n24 10.955
R167 plus.n18 plus.n16 10.955
R168 plus.n7 plus.n6 0.189894
R169 plus.n8 plus.n7 0.189894
R170 plus.n8 plus.n0 0.189894
R171 plus.n14 plus.n0 0.189894
R172 plus.n29 plus.n15 0.189894
R173 plus.n23 plus.n15 0.189894
R174 plus.n23 plus.n22 0.189894
R175 plus.n22 plus.n21 0.189894
R176 drain_left.n6 drain_left.n4 60.113
R177 drain_left.n3 drain_left.n2 60.0575
R178 drain_left.n3 drain_left.n0 60.0575
R179 drain_left.n6 drain_left.n5 59.5527
R180 drain_left.n3 drain_left.n1 59.5525
R181 drain_left.n8 drain_left.n7 59.5525
R182 drain_left drain_left.n3 30.1688
R183 drain_left drain_left.n8 6.21356
R184 drain_left.n1 drain_left.t9 2.5005
R185 drain_left.n1 drain_left.t10 2.5005
R186 drain_left.n2 drain_left.t6 2.5005
R187 drain_left.n2 drain_left.t8 2.5005
R188 drain_left.n0 drain_left.t11 2.5005
R189 drain_left.n0 drain_left.t7 2.5005
R190 drain_left.n7 drain_left.t0 2.5005
R191 drain_left.n7 drain_left.t2 2.5005
R192 drain_left.n5 drain_left.t3 2.5005
R193 drain_left.n5 drain_left.t4 2.5005
R194 drain_left.n4 drain_left.t5 2.5005
R195 drain_left.n4 drain_left.t1 2.5005
R196 drain_left.n8 drain_left.n6 0.560845
C0 plus drain_left 3.01925f
C1 minus drain_right 2.86276f
C2 plus drain_right 0.309819f
C3 source drain_left 24.016802f
C4 minus plus 5.16374f
C5 source drain_right 24.016699f
C6 source minus 2.33202f
C7 source plus 2.34606f
C8 drain_right drain_left 0.801529f
C9 minus drain_left 0.170585f
C10 drain_right a_n1626_n3288# 5.698009f
C11 drain_left a_n1626_n3288# 5.94005f
C12 source a_n1626_n3288# 8.68202f
C13 minus a_n1626_n3288# 5.980671f
C14 plus a_n1626_n3288# 8.13156f
C15 drain_left.t11 a_n1626_n3288# 0.4041f
C16 drain_left.t7 a_n1626_n3288# 0.4041f
C17 drain_left.n0 a_n1626_n3288# 2.65096f
C18 drain_left.t9 a_n1626_n3288# 0.4041f
C19 drain_left.t10 a_n1626_n3288# 0.4041f
C20 drain_left.n1 a_n1626_n3288# 2.64806f
C21 drain_left.t6 a_n1626_n3288# 0.4041f
C22 drain_left.t8 a_n1626_n3288# 0.4041f
C23 drain_left.n2 a_n1626_n3288# 2.65096f
C24 drain_left.n3 a_n1626_n3288# 2.2892f
C25 drain_left.t5 a_n1626_n3288# 0.4041f
C26 drain_left.t1 a_n1626_n3288# 0.4041f
C27 drain_left.n4 a_n1626_n3288# 2.65132f
C28 drain_left.t3 a_n1626_n3288# 0.4041f
C29 drain_left.t4 a_n1626_n3288# 0.4041f
C30 drain_left.n5 a_n1626_n3288# 2.64807f
C31 drain_left.n6 a_n1626_n3288# 0.68327f
C32 drain_left.t0 a_n1626_n3288# 0.4041f
C33 drain_left.t2 a_n1626_n3288# 0.4041f
C34 drain_left.n7 a_n1626_n3288# 2.64806f
C35 drain_left.n8 a_n1626_n3288# 0.572483f
C36 plus.n0 a_n1626_n3288# 0.057282f
C37 plus.t11 a_n1626_n3288# 0.291362f
C38 plus.t7 a_n1626_n3288# 0.291362f
C39 plus.n1 a_n1626_n3288# 0.021651f
C40 plus.t6 a_n1626_n3288# 0.294494f
C41 plus.n2 a_n1626_n3288# 0.146546f
C42 plus.t10 a_n1626_n3288# 0.291362f
C43 plus.n3 a_n1626_n3288# 0.124411f
C44 plus.t8 a_n1626_n3288# 0.291362f
C45 plus.n4 a_n1626_n3288# 0.124411f
C46 plus.n5 a_n1626_n3288# 0.0243f
C47 plus.n6 a_n1626_n3288# 0.128606f
C48 plus.n7 a_n1626_n3288# 0.057282f
C49 plus.n8 a_n1626_n3288# 0.057282f
C50 plus.n9 a_n1626_n3288# 0.021651f
C51 plus.n10 a_n1626_n3288# 0.124411f
C52 plus.n11 a_n1626_n3288# 0.0243f
C53 plus.n12 a_n1626_n3288# 0.124411f
C54 plus.t9 a_n1626_n3288# 0.294494f
C55 plus.n13 a_n1626_n3288# 0.146462f
C56 plus.n14 a_n1626_n3288# 0.646664f
C57 plus.n15 a_n1626_n3288# 0.057282f
C58 plus.t0 a_n1626_n3288# 0.294494f
C59 plus.t4 a_n1626_n3288# 0.291362f
C60 plus.t2 a_n1626_n3288# 0.291362f
C61 plus.n16 a_n1626_n3288# 0.021651f
C62 plus.t3 a_n1626_n3288# 0.294494f
C63 plus.n17 a_n1626_n3288# 0.146546f
C64 plus.t1 a_n1626_n3288# 0.291362f
C65 plus.n18 a_n1626_n3288# 0.124411f
C66 plus.t5 a_n1626_n3288# 0.291362f
C67 plus.n19 a_n1626_n3288# 0.124411f
C68 plus.n20 a_n1626_n3288# 0.0243f
C69 plus.n21 a_n1626_n3288# 0.128606f
C70 plus.n22 a_n1626_n3288# 0.057282f
C71 plus.n23 a_n1626_n3288# 0.057282f
C72 plus.n24 a_n1626_n3288# 0.021651f
C73 plus.n25 a_n1626_n3288# 0.124411f
C74 plus.n26 a_n1626_n3288# 0.0243f
C75 plus.n27 a_n1626_n3288# 0.124411f
C76 plus.n28 a_n1626_n3288# 0.146462f
C77 plus.n29 a_n1626_n3288# 1.6471f
C78 source.t2 a_n1626_n3288# 2.51896f
C79 source.n0 a_n1626_n3288# 1.25619f
C80 source.t1 a_n1626_n3288# 0.325531f
C81 source.t11 a_n1626_n3288# 0.325531f
C82 source.n1 a_n1626_n3288# 2.06091f
C83 source.n2 a_n1626_n3288# 0.313455f
C84 source.t9 a_n1626_n3288# 0.325531f
C85 source.t5 a_n1626_n3288# 0.325531f
C86 source.n3 a_n1626_n3288# 2.06091f
C87 source.n4 a_n1626_n3288# 0.313455f
C88 source.t10 a_n1626_n3288# 2.51897f
C89 source.n5 a_n1626_n3288# 0.434749f
C90 source.t20 a_n1626_n3288# 2.51897f
C91 source.n6 a_n1626_n3288# 0.434749f
C92 source.t15 a_n1626_n3288# 0.325531f
C93 source.t21 a_n1626_n3288# 0.325531f
C94 source.n7 a_n1626_n3288# 2.06091f
C95 source.n8 a_n1626_n3288# 0.313455f
C96 source.t19 a_n1626_n3288# 0.325531f
C97 source.t17 a_n1626_n3288# 0.325531f
C98 source.n9 a_n1626_n3288# 2.06091f
C99 source.n10 a_n1626_n3288# 0.313455f
C100 source.t14 a_n1626_n3288# 2.51897f
C101 source.n11 a_n1626_n3288# 1.61289f
C102 source.t3 a_n1626_n3288# 2.51896f
C103 source.n12 a_n1626_n3288# 1.6129f
C104 source.t8 a_n1626_n3288# 0.325531f
C105 source.t4 a_n1626_n3288# 0.325531f
C106 source.n13 a_n1626_n3288# 2.0609f
C107 source.n14 a_n1626_n3288# 0.313466f
C108 source.t7 a_n1626_n3288# 0.325531f
C109 source.t0 a_n1626_n3288# 0.325531f
C110 source.n15 a_n1626_n3288# 2.0609f
C111 source.n16 a_n1626_n3288# 0.313466f
C112 source.t6 a_n1626_n3288# 2.51896f
C113 source.n17 a_n1626_n3288# 0.43476f
C114 source.t23 a_n1626_n3288# 2.51896f
C115 source.n18 a_n1626_n3288# 0.43476f
C116 source.t18 a_n1626_n3288# 0.325531f
C117 source.t13 a_n1626_n3288# 0.325531f
C118 source.n19 a_n1626_n3288# 2.0609f
C119 source.n20 a_n1626_n3288# 0.313466f
C120 source.t12 a_n1626_n3288# 0.325531f
C121 source.t22 a_n1626_n3288# 0.325531f
C122 source.n21 a_n1626_n3288# 2.0609f
C123 source.n22 a_n1626_n3288# 0.313466f
C124 source.t16 a_n1626_n3288# 2.51896f
C125 source.n23 a_n1626_n3288# 0.563664f
C126 source.n24 a_n1626_n3288# 1.42207f
C127 drain_right.t5 a_n1626_n3288# 0.40425f
C128 drain_right.t7 a_n1626_n3288# 0.40425f
C129 drain_right.n0 a_n1626_n3288# 2.65195f
C130 drain_right.t2 a_n1626_n3288# 0.40425f
C131 drain_right.t0 a_n1626_n3288# 0.40425f
C132 drain_right.n1 a_n1626_n3288# 2.64904f
C133 drain_right.t11 a_n1626_n3288# 0.40425f
C134 drain_right.t8 a_n1626_n3288# 0.40425f
C135 drain_right.n2 a_n1626_n3288# 2.65195f
C136 drain_right.n3 a_n1626_n3288# 2.23147f
C137 drain_right.t4 a_n1626_n3288# 0.40425f
C138 drain_right.t9 a_n1626_n3288# 0.40425f
C139 drain_right.n4 a_n1626_n3288# 2.6523f
C140 drain_right.t10 a_n1626_n3288# 0.40425f
C141 drain_right.t6 a_n1626_n3288# 0.40425f
C142 drain_right.n5 a_n1626_n3288# 2.64905f
C143 drain_right.n6 a_n1626_n3288# 0.683535f
C144 drain_right.t3 a_n1626_n3288# 0.40425f
C145 drain_right.t1 a_n1626_n3288# 0.40425f
C146 drain_right.n7 a_n1626_n3288# 2.64905f
C147 drain_right.n8 a_n1626_n3288# 0.572687f
C148 minus.n0 a_n1626_n3288# 0.056117f
C149 minus.t9 a_n1626_n3288# 0.288506f
C150 minus.t4 a_n1626_n3288# 0.285438f
C151 minus.t6 a_n1626_n3288# 0.285438f
C152 minus.n1 a_n1626_n3288# 0.021211f
C153 minus.t3 a_n1626_n3288# 0.288506f
C154 minus.n2 a_n1626_n3288# 0.143566f
C155 minus.t8 a_n1626_n3288# 0.285438f
C156 minus.n3 a_n1626_n3288# 0.121881f
C157 minus.t2 a_n1626_n3288# 0.285438f
C158 minus.n4 a_n1626_n3288# 0.121881f
C159 minus.n5 a_n1626_n3288# 0.023806f
C160 minus.n6 a_n1626_n3288# 0.125992f
C161 minus.n7 a_n1626_n3288# 0.056117f
C162 minus.n8 a_n1626_n3288# 0.056117f
C163 minus.n9 a_n1626_n3288# 0.021211f
C164 minus.n10 a_n1626_n3288# 0.121881f
C165 minus.n11 a_n1626_n3288# 0.023806f
C166 minus.n12 a_n1626_n3288# 0.121881f
C167 minus.n13 a_n1626_n3288# 0.143484f
C168 minus.n14 a_n1626_n3288# 1.91058f
C169 minus.n15 a_n1626_n3288# 0.056117f
C170 minus.t1 a_n1626_n3288# 0.285438f
C171 minus.t11 a_n1626_n3288# 0.285438f
C172 minus.n16 a_n1626_n3288# 0.021211f
C173 minus.t0 a_n1626_n3288# 0.288506f
C174 minus.n17 a_n1626_n3288# 0.143566f
C175 minus.t5 a_n1626_n3288# 0.285438f
C176 minus.n18 a_n1626_n3288# 0.121881f
C177 minus.t10 a_n1626_n3288# 0.285438f
C178 minus.n19 a_n1626_n3288# 0.121881f
C179 minus.n20 a_n1626_n3288# 0.023806f
C180 minus.n21 a_n1626_n3288# 0.125992f
C181 minus.n22 a_n1626_n3288# 0.056117f
C182 minus.n23 a_n1626_n3288# 0.056117f
C183 minus.n24 a_n1626_n3288# 0.021211f
C184 minus.n25 a_n1626_n3288# 0.121881f
C185 minus.n26 a_n1626_n3288# 0.023806f
C186 minus.n27 a_n1626_n3288# 0.121881f
C187 minus.t7 a_n1626_n3288# 0.288506f
C188 minus.n28 a_n1626_n3288# 0.143484f
C189 minus.n29 a_n1626_n3288# 0.372443f
C190 minus.n30 a_n1626_n3288# 2.32469f
.ends

