* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t24 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X1 drain_left.t18 plus.t1 source.t25 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X2 drain_left.t17 plus.t2 source.t32 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X3 source.t36 plus.t3 drain_left.t16 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X4 a_n1992_n1288# a_n1992_n1288# a_n1992_n1288# a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.25
X5 drain_left.t15 plus.t4 source.t27 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X6 source.t15 minus.t0 drain_right.t19 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X7 drain_left.t14 plus.t5 source.t37 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X8 source.t9 minus.t1 drain_right.t18 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X9 a_n1992_n1288# a_n1992_n1288# a_n1992_n1288# a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X10 source.t20 plus.t6 drain_left.t13 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X11 source.t30 plus.t7 drain_left.t12 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X12 source.t22 plus.t8 drain_left.t11 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X13 source.t34 plus.t9 drain_left.t10 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X14 drain_right.t17 minus.t2 source.t8 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X15 source.t2 minus.t3 drain_right.t16 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X16 drain_left.t9 plus.t10 source.t29 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X17 source.t6 minus.t4 drain_right.t15 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X18 drain_right.t14 minus.t5 source.t10 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X19 source.t11 minus.t6 drain_right.t13 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X20 source.t16 minus.t7 drain_right.t12 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X21 source.t31 plus.t11 drain_left.t8 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X22 source.t33 plus.t12 drain_left.t7 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X23 source.t23 plus.t13 drain_left.t6 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X24 source.t1 minus.t8 drain_right.t11 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X25 source.t3 minus.t9 drain_right.t10 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X26 source.t39 minus.t10 drain_right.t9 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.25
X27 drain_right.t8 minus.t11 source.t5 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X28 a_n1992_n1288# a_n1992_n1288# a_n1992_n1288# a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X29 source.t26 plus.t14 drain_left.t5 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X30 drain_right.t7 minus.t12 source.t0 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X31 drain_right.t6 minus.t13 source.t4 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X32 source.t14 minus.t14 drain_right.t5 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X33 a_n1992_n1288# a_n1992_n1288# a_n1992_n1288# a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.25
X34 drain_right.t4 minus.t15 source.t12 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X35 drain_right.t3 minus.t16 source.t17 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X36 source.t18 plus.t15 drain_left.t4 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X37 drain_right.t2 minus.t17 source.t38 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X38 drain_right.t1 minus.t18 source.t13 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X39 drain_right.t0 minus.t19 source.t7 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X40 drain_left.t3 plus.t16 source.t35 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X41 drain_left.t2 plus.t17 source.t28 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.25
X42 drain_left.t1 plus.t18 source.t21 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
X43 drain_left.t0 plus.t19 source.t19 a_n1992_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.25
R0 plus.n6 plus.t8 370.702
R1 plus.n25 plus.t4 370.702
R2 plus.n33 plus.t17 370.702
R3 plus.n52 plus.t9 370.702
R4 plus.n5 plus.t1 318.12
R5 plus.n9 plus.t13 318.12
R6 plus.n11 plus.t0 318.12
R7 plus.n3 plus.t12 318.12
R8 plus.n17 plus.t18 318.12
R9 plus.n1 plus.t11 318.12
R10 plus.n22 plus.t5 318.12
R11 plus.n24 plus.t14 318.12
R12 plus.n32 plus.t15 318.12
R13 plus.n36 plus.t2 318.12
R14 plus.n38 plus.t7 318.12
R15 plus.n30 plus.t16 318.12
R16 plus.n44 plus.t3 318.12
R17 plus.n28 plus.t19 318.12
R18 plus.n49 plus.t6 318.12
R19 plus.n51 plus.t10 318.12
R20 plus.n7 plus.n6 161.489
R21 plus.n34 plus.n33 161.489
R22 plus.n8 plus.n7 161.3
R23 plus.n10 plus.n4 161.3
R24 plus.n13 plus.n12 161.3
R25 plus.n15 plus.n14 161.3
R26 plus.n16 plus.n2 161.3
R27 plus.n19 plus.n18 161.3
R28 plus.n21 plus.n20 161.3
R29 plus.n23 plus.n0 161.3
R30 plus.n26 plus.n25 161.3
R31 plus.n35 plus.n34 161.3
R32 plus.n37 plus.n31 161.3
R33 plus.n40 plus.n39 161.3
R34 plus.n42 plus.n41 161.3
R35 plus.n43 plus.n29 161.3
R36 plus.n46 plus.n45 161.3
R37 plus.n48 plus.n47 161.3
R38 plus.n50 plus.n27 161.3
R39 plus.n53 plus.n52 161.3
R40 plus.n16 plus.n15 73.0308
R41 plus.n43 plus.n42 73.0308
R42 plus.n12 plus.n3 67.1884
R43 plus.n18 plus.n17 67.1884
R44 plus.n45 plus.n44 67.1884
R45 plus.n39 plus.n30 67.1884
R46 plus.n11 plus.n10 55.5035
R47 plus.n21 plus.n1 55.5035
R48 plus.n48 plus.n28 55.5035
R49 plus.n38 plus.n37 55.5035
R50 plus.n9 plus.n8 43.8187
R51 plus.n23 plus.n22 43.8187
R52 plus.n50 plus.n49 43.8187
R53 plus.n36 plus.n35 43.8187
R54 plus.n8 plus.n5 40.8975
R55 plus.n24 plus.n23 40.8975
R56 plus.n51 plus.n50 40.8975
R57 plus.n35 plus.n32 40.8975
R58 plus.n6 plus.n5 32.1338
R59 plus.n25 plus.n24 32.1338
R60 plus.n52 plus.n51 32.1338
R61 plus.n33 plus.n32 32.1338
R62 plus.n10 plus.n9 29.2126
R63 plus.n22 plus.n21 29.2126
R64 plus.n49 plus.n48 29.2126
R65 plus.n37 plus.n36 29.2126
R66 plus plus.n53 26.7566
R67 plus.n12 plus.n11 17.5278
R68 plus.n18 plus.n1 17.5278
R69 plus.n45 plus.n28 17.5278
R70 plus.n39 plus.n38 17.5278
R71 plus plus.n26 8.35277
R72 plus.n15 plus.n3 5.84292
R73 plus.n17 plus.n16 5.84292
R74 plus.n44 plus.n43 5.84292
R75 plus.n42 plus.n30 5.84292
R76 plus.n7 plus.n4 0.189894
R77 plus.n13 plus.n4 0.189894
R78 plus.n14 plus.n13 0.189894
R79 plus.n14 plus.n2 0.189894
R80 plus.n19 plus.n2 0.189894
R81 plus.n20 plus.n19 0.189894
R82 plus.n20 plus.n0 0.189894
R83 plus.n26 plus.n0 0.189894
R84 plus.n53 plus.n27 0.189894
R85 plus.n47 plus.n27 0.189894
R86 plus.n47 plus.n46 0.189894
R87 plus.n46 plus.n29 0.189894
R88 plus.n41 plus.n29 0.189894
R89 plus.n41 plus.n40 0.189894
R90 plus.n40 plus.n31 0.189894
R91 plus.n34 plus.n31 0.189894
R92 source.n90 source.n88 289.615
R93 source.n74 source.n72 289.615
R94 source.n66 source.n64 289.615
R95 source.n50 source.n48 289.615
R96 source.n2 source.n0 289.615
R97 source.n18 source.n16 289.615
R98 source.n26 source.n24 289.615
R99 source.n42 source.n40 289.615
R100 source.n91 source.n90 185
R101 source.n75 source.n74 185
R102 source.n67 source.n66 185
R103 source.n51 source.n50 185
R104 source.n3 source.n2 185
R105 source.n19 source.n18 185
R106 source.n27 source.n26 185
R107 source.n43 source.n42 185
R108 source.t12 source.n89 167.117
R109 source.t39 source.n73 167.117
R110 source.t28 source.n65 167.117
R111 source.t34 source.n49 167.117
R112 source.t27 source.n1 167.117
R113 source.t22 source.n17 167.117
R114 source.t0 source.n25 167.117
R115 source.t11 source.n41 167.117
R116 source.n9 source.n8 84.1169
R117 source.n11 source.n10 84.1169
R118 source.n13 source.n12 84.1169
R119 source.n15 source.n14 84.1169
R120 source.n33 source.n32 84.1169
R121 source.n35 source.n34 84.1169
R122 source.n37 source.n36 84.1169
R123 source.n39 source.n38 84.1169
R124 source.n87 source.n86 84.1168
R125 source.n85 source.n84 84.1168
R126 source.n83 source.n82 84.1168
R127 source.n81 source.n80 84.1168
R128 source.n63 source.n62 84.1168
R129 source.n61 source.n60 84.1168
R130 source.n59 source.n58 84.1168
R131 source.n57 source.n56 84.1168
R132 source.n90 source.t12 52.3082
R133 source.n74 source.t39 52.3082
R134 source.n66 source.t28 52.3082
R135 source.n50 source.t34 52.3082
R136 source.n2 source.t27 52.3082
R137 source.n18 source.t22 52.3082
R138 source.n26 source.t0 52.3082
R139 source.n42 source.t11 52.3082
R140 source.n95 source.n94 31.4096
R141 source.n79 source.n78 31.4096
R142 source.n71 source.n70 31.4096
R143 source.n55 source.n54 31.4096
R144 source.n7 source.n6 31.4096
R145 source.n23 source.n22 31.4096
R146 source.n31 source.n30 31.4096
R147 source.n47 source.n46 31.4096
R148 source.n55 source.n47 14.212
R149 source.n86 source.t4 9.9005
R150 source.n86 source.t1 9.9005
R151 source.n84 source.t17 9.9005
R152 source.n84 source.t14 9.9005
R153 source.n82 source.t10 9.9005
R154 source.n82 source.t3 9.9005
R155 source.n80 source.t8 9.9005
R156 source.n80 source.t16 9.9005
R157 source.n62 source.t32 9.9005
R158 source.n62 source.t18 9.9005
R159 source.n60 source.t35 9.9005
R160 source.n60 source.t30 9.9005
R161 source.n58 source.t19 9.9005
R162 source.n58 source.t36 9.9005
R163 source.n56 source.t29 9.9005
R164 source.n56 source.t20 9.9005
R165 source.n8 source.t37 9.9005
R166 source.n8 source.t26 9.9005
R167 source.n10 source.t21 9.9005
R168 source.n10 source.t31 9.9005
R169 source.n12 source.t24 9.9005
R170 source.n12 source.t33 9.9005
R171 source.n14 source.t25 9.9005
R172 source.n14 source.t23 9.9005
R173 source.n32 source.t5 9.9005
R174 source.n32 source.t9 9.9005
R175 source.n34 source.t38 9.9005
R176 source.n34 source.t15 9.9005
R177 source.n36 source.t13 9.9005
R178 source.n36 source.t6 9.9005
R179 source.n38 source.t7 9.9005
R180 source.n38 source.t2 9.9005
R181 source.n91 source.n89 9.71174
R182 source.n75 source.n73 9.71174
R183 source.n67 source.n65 9.71174
R184 source.n51 source.n49 9.71174
R185 source.n3 source.n1 9.71174
R186 source.n19 source.n17 9.71174
R187 source.n27 source.n25 9.71174
R188 source.n43 source.n41 9.71174
R189 source.n94 source.n93 9.45567
R190 source.n78 source.n77 9.45567
R191 source.n70 source.n69 9.45567
R192 source.n54 source.n53 9.45567
R193 source.n6 source.n5 9.45567
R194 source.n22 source.n21 9.45567
R195 source.n30 source.n29 9.45567
R196 source.n46 source.n45 9.45567
R197 source.n93 source.n92 9.3005
R198 source.n77 source.n76 9.3005
R199 source.n69 source.n68 9.3005
R200 source.n53 source.n52 9.3005
R201 source.n5 source.n4 9.3005
R202 source.n21 source.n20 9.3005
R203 source.n29 source.n28 9.3005
R204 source.n45 source.n44 9.3005
R205 source.n96 source.n7 8.69904
R206 source.n94 source.n88 8.14595
R207 source.n78 source.n72 8.14595
R208 source.n70 source.n64 8.14595
R209 source.n54 source.n48 8.14595
R210 source.n6 source.n0 8.14595
R211 source.n22 source.n16 8.14595
R212 source.n30 source.n24 8.14595
R213 source.n46 source.n40 8.14595
R214 source.n92 source.n91 7.3702
R215 source.n76 source.n75 7.3702
R216 source.n68 source.n67 7.3702
R217 source.n52 source.n51 7.3702
R218 source.n4 source.n3 7.3702
R219 source.n20 source.n19 7.3702
R220 source.n28 source.n27 7.3702
R221 source.n44 source.n43 7.3702
R222 source.n92 source.n88 5.81868
R223 source.n76 source.n72 5.81868
R224 source.n68 source.n64 5.81868
R225 source.n52 source.n48 5.81868
R226 source.n4 source.n0 5.81868
R227 source.n20 source.n16 5.81868
R228 source.n28 source.n24 5.81868
R229 source.n44 source.n40 5.81868
R230 source.n96 source.n95 5.51343
R231 source.n93 source.n89 3.44771
R232 source.n77 source.n73 3.44771
R233 source.n69 source.n65 3.44771
R234 source.n53 source.n49 3.44771
R235 source.n5 source.n1 3.44771
R236 source.n21 source.n17 3.44771
R237 source.n29 source.n25 3.44771
R238 source.n45 source.n41 3.44771
R239 source.n47 source.n39 0.5005
R240 source.n39 source.n37 0.5005
R241 source.n37 source.n35 0.5005
R242 source.n35 source.n33 0.5005
R243 source.n33 source.n31 0.5005
R244 source.n23 source.n15 0.5005
R245 source.n15 source.n13 0.5005
R246 source.n13 source.n11 0.5005
R247 source.n11 source.n9 0.5005
R248 source.n9 source.n7 0.5005
R249 source.n57 source.n55 0.5005
R250 source.n59 source.n57 0.5005
R251 source.n61 source.n59 0.5005
R252 source.n63 source.n61 0.5005
R253 source.n71 source.n63 0.5005
R254 source.n81 source.n79 0.5005
R255 source.n83 source.n81 0.5005
R256 source.n85 source.n83 0.5005
R257 source.n87 source.n85 0.5005
R258 source.n95 source.n87 0.5005
R259 source.n31 source.n23 0.470328
R260 source.n79 source.n71 0.470328
R261 source source.n96 0.188
R262 drain_left.n10 drain_left.n8 101.296
R263 drain_left.n6 drain_left.n4 101.296
R264 drain_left.n2 drain_left.n0 101.296
R265 drain_left.n16 drain_left.n15 100.796
R266 drain_left.n14 drain_left.n13 100.796
R267 drain_left.n12 drain_left.n11 100.796
R268 drain_left.n10 drain_left.n9 100.796
R269 drain_left.n7 drain_left.n3 100.796
R270 drain_left.n6 drain_left.n5 100.796
R271 drain_left.n2 drain_left.n1 100.796
R272 drain_left drain_left.n7 23.7913
R273 drain_left.n3 drain_left.t16 9.9005
R274 drain_left.n3 drain_left.t3 9.9005
R275 drain_left.n4 drain_left.t4 9.9005
R276 drain_left.n4 drain_left.t2 9.9005
R277 drain_left.n5 drain_left.t12 9.9005
R278 drain_left.n5 drain_left.t17 9.9005
R279 drain_left.n1 drain_left.t13 9.9005
R280 drain_left.n1 drain_left.t0 9.9005
R281 drain_left.n0 drain_left.t10 9.9005
R282 drain_left.n0 drain_left.t9 9.9005
R283 drain_left.n15 drain_left.t5 9.9005
R284 drain_left.n15 drain_left.t15 9.9005
R285 drain_left.n13 drain_left.t8 9.9005
R286 drain_left.n13 drain_left.t14 9.9005
R287 drain_left.n11 drain_left.t7 9.9005
R288 drain_left.n11 drain_left.t1 9.9005
R289 drain_left.n9 drain_left.t6 9.9005
R290 drain_left.n9 drain_left.t19 9.9005
R291 drain_left.n8 drain_left.t11 9.9005
R292 drain_left.n8 drain_left.t18 9.9005
R293 drain_left drain_left.n16 6.15322
R294 drain_left.n12 drain_left.n10 0.5005
R295 drain_left.n14 drain_left.n12 0.5005
R296 drain_left.n16 drain_left.n14 0.5005
R297 drain_left.n7 drain_left.n6 0.445154
R298 drain_left.n7 drain_left.n2 0.445154
R299 minus.n25 minus.t6 370.702
R300 minus.n6 minus.t12 370.702
R301 minus.n52 minus.t15 370.702
R302 minus.n33 minus.t10 370.702
R303 minus.n24 minus.t19 318.12
R304 minus.n22 minus.t3 318.12
R305 minus.n1 minus.t18 318.12
R306 minus.n17 minus.t4 318.12
R307 minus.n3 minus.t17 318.12
R308 minus.n11 minus.t0 318.12
R309 minus.n9 minus.t11 318.12
R310 minus.n5 minus.t1 318.12
R311 minus.n51 minus.t8 318.12
R312 minus.n49 minus.t13 318.12
R313 minus.n28 minus.t14 318.12
R314 minus.n44 minus.t16 318.12
R315 minus.n30 minus.t9 318.12
R316 minus.n38 minus.t5 318.12
R317 minus.n36 minus.t7 318.12
R318 minus.n32 minus.t2 318.12
R319 minus.n7 minus.n6 161.489
R320 minus.n34 minus.n33 161.489
R321 minus.n26 minus.n25 161.3
R322 minus.n23 minus.n0 161.3
R323 minus.n21 minus.n20 161.3
R324 minus.n19 minus.n18 161.3
R325 minus.n16 minus.n2 161.3
R326 minus.n15 minus.n14 161.3
R327 minus.n13 minus.n12 161.3
R328 minus.n10 minus.n4 161.3
R329 minus.n8 minus.n7 161.3
R330 minus.n53 minus.n52 161.3
R331 minus.n50 minus.n27 161.3
R332 minus.n48 minus.n47 161.3
R333 minus.n46 minus.n45 161.3
R334 minus.n43 minus.n29 161.3
R335 minus.n42 minus.n41 161.3
R336 minus.n40 minus.n39 161.3
R337 minus.n37 minus.n31 161.3
R338 minus.n35 minus.n34 161.3
R339 minus.n16 minus.n15 73.0308
R340 minus.n43 minus.n42 73.0308
R341 minus.n18 minus.n17 67.1884
R342 minus.n12 minus.n3 67.1884
R343 minus.n39 minus.n30 67.1884
R344 minus.n45 minus.n44 67.1884
R345 minus.n21 minus.n1 55.5035
R346 minus.n11 minus.n10 55.5035
R347 minus.n38 minus.n37 55.5035
R348 minus.n48 minus.n28 55.5035
R349 minus.n23 minus.n22 43.8187
R350 minus.n9 minus.n8 43.8187
R351 minus.n36 minus.n35 43.8187
R352 minus.n50 minus.n49 43.8187
R353 minus.n24 minus.n23 40.8975
R354 minus.n8 minus.n5 40.8975
R355 minus.n35 minus.n32 40.8975
R356 minus.n51 minus.n50 40.8975
R357 minus.n25 minus.n24 32.1338
R358 minus.n6 minus.n5 32.1338
R359 minus.n33 minus.n32 32.1338
R360 minus.n52 minus.n51 32.1338
R361 minus.n22 minus.n21 29.2126
R362 minus.n10 minus.n9 29.2126
R363 minus.n37 minus.n36 29.2126
R364 minus.n49 minus.n48 29.2126
R365 minus.n54 minus.n26 29.0876
R366 minus.n18 minus.n1 17.5278
R367 minus.n12 minus.n11 17.5278
R368 minus.n39 minus.n38 17.5278
R369 minus.n45 minus.n28 17.5278
R370 minus.n54 minus.n53 6.49671
R371 minus.n17 minus.n16 5.84292
R372 minus.n15 minus.n3 5.84292
R373 minus.n42 minus.n30 5.84292
R374 minus.n44 minus.n43 5.84292
R375 minus.n26 minus.n0 0.189894
R376 minus.n20 minus.n0 0.189894
R377 minus.n20 minus.n19 0.189894
R378 minus.n19 minus.n2 0.189894
R379 minus.n14 minus.n2 0.189894
R380 minus.n14 minus.n13 0.189894
R381 minus.n13 minus.n4 0.189894
R382 minus.n7 minus.n4 0.189894
R383 minus.n34 minus.n31 0.189894
R384 minus.n40 minus.n31 0.189894
R385 minus.n41 minus.n40 0.189894
R386 minus.n41 minus.n29 0.189894
R387 minus.n46 minus.n29 0.189894
R388 minus.n47 minus.n46 0.189894
R389 minus.n47 minus.n27 0.189894
R390 minus.n53 minus.n27 0.189894
R391 minus minus.n54 0.188
R392 drain_right.n10 drain_right.n8 101.296
R393 drain_right.n6 drain_right.n4 101.296
R394 drain_right.n2 drain_right.n0 101.296
R395 drain_right.n10 drain_right.n9 100.796
R396 drain_right.n12 drain_right.n11 100.796
R397 drain_right.n14 drain_right.n13 100.796
R398 drain_right.n16 drain_right.n15 100.796
R399 drain_right.n7 drain_right.n3 100.796
R400 drain_right.n6 drain_right.n5 100.796
R401 drain_right.n2 drain_right.n1 100.796
R402 drain_right drain_right.n7 23.2381
R403 drain_right.n3 drain_right.t10 9.9005
R404 drain_right.n3 drain_right.t3 9.9005
R405 drain_right.n4 drain_right.t11 9.9005
R406 drain_right.n4 drain_right.t4 9.9005
R407 drain_right.n5 drain_right.t5 9.9005
R408 drain_right.n5 drain_right.t6 9.9005
R409 drain_right.n1 drain_right.t12 9.9005
R410 drain_right.n1 drain_right.t14 9.9005
R411 drain_right.n0 drain_right.t9 9.9005
R412 drain_right.n0 drain_right.t17 9.9005
R413 drain_right.n8 drain_right.t18 9.9005
R414 drain_right.n8 drain_right.t7 9.9005
R415 drain_right.n9 drain_right.t19 9.9005
R416 drain_right.n9 drain_right.t8 9.9005
R417 drain_right.n11 drain_right.t15 9.9005
R418 drain_right.n11 drain_right.t2 9.9005
R419 drain_right.n13 drain_right.t16 9.9005
R420 drain_right.n13 drain_right.t1 9.9005
R421 drain_right.n15 drain_right.t13 9.9005
R422 drain_right.n15 drain_right.t0 9.9005
R423 drain_right drain_right.n16 6.15322
R424 drain_right.n16 drain_right.n14 0.5005
R425 drain_right.n14 drain_right.n12 0.5005
R426 drain_right.n12 drain_right.n10 0.5005
R427 drain_right.n7 drain_right.n6 0.445154
R428 drain_right.n7 drain_right.n2 0.445154
C0 plus drain_left 1.72704f
C1 source drain_left 9.51204f
C2 plus minus 3.79425f
C3 minus source 1.75935f
C4 plus drain_right 0.355923f
C5 source drain_right 9.51227f
C6 minus drain_left 0.177702f
C7 drain_right drain_left 1.04677f
C8 minus drain_right 1.53257f
C9 plus source 1.77332f
C10 drain_right a_n1992_n1288# 4.28383f
C11 drain_left a_n1992_n1288# 4.56005f
C12 source a_n1992_n1288# 3.185815f
C13 minus a_n1992_n1288# 6.967883f
C14 plus a_n1992_n1288# 7.588521f
C15 drain_right.t9 a_n1992_n1288# 0.045402f
C16 drain_right.t17 a_n1992_n1288# 0.045402f
C17 drain_right.n0 a_n1992_n1288# 0.286829f
C18 drain_right.t12 a_n1992_n1288# 0.045402f
C19 drain_right.t14 a_n1992_n1288# 0.045402f
C20 drain_right.n1 a_n1992_n1288# 0.28523f
C21 drain_right.n2 a_n1992_n1288# 0.631226f
C22 drain_right.t10 a_n1992_n1288# 0.045402f
C23 drain_right.t3 a_n1992_n1288# 0.045402f
C24 drain_right.n3 a_n1992_n1288# 0.28523f
C25 drain_right.t11 a_n1992_n1288# 0.045402f
C26 drain_right.t4 a_n1992_n1288# 0.045402f
C27 drain_right.n4 a_n1992_n1288# 0.286829f
C28 drain_right.t5 a_n1992_n1288# 0.045402f
C29 drain_right.t6 a_n1992_n1288# 0.045402f
C30 drain_right.n5 a_n1992_n1288# 0.28523f
C31 drain_right.n6 a_n1992_n1288# 0.631226f
C32 drain_right.n7 a_n1992_n1288# 1.07099f
C33 drain_right.t18 a_n1992_n1288# 0.045402f
C34 drain_right.t7 a_n1992_n1288# 0.045402f
C35 drain_right.n8 a_n1992_n1288# 0.28683f
C36 drain_right.t19 a_n1992_n1288# 0.045402f
C37 drain_right.t8 a_n1992_n1288# 0.045402f
C38 drain_right.n9 a_n1992_n1288# 0.285231f
C39 drain_right.n10 a_n1992_n1288# 0.634849f
C40 drain_right.t15 a_n1992_n1288# 0.045402f
C41 drain_right.t2 a_n1992_n1288# 0.045402f
C42 drain_right.n11 a_n1992_n1288# 0.285231f
C43 drain_right.n12 a_n1992_n1288# 0.312439f
C44 drain_right.t16 a_n1992_n1288# 0.045402f
C45 drain_right.t1 a_n1992_n1288# 0.045402f
C46 drain_right.n13 a_n1992_n1288# 0.285231f
C47 drain_right.n14 a_n1992_n1288# 0.312439f
C48 drain_right.t13 a_n1992_n1288# 0.045402f
C49 drain_right.t0 a_n1992_n1288# 0.045402f
C50 drain_right.n15 a_n1992_n1288# 0.285231f
C51 drain_right.n16 a_n1992_n1288# 0.549561f
C52 minus.n0 a_n1992_n1288# 0.027201f
C53 minus.t6 a_n1992_n1288# 0.044446f
C54 minus.t19 a_n1992_n1288# 0.040021f
C55 minus.t3 a_n1992_n1288# 0.040021f
C56 minus.t18 a_n1992_n1288# 0.040021f
C57 minus.n1 a_n1992_n1288# 0.029349f
C58 minus.n2 a_n1992_n1288# 0.027201f
C59 minus.t4 a_n1992_n1288# 0.040021f
C60 minus.t17 a_n1992_n1288# 0.040021f
C61 minus.n3 a_n1992_n1288# 0.029349f
C62 minus.n4 a_n1992_n1288# 0.027201f
C63 minus.t0 a_n1992_n1288# 0.040021f
C64 minus.t11 a_n1992_n1288# 0.040021f
C65 minus.t1 a_n1992_n1288# 0.040021f
C66 minus.n5 a_n1992_n1288# 0.029349f
C67 minus.t12 a_n1992_n1288# 0.044446f
C68 minus.n6 a_n1992_n1288# 0.037175f
C69 minus.n7 a_n1992_n1288# 0.062244f
C70 minus.n8 a_n1992_n1288# 0.010365f
C71 minus.n9 a_n1992_n1288# 0.029349f
C72 minus.n10 a_n1992_n1288# 0.010365f
C73 minus.n11 a_n1992_n1288# 0.029349f
C74 minus.n12 a_n1992_n1288# 0.010365f
C75 minus.n13 a_n1992_n1288# 0.027201f
C76 minus.n14 a_n1992_n1288# 0.027201f
C77 minus.n15 a_n1992_n1288# 0.009694f
C78 minus.n16 a_n1992_n1288# 0.009694f
C79 minus.n17 a_n1992_n1288# 0.029349f
C80 minus.n18 a_n1992_n1288# 0.010365f
C81 minus.n19 a_n1992_n1288# 0.027201f
C82 minus.n20 a_n1992_n1288# 0.027201f
C83 minus.n21 a_n1992_n1288# 0.010365f
C84 minus.n22 a_n1992_n1288# 0.029349f
C85 minus.n23 a_n1992_n1288# 0.010365f
C86 minus.n24 a_n1992_n1288# 0.029349f
C87 minus.n25 a_n1992_n1288# 0.037134f
C88 minus.n26 a_n1992_n1288# 0.670901f
C89 minus.n27 a_n1992_n1288# 0.027201f
C90 minus.t8 a_n1992_n1288# 0.040021f
C91 minus.t13 a_n1992_n1288# 0.040021f
C92 minus.t14 a_n1992_n1288# 0.040021f
C93 minus.n28 a_n1992_n1288# 0.029349f
C94 minus.n29 a_n1992_n1288# 0.027201f
C95 minus.t16 a_n1992_n1288# 0.040021f
C96 minus.t9 a_n1992_n1288# 0.040021f
C97 minus.n30 a_n1992_n1288# 0.029349f
C98 minus.n31 a_n1992_n1288# 0.027201f
C99 minus.t5 a_n1992_n1288# 0.040021f
C100 minus.t7 a_n1992_n1288# 0.040021f
C101 minus.t2 a_n1992_n1288# 0.040021f
C102 minus.n32 a_n1992_n1288# 0.029349f
C103 minus.t10 a_n1992_n1288# 0.044446f
C104 minus.n33 a_n1992_n1288# 0.037175f
C105 minus.n34 a_n1992_n1288# 0.062244f
C106 minus.n35 a_n1992_n1288# 0.010365f
C107 minus.n36 a_n1992_n1288# 0.029349f
C108 minus.n37 a_n1992_n1288# 0.010365f
C109 minus.n38 a_n1992_n1288# 0.029349f
C110 minus.n39 a_n1992_n1288# 0.010365f
C111 minus.n40 a_n1992_n1288# 0.027201f
C112 minus.n41 a_n1992_n1288# 0.027201f
C113 minus.n42 a_n1992_n1288# 0.009694f
C114 minus.n43 a_n1992_n1288# 0.009694f
C115 minus.n44 a_n1992_n1288# 0.029349f
C116 minus.n45 a_n1992_n1288# 0.010365f
C117 minus.n46 a_n1992_n1288# 0.027201f
C118 minus.n47 a_n1992_n1288# 0.027201f
C119 minus.n48 a_n1992_n1288# 0.010365f
C120 minus.n49 a_n1992_n1288# 0.029349f
C121 minus.n50 a_n1992_n1288# 0.010365f
C122 minus.n51 a_n1992_n1288# 0.029349f
C123 minus.t15 a_n1992_n1288# 0.044446f
C124 minus.n52 a_n1992_n1288# 0.037134f
C125 minus.n53 a_n1992_n1288# 0.177624f
C126 minus.n54 a_n1992_n1288# 0.828825f
C127 drain_left.t10 a_n1992_n1288# 0.044871f
C128 drain_left.t9 a_n1992_n1288# 0.044871f
C129 drain_left.n0 a_n1992_n1288# 0.283476f
C130 drain_left.t13 a_n1992_n1288# 0.044871f
C131 drain_left.t0 a_n1992_n1288# 0.044871f
C132 drain_left.n1 a_n1992_n1288# 0.281895f
C133 drain_left.n2 a_n1992_n1288# 0.623846f
C134 drain_left.t16 a_n1992_n1288# 0.044871f
C135 drain_left.t3 a_n1992_n1288# 0.044871f
C136 drain_left.n3 a_n1992_n1288# 0.281895f
C137 drain_left.t4 a_n1992_n1288# 0.044871f
C138 drain_left.t2 a_n1992_n1288# 0.044871f
C139 drain_left.n4 a_n1992_n1288# 0.283476f
C140 drain_left.t12 a_n1992_n1288# 0.044871f
C141 drain_left.t17 a_n1992_n1288# 0.044871f
C142 drain_left.n5 a_n1992_n1288# 0.281895f
C143 drain_left.n6 a_n1992_n1288# 0.623846f
C144 drain_left.n7 a_n1992_n1288# 1.11401f
C145 drain_left.t11 a_n1992_n1288# 0.044871f
C146 drain_left.t18 a_n1992_n1288# 0.044871f
C147 drain_left.n8 a_n1992_n1288# 0.283477f
C148 drain_left.t6 a_n1992_n1288# 0.044871f
C149 drain_left.t19 a_n1992_n1288# 0.044871f
C150 drain_left.n9 a_n1992_n1288# 0.281896f
C151 drain_left.n10 a_n1992_n1288# 0.627426f
C152 drain_left.t7 a_n1992_n1288# 0.044871f
C153 drain_left.t1 a_n1992_n1288# 0.044871f
C154 drain_left.n11 a_n1992_n1288# 0.281896f
C155 drain_left.n12 a_n1992_n1288# 0.308786f
C156 drain_left.t8 a_n1992_n1288# 0.044871f
C157 drain_left.t14 a_n1992_n1288# 0.044871f
C158 drain_left.n13 a_n1992_n1288# 0.281896f
C159 drain_left.n14 a_n1992_n1288# 0.308786f
C160 drain_left.t5 a_n1992_n1288# 0.044871f
C161 drain_left.t15 a_n1992_n1288# 0.044871f
C162 drain_left.n15 a_n1992_n1288# 0.281896f
C163 drain_left.n16 a_n1992_n1288# 0.543136f
C164 source.n0 a_n1992_n1288# 0.04373f
C165 source.n1 a_n1992_n1288# 0.096758f
C166 source.t27 a_n1992_n1288# 0.072612f
C167 source.n2 a_n1992_n1288# 0.075727f
C168 source.n3 a_n1992_n1288# 0.024411f
C169 source.n4 a_n1992_n1288# 0.0161f
C170 source.n5 a_n1992_n1288# 0.213278f
C171 source.n6 a_n1992_n1288# 0.047938f
C172 source.n7 a_n1992_n1288# 0.444966f
C173 source.t37 a_n1992_n1288# 0.047352f
C174 source.t26 a_n1992_n1288# 0.047352f
C175 source.n8 a_n1992_n1288# 0.253144f
C176 source.n9 a_n1992_n1288# 0.329475f
C177 source.t21 a_n1992_n1288# 0.047352f
C178 source.t31 a_n1992_n1288# 0.047352f
C179 source.n10 a_n1992_n1288# 0.253144f
C180 source.n11 a_n1992_n1288# 0.329475f
C181 source.t24 a_n1992_n1288# 0.047352f
C182 source.t33 a_n1992_n1288# 0.047352f
C183 source.n12 a_n1992_n1288# 0.253144f
C184 source.n13 a_n1992_n1288# 0.329475f
C185 source.t25 a_n1992_n1288# 0.047352f
C186 source.t23 a_n1992_n1288# 0.047352f
C187 source.n14 a_n1992_n1288# 0.253144f
C188 source.n15 a_n1992_n1288# 0.329475f
C189 source.n16 a_n1992_n1288# 0.04373f
C190 source.n17 a_n1992_n1288# 0.096758f
C191 source.t22 a_n1992_n1288# 0.072612f
C192 source.n18 a_n1992_n1288# 0.075727f
C193 source.n19 a_n1992_n1288# 0.024411f
C194 source.n20 a_n1992_n1288# 0.0161f
C195 source.n21 a_n1992_n1288# 0.213278f
C196 source.n22 a_n1992_n1288# 0.047938f
C197 source.n23 a_n1992_n1288# 0.118294f
C198 source.n24 a_n1992_n1288# 0.04373f
C199 source.n25 a_n1992_n1288# 0.096758f
C200 source.t0 a_n1992_n1288# 0.072612f
C201 source.n26 a_n1992_n1288# 0.075727f
C202 source.n27 a_n1992_n1288# 0.024411f
C203 source.n28 a_n1992_n1288# 0.0161f
C204 source.n29 a_n1992_n1288# 0.213278f
C205 source.n30 a_n1992_n1288# 0.047938f
C206 source.n31 a_n1992_n1288# 0.118294f
C207 source.t5 a_n1992_n1288# 0.047352f
C208 source.t9 a_n1992_n1288# 0.047352f
C209 source.n32 a_n1992_n1288# 0.253144f
C210 source.n33 a_n1992_n1288# 0.329475f
C211 source.t38 a_n1992_n1288# 0.047352f
C212 source.t15 a_n1992_n1288# 0.047352f
C213 source.n34 a_n1992_n1288# 0.253144f
C214 source.n35 a_n1992_n1288# 0.329475f
C215 source.t13 a_n1992_n1288# 0.047352f
C216 source.t6 a_n1992_n1288# 0.047352f
C217 source.n36 a_n1992_n1288# 0.253144f
C218 source.n37 a_n1992_n1288# 0.329475f
C219 source.t7 a_n1992_n1288# 0.047352f
C220 source.t2 a_n1992_n1288# 0.047352f
C221 source.n38 a_n1992_n1288# 0.253144f
C222 source.n39 a_n1992_n1288# 0.329475f
C223 source.n40 a_n1992_n1288# 0.04373f
C224 source.n41 a_n1992_n1288# 0.096758f
C225 source.t11 a_n1992_n1288# 0.072612f
C226 source.n42 a_n1992_n1288# 0.075727f
C227 source.n43 a_n1992_n1288# 0.024411f
C228 source.n44 a_n1992_n1288# 0.0161f
C229 source.n45 a_n1992_n1288# 0.213278f
C230 source.n46 a_n1992_n1288# 0.047938f
C231 source.n47 a_n1992_n1288# 0.723369f
C232 source.n48 a_n1992_n1288# 0.04373f
C233 source.n49 a_n1992_n1288# 0.096758f
C234 source.t34 a_n1992_n1288# 0.072612f
C235 source.n50 a_n1992_n1288# 0.075727f
C236 source.n51 a_n1992_n1288# 0.024411f
C237 source.n52 a_n1992_n1288# 0.0161f
C238 source.n53 a_n1992_n1288# 0.213278f
C239 source.n54 a_n1992_n1288# 0.047938f
C240 source.n55 a_n1992_n1288# 0.723369f
C241 source.t29 a_n1992_n1288# 0.047352f
C242 source.t20 a_n1992_n1288# 0.047352f
C243 source.n56 a_n1992_n1288# 0.253142f
C244 source.n57 a_n1992_n1288# 0.329476f
C245 source.t19 a_n1992_n1288# 0.047352f
C246 source.t36 a_n1992_n1288# 0.047352f
C247 source.n58 a_n1992_n1288# 0.253142f
C248 source.n59 a_n1992_n1288# 0.329476f
C249 source.t35 a_n1992_n1288# 0.047352f
C250 source.t30 a_n1992_n1288# 0.047352f
C251 source.n60 a_n1992_n1288# 0.253142f
C252 source.n61 a_n1992_n1288# 0.329476f
C253 source.t32 a_n1992_n1288# 0.047352f
C254 source.t18 a_n1992_n1288# 0.047352f
C255 source.n62 a_n1992_n1288# 0.253142f
C256 source.n63 a_n1992_n1288# 0.329476f
C257 source.n64 a_n1992_n1288# 0.04373f
C258 source.n65 a_n1992_n1288# 0.096758f
C259 source.t28 a_n1992_n1288# 0.072612f
C260 source.n66 a_n1992_n1288# 0.075727f
C261 source.n67 a_n1992_n1288# 0.024411f
C262 source.n68 a_n1992_n1288# 0.0161f
C263 source.n69 a_n1992_n1288# 0.213278f
C264 source.n70 a_n1992_n1288# 0.047938f
C265 source.n71 a_n1992_n1288# 0.118294f
C266 source.n72 a_n1992_n1288# 0.04373f
C267 source.n73 a_n1992_n1288# 0.096758f
C268 source.t39 a_n1992_n1288# 0.072612f
C269 source.n74 a_n1992_n1288# 0.075727f
C270 source.n75 a_n1992_n1288# 0.024411f
C271 source.n76 a_n1992_n1288# 0.0161f
C272 source.n77 a_n1992_n1288# 0.213278f
C273 source.n78 a_n1992_n1288# 0.047938f
C274 source.n79 a_n1992_n1288# 0.118294f
C275 source.t8 a_n1992_n1288# 0.047352f
C276 source.t16 a_n1992_n1288# 0.047352f
C277 source.n80 a_n1992_n1288# 0.253142f
C278 source.n81 a_n1992_n1288# 0.329476f
C279 source.t10 a_n1992_n1288# 0.047352f
C280 source.t3 a_n1992_n1288# 0.047352f
C281 source.n82 a_n1992_n1288# 0.253142f
C282 source.n83 a_n1992_n1288# 0.329476f
C283 source.t17 a_n1992_n1288# 0.047352f
C284 source.t14 a_n1992_n1288# 0.047352f
C285 source.n84 a_n1992_n1288# 0.253142f
C286 source.n85 a_n1992_n1288# 0.329476f
C287 source.t4 a_n1992_n1288# 0.047352f
C288 source.t1 a_n1992_n1288# 0.047352f
C289 source.n86 a_n1992_n1288# 0.253142f
C290 source.n87 a_n1992_n1288# 0.329476f
C291 source.n88 a_n1992_n1288# 0.04373f
C292 source.n89 a_n1992_n1288# 0.096758f
C293 source.t12 a_n1992_n1288# 0.072612f
C294 source.n90 a_n1992_n1288# 0.075727f
C295 source.n91 a_n1992_n1288# 0.024411f
C296 source.n92 a_n1992_n1288# 0.0161f
C297 source.n93 a_n1992_n1288# 0.213278f
C298 source.n94 a_n1992_n1288# 0.047938f
C299 source.n95 a_n1992_n1288# 0.284092f
C300 source.n96 a_n1992_n1288# 0.73899f
C301 plus.n0 a_n1992_n1288# 0.027601f
C302 plus.t14 a_n1992_n1288# 0.040609f
C303 plus.t5 a_n1992_n1288# 0.040609f
C304 plus.t11 a_n1992_n1288# 0.040609f
C305 plus.n1 a_n1992_n1288# 0.02978f
C306 plus.n2 a_n1992_n1288# 0.027601f
C307 plus.t18 a_n1992_n1288# 0.040609f
C308 plus.t12 a_n1992_n1288# 0.040609f
C309 plus.n3 a_n1992_n1288# 0.02978f
C310 plus.n4 a_n1992_n1288# 0.027601f
C311 plus.t0 a_n1992_n1288# 0.040609f
C312 plus.t13 a_n1992_n1288# 0.040609f
C313 plus.t1 a_n1992_n1288# 0.040609f
C314 plus.n5 a_n1992_n1288# 0.02978f
C315 plus.t8 a_n1992_n1288# 0.045099f
C316 plus.n6 a_n1992_n1288# 0.037721f
C317 plus.n7 a_n1992_n1288# 0.063158f
C318 plus.n8 a_n1992_n1288# 0.010517f
C319 plus.n9 a_n1992_n1288# 0.02978f
C320 plus.n10 a_n1992_n1288# 0.010517f
C321 plus.n11 a_n1992_n1288# 0.02978f
C322 plus.n12 a_n1992_n1288# 0.010517f
C323 plus.n13 a_n1992_n1288# 0.027601f
C324 plus.n14 a_n1992_n1288# 0.027601f
C325 plus.n15 a_n1992_n1288# 0.009837f
C326 plus.n16 a_n1992_n1288# 0.009837f
C327 plus.n17 a_n1992_n1288# 0.02978f
C328 plus.n18 a_n1992_n1288# 0.010517f
C329 plus.n19 a_n1992_n1288# 0.027601f
C330 plus.n20 a_n1992_n1288# 0.027601f
C331 plus.n21 a_n1992_n1288# 0.010517f
C332 plus.n22 a_n1992_n1288# 0.02978f
C333 plus.n23 a_n1992_n1288# 0.010517f
C334 plus.n24 a_n1992_n1288# 0.02978f
C335 plus.t4 a_n1992_n1288# 0.045099f
C336 plus.n25 a_n1992_n1288# 0.03768f
C337 plus.n26 a_n1992_n1288# 0.19709f
C338 plus.n27 a_n1992_n1288# 0.027601f
C339 plus.t9 a_n1992_n1288# 0.045099f
C340 plus.t10 a_n1992_n1288# 0.040609f
C341 plus.t6 a_n1992_n1288# 0.040609f
C342 plus.t19 a_n1992_n1288# 0.040609f
C343 plus.n28 a_n1992_n1288# 0.02978f
C344 plus.n29 a_n1992_n1288# 0.027601f
C345 plus.t3 a_n1992_n1288# 0.040609f
C346 plus.t16 a_n1992_n1288# 0.040609f
C347 plus.n30 a_n1992_n1288# 0.02978f
C348 plus.n31 a_n1992_n1288# 0.027601f
C349 plus.t7 a_n1992_n1288# 0.040609f
C350 plus.t2 a_n1992_n1288# 0.040609f
C351 plus.t15 a_n1992_n1288# 0.040609f
C352 plus.n32 a_n1992_n1288# 0.02978f
C353 plus.t17 a_n1992_n1288# 0.045099f
C354 plus.n33 a_n1992_n1288# 0.037721f
C355 plus.n34 a_n1992_n1288# 0.063158f
C356 plus.n35 a_n1992_n1288# 0.010517f
C357 plus.n36 a_n1992_n1288# 0.02978f
C358 plus.n37 a_n1992_n1288# 0.010517f
C359 plus.n38 a_n1992_n1288# 0.02978f
C360 plus.n39 a_n1992_n1288# 0.010517f
C361 plus.n40 a_n1992_n1288# 0.027601f
C362 plus.n41 a_n1992_n1288# 0.027601f
C363 plus.n42 a_n1992_n1288# 0.009837f
C364 plus.n43 a_n1992_n1288# 0.009837f
C365 plus.n44 a_n1992_n1288# 0.02978f
C366 plus.n45 a_n1992_n1288# 0.010517f
C367 plus.n46 a_n1992_n1288# 0.027601f
C368 plus.n47 a_n1992_n1288# 0.027601f
C369 plus.n48 a_n1992_n1288# 0.010517f
C370 plus.n49 a_n1992_n1288# 0.02978f
C371 plus.n50 a_n1992_n1288# 0.010517f
C372 plus.n51 a_n1992_n1288# 0.02978f
C373 plus.n52 a_n1992_n1288# 0.03768f
C374 plus.n53 a_n1992_n1288# 0.649184f
.ends

