* NGSPICE file created from diffpair263.ext - technology: sky130A

.subckt diffpair263 minus drain_right drain_left source plus
X0 a_n1296_n2088# a_n1296_n2088# a_n1296_n2088# a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.25
X1 drain_left.t7 plus.t0 source.t12 a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X2 drain_left.t6 plus.t1 source.t7 a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X3 drain_left.t5 plus.t2 source.t13 a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X4 source.t4 minus.t0 drain_right.t7 a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X5 source.t0 minus.t1 drain_right.t6 a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X6 source.t14 plus.t3 drain_left.t4 a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X7 drain_right.t5 minus.t2 source.t15 a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X8 a_n1296_n2088# a_n1296_n2088# a_n1296_n2088# a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X9 source.t8 plus.t4 drain_left.t3 a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X10 source.t2 minus.t3 drain_right.t4 a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X11 source.t9 plus.t5 drain_left.t2 a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X12 drain_left.t1 plus.t6 source.t10 a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X13 drain_right.t3 minus.t4 source.t1 a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X14 source.t5 minus.t5 drain_right.t2 a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X15 drain_right.t1 minus.t6 source.t6 a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X16 source.t11 plus.t7 drain_left.t0 a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X17 a_n1296_n2088# a_n1296_n2088# a_n1296_n2088# a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X18 drain_right.t0 minus.t7 source.t3 a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X19 a_n1296_n2088# a_n1296_n2088# a_n1296_n2088# a_n1296_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
R0 plus.n1 plus.t3 757.763
R1 plus.n5 plus.t0 757.763
R2 plus.n8 plus.t6 757.763
R3 plus.n12 plus.t7 757.763
R4 plus.n2 plus.t1 703.721
R5 plus.n4 plus.t5 703.721
R6 plus.n9 plus.t4 703.721
R7 plus.n11 plus.t2 703.721
R8 plus.n1 plus.n0 161.489
R9 plus.n8 plus.n7 161.489
R10 plus.n3 plus.n0 161.3
R11 plus.n6 plus.n5 161.3
R12 plus.n10 plus.n7 161.3
R13 plus.n13 plus.n12 161.3
R14 plus.n3 plus.n2 42.3581
R15 plus.n4 plus.n3 42.3581
R16 plus.n11 plus.n10 42.3581
R17 plus.n10 plus.n9 42.3581
R18 plus.n2 plus.n1 30.6732
R19 plus.n5 plus.n4 30.6732
R20 plus.n12 plus.n11 30.6732
R21 plus.n9 plus.n8 30.6732
R22 plus plus.n13 25.6392
R23 plus plus.n6 9.87171
R24 plus.n6 plus.n0 0.189894
R25 plus.n13 plus.n7 0.189894
R26 source.n258 source.n232 289.615
R27 source.n224 source.n198 289.615
R28 source.n192 source.n166 289.615
R29 source.n158 source.n132 289.615
R30 source.n26 source.n0 289.615
R31 source.n60 source.n34 289.615
R32 source.n92 source.n66 289.615
R33 source.n126 source.n100 289.615
R34 source.n243 source.n242 185
R35 source.n240 source.n239 185
R36 source.n249 source.n248 185
R37 source.n251 source.n250 185
R38 source.n236 source.n235 185
R39 source.n257 source.n256 185
R40 source.n259 source.n258 185
R41 source.n209 source.n208 185
R42 source.n206 source.n205 185
R43 source.n215 source.n214 185
R44 source.n217 source.n216 185
R45 source.n202 source.n201 185
R46 source.n223 source.n222 185
R47 source.n225 source.n224 185
R48 source.n177 source.n176 185
R49 source.n174 source.n173 185
R50 source.n183 source.n182 185
R51 source.n185 source.n184 185
R52 source.n170 source.n169 185
R53 source.n191 source.n190 185
R54 source.n193 source.n192 185
R55 source.n143 source.n142 185
R56 source.n140 source.n139 185
R57 source.n149 source.n148 185
R58 source.n151 source.n150 185
R59 source.n136 source.n135 185
R60 source.n157 source.n156 185
R61 source.n159 source.n158 185
R62 source.n27 source.n26 185
R63 source.n25 source.n24 185
R64 source.n4 source.n3 185
R65 source.n19 source.n18 185
R66 source.n17 source.n16 185
R67 source.n8 source.n7 185
R68 source.n11 source.n10 185
R69 source.n61 source.n60 185
R70 source.n59 source.n58 185
R71 source.n38 source.n37 185
R72 source.n53 source.n52 185
R73 source.n51 source.n50 185
R74 source.n42 source.n41 185
R75 source.n45 source.n44 185
R76 source.n93 source.n92 185
R77 source.n91 source.n90 185
R78 source.n70 source.n69 185
R79 source.n85 source.n84 185
R80 source.n83 source.n82 185
R81 source.n74 source.n73 185
R82 source.n77 source.n76 185
R83 source.n127 source.n126 185
R84 source.n125 source.n124 185
R85 source.n104 source.n103 185
R86 source.n119 source.n118 185
R87 source.n117 source.n116 185
R88 source.n108 source.n107 185
R89 source.n111 source.n110 185
R90 source.t15 source.n241 147.661
R91 source.t5 source.n207 147.661
R92 source.t10 source.n175 147.661
R93 source.t11 source.n141 147.661
R94 source.t12 source.n9 147.661
R95 source.t14 source.n43 147.661
R96 source.t6 source.n75 147.661
R97 source.t4 source.n109 147.661
R98 source.n242 source.n239 104.615
R99 source.n249 source.n239 104.615
R100 source.n250 source.n249 104.615
R101 source.n250 source.n235 104.615
R102 source.n257 source.n235 104.615
R103 source.n258 source.n257 104.615
R104 source.n208 source.n205 104.615
R105 source.n215 source.n205 104.615
R106 source.n216 source.n215 104.615
R107 source.n216 source.n201 104.615
R108 source.n223 source.n201 104.615
R109 source.n224 source.n223 104.615
R110 source.n176 source.n173 104.615
R111 source.n183 source.n173 104.615
R112 source.n184 source.n183 104.615
R113 source.n184 source.n169 104.615
R114 source.n191 source.n169 104.615
R115 source.n192 source.n191 104.615
R116 source.n142 source.n139 104.615
R117 source.n149 source.n139 104.615
R118 source.n150 source.n149 104.615
R119 source.n150 source.n135 104.615
R120 source.n157 source.n135 104.615
R121 source.n158 source.n157 104.615
R122 source.n26 source.n25 104.615
R123 source.n25 source.n3 104.615
R124 source.n18 source.n3 104.615
R125 source.n18 source.n17 104.615
R126 source.n17 source.n7 104.615
R127 source.n10 source.n7 104.615
R128 source.n60 source.n59 104.615
R129 source.n59 source.n37 104.615
R130 source.n52 source.n37 104.615
R131 source.n52 source.n51 104.615
R132 source.n51 source.n41 104.615
R133 source.n44 source.n41 104.615
R134 source.n92 source.n91 104.615
R135 source.n91 source.n69 104.615
R136 source.n84 source.n69 104.615
R137 source.n84 source.n83 104.615
R138 source.n83 source.n73 104.615
R139 source.n76 source.n73 104.615
R140 source.n126 source.n125 104.615
R141 source.n125 source.n103 104.615
R142 source.n118 source.n103 104.615
R143 source.n118 source.n117 104.615
R144 source.n117 source.n107 104.615
R145 source.n110 source.n107 104.615
R146 source.n242 source.t15 52.3082
R147 source.n208 source.t5 52.3082
R148 source.n176 source.t10 52.3082
R149 source.n142 source.t11 52.3082
R150 source.n10 source.t12 52.3082
R151 source.n44 source.t14 52.3082
R152 source.n76 source.t6 52.3082
R153 source.n110 source.t4 52.3082
R154 source.n33 source.n32 50.512
R155 source.n99 source.n98 50.512
R156 source.n231 source.n230 50.5119
R157 source.n165 source.n164 50.5119
R158 source.n263 source.n262 32.1853
R159 source.n229 source.n228 32.1853
R160 source.n197 source.n196 32.1853
R161 source.n163 source.n162 32.1853
R162 source.n31 source.n30 32.1853
R163 source.n65 source.n64 32.1853
R164 source.n97 source.n96 32.1853
R165 source.n131 source.n130 32.1853
R166 source.n163 source.n131 17.2423
R167 source.n243 source.n241 15.6674
R168 source.n209 source.n207 15.6674
R169 source.n177 source.n175 15.6674
R170 source.n143 source.n141 15.6674
R171 source.n11 source.n9 15.6674
R172 source.n45 source.n43 15.6674
R173 source.n77 source.n75 15.6674
R174 source.n111 source.n109 15.6674
R175 source.n244 source.n240 12.8005
R176 source.n210 source.n206 12.8005
R177 source.n178 source.n174 12.8005
R178 source.n144 source.n140 12.8005
R179 source.n12 source.n8 12.8005
R180 source.n46 source.n42 12.8005
R181 source.n78 source.n74 12.8005
R182 source.n112 source.n108 12.8005
R183 source.n248 source.n247 12.0247
R184 source.n214 source.n213 12.0247
R185 source.n182 source.n181 12.0247
R186 source.n148 source.n147 12.0247
R187 source.n16 source.n15 12.0247
R188 source.n50 source.n49 12.0247
R189 source.n82 source.n81 12.0247
R190 source.n116 source.n115 12.0247
R191 source.n264 source.n31 11.7293
R192 source.n251 source.n238 11.249
R193 source.n217 source.n204 11.249
R194 source.n185 source.n172 11.249
R195 source.n151 source.n138 11.249
R196 source.n19 source.n6 11.249
R197 source.n53 source.n40 11.249
R198 source.n85 source.n72 11.249
R199 source.n119 source.n106 11.249
R200 source.n252 source.n236 10.4732
R201 source.n218 source.n202 10.4732
R202 source.n186 source.n170 10.4732
R203 source.n152 source.n136 10.4732
R204 source.n20 source.n4 10.4732
R205 source.n54 source.n38 10.4732
R206 source.n86 source.n70 10.4732
R207 source.n120 source.n104 10.4732
R208 source.n256 source.n255 9.69747
R209 source.n222 source.n221 9.69747
R210 source.n190 source.n189 9.69747
R211 source.n156 source.n155 9.69747
R212 source.n24 source.n23 9.69747
R213 source.n58 source.n57 9.69747
R214 source.n90 source.n89 9.69747
R215 source.n124 source.n123 9.69747
R216 source.n262 source.n261 9.45567
R217 source.n228 source.n227 9.45567
R218 source.n196 source.n195 9.45567
R219 source.n162 source.n161 9.45567
R220 source.n30 source.n29 9.45567
R221 source.n64 source.n63 9.45567
R222 source.n96 source.n95 9.45567
R223 source.n130 source.n129 9.45567
R224 source.n261 source.n260 9.3005
R225 source.n234 source.n233 9.3005
R226 source.n255 source.n254 9.3005
R227 source.n253 source.n252 9.3005
R228 source.n238 source.n237 9.3005
R229 source.n247 source.n246 9.3005
R230 source.n245 source.n244 9.3005
R231 source.n227 source.n226 9.3005
R232 source.n200 source.n199 9.3005
R233 source.n221 source.n220 9.3005
R234 source.n219 source.n218 9.3005
R235 source.n204 source.n203 9.3005
R236 source.n213 source.n212 9.3005
R237 source.n211 source.n210 9.3005
R238 source.n195 source.n194 9.3005
R239 source.n168 source.n167 9.3005
R240 source.n189 source.n188 9.3005
R241 source.n187 source.n186 9.3005
R242 source.n172 source.n171 9.3005
R243 source.n181 source.n180 9.3005
R244 source.n179 source.n178 9.3005
R245 source.n161 source.n160 9.3005
R246 source.n134 source.n133 9.3005
R247 source.n155 source.n154 9.3005
R248 source.n153 source.n152 9.3005
R249 source.n138 source.n137 9.3005
R250 source.n147 source.n146 9.3005
R251 source.n145 source.n144 9.3005
R252 source.n29 source.n28 9.3005
R253 source.n2 source.n1 9.3005
R254 source.n23 source.n22 9.3005
R255 source.n21 source.n20 9.3005
R256 source.n6 source.n5 9.3005
R257 source.n15 source.n14 9.3005
R258 source.n13 source.n12 9.3005
R259 source.n63 source.n62 9.3005
R260 source.n36 source.n35 9.3005
R261 source.n57 source.n56 9.3005
R262 source.n55 source.n54 9.3005
R263 source.n40 source.n39 9.3005
R264 source.n49 source.n48 9.3005
R265 source.n47 source.n46 9.3005
R266 source.n95 source.n94 9.3005
R267 source.n68 source.n67 9.3005
R268 source.n89 source.n88 9.3005
R269 source.n87 source.n86 9.3005
R270 source.n72 source.n71 9.3005
R271 source.n81 source.n80 9.3005
R272 source.n79 source.n78 9.3005
R273 source.n129 source.n128 9.3005
R274 source.n102 source.n101 9.3005
R275 source.n123 source.n122 9.3005
R276 source.n121 source.n120 9.3005
R277 source.n106 source.n105 9.3005
R278 source.n115 source.n114 9.3005
R279 source.n113 source.n112 9.3005
R280 source.n259 source.n234 8.92171
R281 source.n225 source.n200 8.92171
R282 source.n193 source.n168 8.92171
R283 source.n159 source.n134 8.92171
R284 source.n27 source.n2 8.92171
R285 source.n61 source.n36 8.92171
R286 source.n93 source.n68 8.92171
R287 source.n127 source.n102 8.92171
R288 source.n260 source.n232 8.14595
R289 source.n226 source.n198 8.14595
R290 source.n194 source.n166 8.14595
R291 source.n160 source.n132 8.14595
R292 source.n28 source.n0 8.14595
R293 source.n62 source.n34 8.14595
R294 source.n94 source.n66 8.14595
R295 source.n128 source.n100 8.14595
R296 source.n262 source.n232 5.81868
R297 source.n228 source.n198 5.81868
R298 source.n196 source.n166 5.81868
R299 source.n162 source.n132 5.81868
R300 source.n30 source.n0 5.81868
R301 source.n64 source.n34 5.81868
R302 source.n96 source.n66 5.81868
R303 source.n130 source.n100 5.81868
R304 source.n264 source.n263 5.51343
R305 source.n260 source.n259 5.04292
R306 source.n226 source.n225 5.04292
R307 source.n194 source.n193 5.04292
R308 source.n160 source.n159 5.04292
R309 source.n28 source.n27 5.04292
R310 source.n62 source.n61 5.04292
R311 source.n94 source.n93 5.04292
R312 source.n128 source.n127 5.04292
R313 source.n245 source.n241 4.38594
R314 source.n211 source.n207 4.38594
R315 source.n179 source.n175 4.38594
R316 source.n145 source.n141 4.38594
R317 source.n13 source.n9 4.38594
R318 source.n47 source.n43 4.38594
R319 source.n79 source.n75 4.38594
R320 source.n113 source.n109 4.38594
R321 source.n256 source.n234 4.26717
R322 source.n222 source.n200 4.26717
R323 source.n190 source.n168 4.26717
R324 source.n156 source.n134 4.26717
R325 source.n24 source.n2 4.26717
R326 source.n58 source.n36 4.26717
R327 source.n90 source.n68 4.26717
R328 source.n124 source.n102 4.26717
R329 source.n255 source.n236 3.49141
R330 source.n221 source.n202 3.49141
R331 source.n189 source.n170 3.49141
R332 source.n155 source.n136 3.49141
R333 source.n23 source.n4 3.49141
R334 source.n57 source.n38 3.49141
R335 source.n89 source.n70 3.49141
R336 source.n123 source.n104 3.49141
R337 source.n230 source.t3 3.3005
R338 source.n230 source.t2 3.3005
R339 source.n164 source.t13 3.3005
R340 source.n164 source.t8 3.3005
R341 source.n32 source.t7 3.3005
R342 source.n32 source.t9 3.3005
R343 source.n98 source.t1 3.3005
R344 source.n98 source.t0 3.3005
R345 source.n252 source.n251 2.71565
R346 source.n218 source.n217 2.71565
R347 source.n186 source.n185 2.71565
R348 source.n152 source.n151 2.71565
R349 source.n20 source.n19 2.71565
R350 source.n54 source.n53 2.71565
R351 source.n86 source.n85 2.71565
R352 source.n120 source.n119 2.71565
R353 source.n248 source.n238 1.93989
R354 source.n214 source.n204 1.93989
R355 source.n182 source.n172 1.93989
R356 source.n148 source.n138 1.93989
R357 source.n16 source.n6 1.93989
R358 source.n50 source.n40 1.93989
R359 source.n82 source.n72 1.93989
R360 source.n116 source.n106 1.93989
R361 source.n247 source.n240 1.16414
R362 source.n213 source.n206 1.16414
R363 source.n181 source.n174 1.16414
R364 source.n147 source.n140 1.16414
R365 source.n15 source.n8 1.16414
R366 source.n49 source.n42 1.16414
R367 source.n81 source.n74 1.16414
R368 source.n115 source.n108 1.16414
R369 source.n131 source.n99 0.5005
R370 source.n99 source.n97 0.5005
R371 source.n65 source.n33 0.5005
R372 source.n33 source.n31 0.5005
R373 source.n165 source.n163 0.5005
R374 source.n197 source.n165 0.5005
R375 source.n231 source.n229 0.5005
R376 source.n263 source.n231 0.5005
R377 source.n97 source.n65 0.470328
R378 source.n229 source.n197 0.470328
R379 source.n244 source.n243 0.388379
R380 source.n210 source.n209 0.388379
R381 source.n178 source.n177 0.388379
R382 source.n144 source.n143 0.388379
R383 source.n12 source.n11 0.388379
R384 source.n46 source.n45 0.388379
R385 source.n78 source.n77 0.388379
R386 source.n112 source.n111 0.388379
R387 source source.n264 0.188
R388 source.n246 source.n245 0.155672
R389 source.n246 source.n237 0.155672
R390 source.n253 source.n237 0.155672
R391 source.n254 source.n253 0.155672
R392 source.n254 source.n233 0.155672
R393 source.n261 source.n233 0.155672
R394 source.n212 source.n211 0.155672
R395 source.n212 source.n203 0.155672
R396 source.n219 source.n203 0.155672
R397 source.n220 source.n219 0.155672
R398 source.n220 source.n199 0.155672
R399 source.n227 source.n199 0.155672
R400 source.n180 source.n179 0.155672
R401 source.n180 source.n171 0.155672
R402 source.n187 source.n171 0.155672
R403 source.n188 source.n187 0.155672
R404 source.n188 source.n167 0.155672
R405 source.n195 source.n167 0.155672
R406 source.n146 source.n145 0.155672
R407 source.n146 source.n137 0.155672
R408 source.n153 source.n137 0.155672
R409 source.n154 source.n153 0.155672
R410 source.n154 source.n133 0.155672
R411 source.n161 source.n133 0.155672
R412 source.n29 source.n1 0.155672
R413 source.n22 source.n1 0.155672
R414 source.n22 source.n21 0.155672
R415 source.n21 source.n5 0.155672
R416 source.n14 source.n5 0.155672
R417 source.n14 source.n13 0.155672
R418 source.n63 source.n35 0.155672
R419 source.n56 source.n35 0.155672
R420 source.n56 source.n55 0.155672
R421 source.n55 source.n39 0.155672
R422 source.n48 source.n39 0.155672
R423 source.n48 source.n47 0.155672
R424 source.n95 source.n67 0.155672
R425 source.n88 source.n67 0.155672
R426 source.n88 source.n87 0.155672
R427 source.n87 source.n71 0.155672
R428 source.n80 source.n71 0.155672
R429 source.n80 source.n79 0.155672
R430 source.n129 source.n101 0.155672
R431 source.n122 source.n101 0.155672
R432 source.n122 source.n121 0.155672
R433 source.n121 source.n105 0.155672
R434 source.n114 source.n105 0.155672
R435 source.n114 source.n113 0.155672
R436 drain_left.n5 drain_left.n3 67.6908
R437 drain_left.n2 drain_left.n1 67.3853
R438 drain_left.n2 drain_left.n0 67.3853
R439 drain_left.n5 drain_left.n4 67.1907
R440 drain_left drain_left.n2 24.5716
R441 drain_left drain_left.n5 6.15322
R442 drain_left.n1 drain_left.t3 3.3005
R443 drain_left.n1 drain_left.t1 3.3005
R444 drain_left.n0 drain_left.t0 3.3005
R445 drain_left.n0 drain_left.t5 3.3005
R446 drain_left.n4 drain_left.t2 3.3005
R447 drain_left.n4 drain_left.t7 3.3005
R448 drain_left.n3 drain_left.t4 3.3005
R449 drain_left.n3 drain_left.t6 3.3005
R450 minus.n5 minus.t0 757.763
R451 minus.n1 minus.t6 757.763
R452 minus.n12 minus.t2 757.763
R453 minus.n8 minus.t5 757.763
R454 minus.n4 minus.t4 703.721
R455 minus.n2 minus.t1 703.721
R456 minus.n11 minus.t3 703.721
R457 minus.n9 minus.t7 703.721
R458 minus.n1 minus.n0 161.489
R459 minus.n8 minus.n7 161.489
R460 minus.n6 minus.n5 161.3
R461 minus.n3 minus.n0 161.3
R462 minus.n13 minus.n12 161.3
R463 minus.n10 minus.n7 161.3
R464 minus.n4 minus.n3 42.3581
R465 minus.n3 minus.n2 42.3581
R466 minus.n10 minus.n9 42.3581
R467 minus.n11 minus.n10 42.3581
R468 minus.n5 minus.n4 30.6732
R469 minus.n2 minus.n1 30.6732
R470 minus.n9 minus.n8 30.6732
R471 minus.n12 minus.n11 30.6732
R472 minus.n14 minus.n6 29.4853
R473 minus.n14 minus.n13 6.5005
R474 minus.n6 minus.n0 0.189894
R475 minus.n13 minus.n7 0.189894
R476 minus minus.n14 0.188
R477 drain_right.n5 drain_right.n3 67.6907
R478 drain_right.n2 drain_right.n1 67.3853
R479 drain_right.n2 drain_right.n0 67.3853
R480 drain_right.n5 drain_right.n4 67.1908
R481 drain_right drain_right.n2 24.0184
R482 drain_right drain_right.n5 6.15322
R483 drain_right.n1 drain_right.t4 3.3005
R484 drain_right.n1 drain_right.t5 3.3005
R485 drain_right.n0 drain_right.t2 3.3005
R486 drain_right.n0 drain_right.t0 3.3005
R487 drain_right.n3 drain_right.t6 3.3005
R488 drain_right.n3 drain_right.t1 3.3005
R489 drain_right.n4 drain_right.t7 3.3005
R490 drain_right.n4 drain_right.t3 3.3005
C0 drain_right minus 1.67696f
C1 drain_left minus 0.170438f
C2 minus plus 3.65502f
C3 drain_right drain_left 0.605638f
C4 drain_right plus 0.275273f
C5 drain_left plus 1.79896f
C6 source minus 1.51727f
C7 source drain_right 9.862201f
C8 source drain_left 9.86333f
C9 source plus 1.53129f
C10 drain_right a_n1296_n2088# 4.10826f
C11 drain_left a_n1296_n2088# 4.27614f
C12 source a_n1296_n2088# 5.087322f
C13 minus a_n1296_n2088# 4.504012f
C14 plus a_n1296_n2088# 5.288948f
C15 drain_right.t2 a_n1296_n2088# 0.136737f
C16 drain_right.t0 a_n1296_n2088# 0.136737f
C17 drain_right.n0 a_n1296_n2088# 1.1413f
C18 drain_right.t4 a_n1296_n2088# 0.136737f
C19 drain_right.t5 a_n1296_n2088# 0.136737f
C20 drain_right.n1 a_n1296_n2088# 1.1413f
C21 drain_right.n2 a_n1296_n2088# 1.43781f
C22 drain_right.t6 a_n1296_n2088# 0.136737f
C23 drain_right.t1 a_n1296_n2088# 0.136737f
C24 drain_right.n3 a_n1296_n2088# 1.14289f
C25 drain_right.t7 a_n1296_n2088# 0.136737f
C26 drain_right.t3 a_n1296_n2088# 0.136737f
C27 drain_right.n4 a_n1296_n2088# 1.1404f
C28 drain_right.n5 a_n1296_n2088# 0.901146f
C29 minus.n0 a_n1296_n2088# 0.070285f
C30 minus.t0 a_n1296_n2088# 0.135115f
C31 minus.t4 a_n1296_n2088# 0.130567f
C32 minus.t1 a_n1296_n2088# 0.130567f
C33 minus.t6 a_n1296_n2088# 0.135115f
C34 minus.n1 a_n1296_n2088# 0.070903f
C35 minus.n2 a_n1296_n2088# 0.061502f
C36 minus.n3 a_n1296_n2088# 0.011642f
C37 minus.n4 a_n1296_n2088# 0.061502f
C38 minus.n5 a_n1296_n2088# 0.070857f
C39 minus.n6 a_n1296_n2088# 0.77153f
C40 minus.n7 a_n1296_n2088# 0.070285f
C41 minus.t3 a_n1296_n2088# 0.130567f
C42 minus.t7 a_n1296_n2088# 0.130567f
C43 minus.t5 a_n1296_n2088# 0.135115f
C44 minus.n8 a_n1296_n2088# 0.070903f
C45 minus.n9 a_n1296_n2088# 0.061502f
C46 minus.n10 a_n1296_n2088# 0.011642f
C47 minus.n11 a_n1296_n2088# 0.061502f
C48 minus.t2 a_n1296_n2088# 0.135115f
C49 minus.n12 a_n1296_n2088# 0.070857f
C50 minus.n13 a_n1296_n2088# 0.19977f
C51 minus.n14 a_n1296_n2088# 0.952532f
C52 drain_left.t0 a_n1296_n2088# 0.135197f
C53 drain_left.t5 a_n1296_n2088# 0.135197f
C54 drain_left.n0 a_n1296_n2088# 1.12844f
C55 drain_left.t3 a_n1296_n2088# 0.135197f
C56 drain_left.t1 a_n1296_n2088# 0.135197f
C57 drain_left.n1 a_n1296_n2088# 1.12844f
C58 drain_left.n2 a_n1296_n2088# 1.48005f
C59 drain_left.t4 a_n1296_n2088# 0.135197f
C60 drain_left.t6 a_n1296_n2088# 0.135197f
C61 drain_left.n3 a_n1296_n2088# 1.13002f
C62 drain_left.t2 a_n1296_n2088# 0.135197f
C63 drain_left.t7 a_n1296_n2088# 0.135197f
C64 drain_left.n4 a_n1296_n2088# 1.12754f
C65 drain_left.n5 a_n1296_n2088# 0.890993f
C66 source.n0 a_n1296_n2088# 0.03204f
C67 source.n1 a_n1296_n2088# 0.022795f
C68 source.n2 a_n1296_n2088# 0.012249f
C69 source.n3 a_n1296_n2088# 0.028952f
C70 source.n4 a_n1296_n2088# 0.012969f
C71 source.n5 a_n1296_n2088# 0.022795f
C72 source.n6 a_n1296_n2088# 0.012249f
C73 source.n7 a_n1296_n2088# 0.028952f
C74 source.n8 a_n1296_n2088# 0.012969f
C75 source.n9 a_n1296_n2088# 0.097545f
C76 source.t12 a_n1296_n2088# 0.047188f
C77 source.n10 a_n1296_n2088# 0.021714f
C78 source.n11 a_n1296_n2088# 0.017102f
C79 source.n12 a_n1296_n2088# 0.012249f
C80 source.n13 a_n1296_n2088# 0.542378f
C81 source.n14 a_n1296_n2088# 0.022795f
C82 source.n15 a_n1296_n2088# 0.012249f
C83 source.n16 a_n1296_n2088# 0.012969f
C84 source.n17 a_n1296_n2088# 0.028952f
C85 source.n18 a_n1296_n2088# 0.028952f
C86 source.n19 a_n1296_n2088# 0.012969f
C87 source.n20 a_n1296_n2088# 0.012249f
C88 source.n21 a_n1296_n2088# 0.022795f
C89 source.n22 a_n1296_n2088# 0.022795f
C90 source.n23 a_n1296_n2088# 0.012249f
C91 source.n24 a_n1296_n2088# 0.012969f
C92 source.n25 a_n1296_n2088# 0.028952f
C93 source.n26 a_n1296_n2088# 0.062676f
C94 source.n27 a_n1296_n2088# 0.012969f
C95 source.n28 a_n1296_n2088# 0.012249f
C96 source.n29 a_n1296_n2088# 0.052689f
C97 source.n30 a_n1296_n2088# 0.03507f
C98 source.n31 a_n1296_n2088# 0.546704f
C99 source.t7 a_n1296_n2088# 0.108078f
C100 source.t9 a_n1296_n2088# 0.108078f
C101 source.n32 a_n1296_n2088# 0.841723f
C102 source.n33 a_n1296_n2088# 0.287128f
C103 source.n34 a_n1296_n2088# 0.03204f
C104 source.n35 a_n1296_n2088# 0.022795f
C105 source.n36 a_n1296_n2088# 0.012249f
C106 source.n37 a_n1296_n2088# 0.028952f
C107 source.n38 a_n1296_n2088# 0.012969f
C108 source.n39 a_n1296_n2088# 0.022795f
C109 source.n40 a_n1296_n2088# 0.012249f
C110 source.n41 a_n1296_n2088# 0.028952f
C111 source.n42 a_n1296_n2088# 0.012969f
C112 source.n43 a_n1296_n2088# 0.097545f
C113 source.t14 a_n1296_n2088# 0.047188f
C114 source.n44 a_n1296_n2088# 0.021714f
C115 source.n45 a_n1296_n2088# 0.017102f
C116 source.n46 a_n1296_n2088# 0.012249f
C117 source.n47 a_n1296_n2088# 0.542378f
C118 source.n48 a_n1296_n2088# 0.022795f
C119 source.n49 a_n1296_n2088# 0.012249f
C120 source.n50 a_n1296_n2088# 0.012969f
C121 source.n51 a_n1296_n2088# 0.028952f
C122 source.n52 a_n1296_n2088# 0.028952f
C123 source.n53 a_n1296_n2088# 0.012969f
C124 source.n54 a_n1296_n2088# 0.012249f
C125 source.n55 a_n1296_n2088# 0.022795f
C126 source.n56 a_n1296_n2088# 0.022795f
C127 source.n57 a_n1296_n2088# 0.012249f
C128 source.n58 a_n1296_n2088# 0.012969f
C129 source.n59 a_n1296_n2088# 0.028952f
C130 source.n60 a_n1296_n2088# 0.062676f
C131 source.n61 a_n1296_n2088# 0.012969f
C132 source.n62 a_n1296_n2088# 0.012249f
C133 source.n63 a_n1296_n2088# 0.052689f
C134 source.n64 a_n1296_n2088# 0.03507f
C135 source.n65 a_n1296_n2088# 0.090702f
C136 source.n66 a_n1296_n2088# 0.03204f
C137 source.n67 a_n1296_n2088# 0.022795f
C138 source.n68 a_n1296_n2088# 0.012249f
C139 source.n69 a_n1296_n2088# 0.028952f
C140 source.n70 a_n1296_n2088# 0.012969f
C141 source.n71 a_n1296_n2088# 0.022795f
C142 source.n72 a_n1296_n2088# 0.012249f
C143 source.n73 a_n1296_n2088# 0.028952f
C144 source.n74 a_n1296_n2088# 0.012969f
C145 source.n75 a_n1296_n2088# 0.097545f
C146 source.t6 a_n1296_n2088# 0.047188f
C147 source.n76 a_n1296_n2088# 0.021714f
C148 source.n77 a_n1296_n2088# 0.017102f
C149 source.n78 a_n1296_n2088# 0.012249f
C150 source.n79 a_n1296_n2088# 0.542378f
C151 source.n80 a_n1296_n2088# 0.022795f
C152 source.n81 a_n1296_n2088# 0.012249f
C153 source.n82 a_n1296_n2088# 0.012969f
C154 source.n83 a_n1296_n2088# 0.028952f
C155 source.n84 a_n1296_n2088# 0.028952f
C156 source.n85 a_n1296_n2088# 0.012969f
C157 source.n86 a_n1296_n2088# 0.012249f
C158 source.n87 a_n1296_n2088# 0.022795f
C159 source.n88 a_n1296_n2088# 0.022795f
C160 source.n89 a_n1296_n2088# 0.012249f
C161 source.n90 a_n1296_n2088# 0.012969f
C162 source.n91 a_n1296_n2088# 0.028952f
C163 source.n92 a_n1296_n2088# 0.062676f
C164 source.n93 a_n1296_n2088# 0.012969f
C165 source.n94 a_n1296_n2088# 0.012249f
C166 source.n95 a_n1296_n2088# 0.052689f
C167 source.n96 a_n1296_n2088# 0.03507f
C168 source.n97 a_n1296_n2088# 0.090702f
C169 source.t1 a_n1296_n2088# 0.108078f
C170 source.t0 a_n1296_n2088# 0.108078f
C171 source.n98 a_n1296_n2088# 0.841723f
C172 source.n99 a_n1296_n2088# 0.287128f
C173 source.n100 a_n1296_n2088# 0.03204f
C174 source.n101 a_n1296_n2088# 0.022795f
C175 source.n102 a_n1296_n2088# 0.012249f
C176 source.n103 a_n1296_n2088# 0.028952f
C177 source.n104 a_n1296_n2088# 0.012969f
C178 source.n105 a_n1296_n2088# 0.022795f
C179 source.n106 a_n1296_n2088# 0.012249f
C180 source.n107 a_n1296_n2088# 0.028952f
C181 source.n108 a_n1296_n2088# 0.012969f
C182 source.n109 a_n1296_n2088# 0.097545f
C183 source.t4 a_n1296_n2088# 0.047188f
C184 source.n110 a_n1296_n2088# 0.021714f
C185 source.n111 a_n1296_n2088# 0.017102f
C186 source.n112 a_n1296_n2088# 0.012249f
C187 source.n113 a_n1296_n2088# 0.542378f
C188 source.n114 a_n1296_n2088# 0.022795f
C189 source.n115 a_n1296_n2088# 0.012249f
C190 source.n116 a_n1296_n2088# 0.012969f
C191 source.n117 a_n1296_n2088# 0.028952f
C192 source.n118 a_n1296_n2088# 0.028952f
C193 source.n119 a_n1296_n2088# 0.012969f
C194 source.n120 a_n1296_n2088# 0.012249f
C195 source.n121 a_n1296_n2088# 0.022795f
C196 source.n122 a_n1296_n2088# 0.022795f
C197 source.n123 a_n1296_n2088# 0.012249f
C198 source.n124 a_n1296_n2088# 0.012969f
C199 source.n125 a_n1296_n2088# 0.028952f
C200 source.n126 a_n1296_n2088# 0.062676f
C201 source.n127 a_n1296_n2088# 0.012969f
C202 source.n128 a_n1296_n2088# 0.012249f
C203 source.n129 a_n1296_n2088# 0.052689f
C204 source.n130 a_n1296_n2088# 0.03507f
C205 source.n131 a_n1296_n2088# 0.839259f
C206 source.n132 a_n1296_n2088# 0.03204f
C207 source.n133 a_n1296_n2088# 0.022795f
C208 source.n134 a_n1296_n2088# 0.012249f
C209 source.n135 a_n1296_n2088# 0.028952f
C210 source.n136 a_n1296_n2088# 0.012969f
C211 source.n137 a_n1296_n2088# 0.022795f
C212 source.n138 a_n1296_n2088# 0.012249f
C213 source.n139 a_n1296_n2088# 0.028952f
C214 source.n140 a_n1296_n2088# 0.012969f
C215 source.n141 a_n1296_n2088# 0.097545f
C216 source.t11 a_n1296_n2088# 0.047188f
C217 source.n142 a_n1296_n2088# 0.021714f
C218 source.n143 a_n1296_n2088# 0.017102f
C219 source.n144 a_n1296_n2088# 0.012249f
C220 source.n145 a_n1296_n2088# 0.542378f
C221 source.n146 a_n1296_n2088# 0.022795f
C222 source.n147 a_n1296_n2088# 0.012249f
C223 source.n148 a_n1296_n2088# 0.012969f
C224 source.n149 a_n1296_n2088# 0.028952f
C225 source.n150 a_n1296_n2088# 0.028952f
C226 source.n151 a_n1296_n2088# 0.012969f
C227 source.n152 a_n1296_n2088# 0.012249f
C228 source.n153 a_n1296_n2088# 0.022795f
C229 source.n154 a_n1296_n2088# 0.022795f
C230 source.n155 a_n1296_n2088# 0.012249f
C231 source.n156 a_n1296_n2088# 0.012969f
C232 source.n157 a_n1296_n2088# 0.028952f
C233 source.n158 a_n1296_n2088# 0.062676f
C234 source.n159 a_n1296_n2088# 0.012969f
C235 source.n160 a_n1296_n2088# 0.012249f
C236 source.n161 a_n1296_n2088# 0.052689f
C237 source.n162 a_n1296_n2088# 0.03507f
C238 source.n163 a_n1296_n2088# 0.839259f
C239 source.t13 a_n1296_n2088# 0.108078f
C240 source.t8 a_n1296_n2088# 0.108078f
C241 source.n164 a_n1296_n2088# 0.841718f
C242 source.n165 a_n1296_n2088# 0.287134f
C243 source.n166 a_n1296_n2088# 0.03204f
C244 source.n167 a_n1296_n2088# 0.022795f
C245 source.n168 a_n1296_n2088# 0.012249f
C246 source.n169 a_n1296_n2088# 0.028952f
C247 source.n170 a_n1296_n2088# 0.012969f
C248 source.n171 a_n1296_n2088# 0.022795f
C249 source.n172 a_n1296_n2088# 0.012249f
C250 source.n173 a_n1296_n2088# 0.028952f
C251 source.n174 a_n1296_n2088# 0.012969f
C252 source.n175 a_n1296_n2088# 0.097545f
C253 source.t10 a_n1296_n2088# 0.047188f
C254 source.n176 a_n1296_n2088# 0.021714f
C255 source.n177 a_n1296_n2088# 0.017102f
C256 source.n178 a_n1296_n2088# 0.012249f
C257 source.n179 a_n1296_n2088# 0.542378f
C258 source.n180 a_n1296_n2088# 0.022795f
C259 source.n181 a_n1296_n2088# 0.012249f
C260 source.n182 a_n1296_n2088# 0.012969f
C261 source.n183 a_n1296_n2088# 0.028952f
C262 source.n184 a_n1296_n2088# 0.028952f
C263 source.n185 a_n1296_n2088# 0.012969f
C264 source.n186 a_n1296_n2088# 0.012249f
C265 source.n187 a_n1296_n2088# 0.022795f
C266 source.n188 a_n1296_n2088# 0.022795f
C267 source.n189 a_n1296_n2088# 0.012249f
C268 source.n190 a_n1296_n2088# 0.012969f
C269 source.n191 a_n1296_n2088# 0.028952f
C270 source.n192 a_n1296_n2088# 0.062676f
C271 source.n193 a_n1296_n2088# 0.012969f
C272 source.n194 a_n1296_n2088# 0.012249f
C273 source.n195 a_n1296_n2088# 0.052689f
C274 source.n196 a_n1296_n2088# 0.03507f
C275 source.n197 a_n1296_n2088# 0.090702f
C276 source.n198 a_n1296_n2088# 0.03204f
C277 source.n199 a_n1296_n2088# 0.022795f
C278 source.n200 a_n1296_n2088# 0.012249f
C279 source.n201 a_n1296_n2088# 0.028952f
C280 source.n202 a_n1296_n2088# 0.012969f
C281 source.n203 a_n1296_n2088# 0.022795f
C282 source.n204 a_n1296_n2088# 0.012249f
C283 source.n205 a_n1296_n2088# 0.028952f
C284 source.n206 a_n1296_n2088# 0.012969f
C285 source.n207 a_n1296_n2088# 0.097545f
C286 source.t5 a_n1296_n2088# 0.047188f
C287 source.n208 a_n1296_n2088# 0.021714f
C288 source.n209 a_n1296_n2088# 0.017102f
C289 source.n210 a_n1296_n2088# 0.012249f
C290 source.n211 a_n1296_n2088# 0.542378f
C291 source.n212 a_n1296_n2088# 0.022795f
C292 source.n213 a_n1296_n2088# 0.012249f
C293 source.n214 a_n1296_n2088# 0.012969f
C294 source.n215 a_n1296_n2088# 0.028952f
C295 source.n216 a_n1296_n2088# 0.028952f
C296 source.n217 a_n1296_n2088# 0.012969f
C297 source.n218 a_n1296_n2088# 0.012249f
C298 source.n219 a_n1296_n2088# 0.022795f
C299 source.n220 a_n1296_n2088# 0.022795f
C300 source.n221 a_n1296_n2088# 0.012249f
C301 source.n222 a_n1296_n2088# 0.012969f
C302 source.n223 a_n1296_n2088# 0.028952f
C303 source.n224 a_n1296_n2088# 0.062676f
C304 source.n225 a_n1296_n2088# 0.012969f
C305 source.n226 a_n1296_n2088# 0.012249f
C306 source.n227 a_n1296_n2088# 0.052689f
C307 source.n228 a_n1296_n2088# 0.03507f
C308 source.n229 a_n1296_n2088# 0.090702f
C309 source.t3 a_n1296_n2088# 0.108078f
C310 source.t2 a_n1296_n2088# 0.108078f
C311 source.n230 a_n1296_n2088# 0.841718f
C312 source.n231 a_n1296_n2088# 0.287134f
C313 source.n232 a_n1296_n2088# 0.03204f
C314 source.n233 a_n1296_n2088# 0.022795f
C315 source.n234 a_n1296_n2088# 0.012249f
C316 source.n235 a_n1296_n2088# 0.028952f
C317 source.n236 a_n1296_n2088# 0.012969f
C318 source.n237 a_n1296_n2088# 0.022795f
C319 source.n238 a_n1296_n2088# 0.012249f
C320 source.n239 a_n1296_n2088# 0.028952f
C321 source.n240 a_n1296_n2088# 0.012969f
C322 source.n241 a_n1296_n2088# 0.097545f
C323 source.t15 a_n1296_n2088# 0.047188f
C324 source.n242 a_n1296_n2088# 0.021714f
C325 source.n243 a_n1296_n2088# 0.017102f
C326 source.n244 a_n1296_n2088# 0.012249f
C327 source.n245 a_n1296_n2088# 0.542378f
C328 source.n246 a_n1296_n2088# 0.022795f
C329 source.n247 a_n1296_n2088# 0.012249f
C330 source.n248 a_n1296_n2088# 0.012969f
C331 source.n249 a_n1296_n2088# 0.028952f
C332 source.n250 a_n1296_n2088# 0.028952f
C333 source.n251 a_n1296_n2088# 0.012969f
C334 source.n252 a_n1296_n2088# 0.012249f
C335 source.n253 a_n1296_n2088# 0.022795f
C336 source.n254 a_n1296_n2088# 0.022795f
C337 source.n255 a_n1296_n2088# 0.012249f
C338 source.n256 a_n1296_n2088# 0.012969f
C339 source.n257 a_n1296_n2088# 0.028952f
C340 source.n258 a_n1296_n2088# 0.062676f
C341 source.n259 a_n1296_n2088# 0.012969f
C342 source.n260 a_n1296_n2088# 0.012249f
C343 source.n261 a_n1296_n2088# 0.052689f
C344 source.n262 a_n1296_n2088# 0.03507f
C345 source.n263 a_n1296_n2088# 0.216844f
C346 source.n264 a_n1296_n2088# 0.931185f
C347 plus.n0 a_n1296_n2088# 0.071478f
C348 plus.t5 a_n1296_n2088# 0.132784f
C349 plus.t1 a_n1296_n2088# 0.132784f
C350 plus.t3 a_n1296_n2088# 0.137409f
C351 plus.n1 a_n1296_n2088# 0.072107f
C352 plus.n2 a_n1296_n2088# 0.062546f
C353 plus.n3 a_n1296_n2088# 0.011839f
C354 plus.n4 a_n1296_n2088# 0.062546f
C355 plus.t0 a_n1296_n2088# 0.137409f
C356 plus.n5 a_n1296_n2088# 0.07206f
C357 plus.n6 a_n1296_n2088# 0.266272f
C358 plus.n7 a_n1296_n2088# 0.071478f
C359 plus.t7 a_n1296_n2088# 0.137409f
C360 plus.t2 a_n1296_n2088# 0.132784f
C361 plus.t4 a_n1296_n2088# 0.132784f
C362 plus.t6 a_n1296_n2088# 0.137409f
C363 plus.n8 a_n1296_n2088# 0.072107f
C364 plus.n9 a_n1296_n2088# 0.062546f
C365 plus.n10 a_n1296_n2088# 0.011839f
C366 plus.n11 a_n1296_n2088# 0.062546f
C367 plus.n12 a_n1296_n2088# 0.07206f
C368 plus.n13 a_n1296_n2088# 0.709762f
.ends

