* NGSPICE file created from diffpair422.ext - technology: sky130A

.subckt diffpair422 minus drain_right drain_left source plus
X0 source.t11 plus.t0 drain_left.t2 a_n1180_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X1 source.t1 minus.t0 drain_right.t5 a_n1180_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X2 source.t4 minus.t1 drain_right.t4 a_n1180_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X3 drain_left.t1 plus.t1 source.t10 a_n1180_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X4 drain_left.t3 plus.t2 source.t9 a_n1180_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X5 drain_left.t4 plus.t3 source.t8 a_n1180_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X6 a_n1180_n3288# a_n1180_n3288# a_n1180_n3288# a_n1180_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.25
X7 a_n1180_n3288# a_n1180_n3288# a_n1180_n3288# a_n1180_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X8 a_n1180_n3288# a_n1180_n3288# a_n1180_n3288# a_n1180_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X9 drain_right.t3 minus.t2 source.t3 a_n1180_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
X10 drain_right.t2 minus.t3 source.t5 a_n1180_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X11 source.t7 plus.t4 drain_left.t0 a_n1180_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.25
X12 drain_right.t1 minus.t4 source.t2 a_n1180_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X13 drain_left.t5 plus.t5 source.t6 a_n1180_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.25
X14 a_n1180_n3288# a_n1180_n3288# a_n1180_n3288# a_n1180_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.25
X15 drain_right.t0 minus.t5 source.t0 a_n1180_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.25
R0 plus.n0 plus.t1 1330.32
R1 plus.n2 plus.t3 1330.32
R2 plus.n4 plus.t5 1330.32
R3 plus.n6 plus.t2 1330.32
R4 plus.n1 plus.t0 1282.12
R5 plus.n5 plus.t4 1282.12
R6 plus.n3 plus.n0 161.489
R7 plus.n7 plus.n4 161.489
R8 plus.n3 plus.n2 161.3
R9 plus.n7 plus.n6 161.3
R10 plus.n1 plus.n0 36.5157
R11 plus.n2 plus.n1 36.5157
R12 plus.n6 plus.n5 36.5157
R13 plus.n5 plus.n4 36.5157
R14 plus plus.n7 27.4574
R15 plus plus.n3 12.1293
R16 drain_left.n60 drain_left.n0 289.615
R17 drain_left.n127 drain_left.n67 289.615
R18 drain_left.n20 drain_left.n19 185
R19 drain_left.n25 drain_left.n24 185
R20 drain_left.n27 drain_left.n26 185
R21 drain_left.n16 drain_left.n15 185
R22 drain_left.n33 drain_left.n32 185
R23 drain_left.n35 drain_left.n34 185
R24 drain_left.n12 drain_left.n11 185
R25 drain_left.n42 drain_left.n41 185
R26 drain_left.n43 drain_left.n10 185
R27 drain_left.n45 drain_left.n44 185
R28 drain_left.n8 drain_left.n7 185
R29 drain_left.n51 drain_left.n50 185
R30 drain_left.n53 drain_left.n52 185
R31 drain_left.n4 drain_left.n3 185
R32 drain_left.n59 drain_left.n58 185
R33 drain_left.n61 drain_left.n60 185
R34 drain_left.n128 drain_left.n127 185
R35 drain_left.n126 drain_left.n125 185
R36 drain_left.n71 drain_left.n70 185
R37 drain_left.n120 drain_left.n119 185
R38 drain_left.n118 drain_left.n117 185
R39 drain_left.n75 drain_left.n74 185
R40 drain_left.n112 drain_left.n111 185
R41 drain_left.n110 drain_left.n77 185
R42 drain_left.n109 drain_left.n108 185
R43 drain_left.n80 drain_left.n78 185
R44 drain_left.n103 drain_left.n102 185
R45 drain_left.n101 drain_left.n100 185
R46 drain_left.n84 drain_left.n83 185
R47 drain_left.n95 drain_left.n94 185
R48 drain_left.n93 drain_left.n92 185
R49 drain_left.n88 drain_left.n87 185
R50 drain_left.n21 drain_left.t3 149.524
R51 drain_left.n89 drain_left.t1 149.524
R52 drain_left.n25 drain_left.n19 104.615
R53 drain_left.n26 drain_left.n25 104.615
R54 drain_left.n26 drain_left.n15 104.615
R55 drain_left.n33 drain_left.n15 104.615
R56 drain_left.n34 drain_left.n33 104.615
R57 drain_left.n34 drain_left.n11 104.615
R58 drain_left.n42 drain_left.n11 104.615
R59 drain_left.n43 drain_left.n42 104.615
R60 drain_left.n44 drain_left.n43 104.615
R61 drain_left.n44 drain_left.n7 104.615
R62 drain_left.n51 drain_left.n7 104.615
R63 drain_left.n52 drain_left.n51 104.615
R64 drain_left.n52 drain_left.n3 104.615
R65 drain_left.n59 drain_left.n3 104.615
R66 drain_left.n60 drain_left.n59 104.615
R67 drain_left.n127 drain_left.n126 104.615
R68 drain_left.n126 drain_left.n70 104.615
R69 drain_left.n119 drain_left.n70 104.615
R70 drain_left.n119 drain_left.n118 104.615
R71 drain_left.n118 drain_left.n74 104.615
R72 drain_left.n111 drain_left.n74 104.615
R73 drain_left.n111 drain_left.n110 104.615
R74 drain_left.n110 drain_left.n109 104.615
R75 drain_left.n109 drain_left.n78 104.615
R76 drain_left.n102 drain_left.n78 104.615
R77 drain_left.n102 drain_left.n101 104.615
R78 drain_left.n101 drain_left.n83 104.615
R79 drain_left.n94 drain_left.n83 104.615
R80 drain_left.n94 drain_left.n93 104.615
R81 drain_left.n93 drain_left.n87 104.615
R82 drain_left.n66 drain_left.n65 59.6222
R83 drain_left.n133 drain_left.n132 59.5525
R84 drain_left.t3 drain_left.n19 52.3082
R85 drain_left.t1 drain_left.n87 52.3082
R86 drain_left.n133 drain_left.n131 47.0369
R87 drain_left.n66 drain_left.n64 46.8565
R88 drain_left drain_left.n66 28.7421
R89 drain_left.n45 drain_left.n10 13.1884
R90 drain_left.n112 drain_left.n77 13.1884
R91 drain_left.n41 drain_left.n40 12.8005
R92 drain_left.n46 drain_left.n8 12.8005
R93 drain_left.n113 drain_left.n75 12.8005
R94 drain_left.n108 drain_left.n79 12.8005
R95 drain_left.n39 drain_left.n12 12.0247
R96 drain_left.n50 drain_left.n49 12.0247
R97 drain_left.n117 drain_left.n116 12.0247
R98 drain_left.n107 drain_left.n80 12.0247
R99 drain_left.n36 drain_left.n35 11.249
R100 drain_left.n53 drain_left.n6 11.249
R101 drain_left.n120 drain_left.n73 11.249
R102 drain_left.n104 drain_left.n103 11.249
R103 drain_left.n32 drain_left.n14 10.4732
R104 drain_left.n54 drain_left.n4 10.4732
R105 drain_left.n121 drain_left.n71 10.4732
R106 drain_left.n100 drain_left.n82 10.4732
R107 drain_left.n21 drain_left.n20 10.2747
R108 drain_left.n89 drain_left.n88 10.2747
R109 drain_left.n31 drain_left.n16 9.69747
R110 drain_left.n58 drain_left.n57 9.69747
R111 drain_left.n125 drain_left.n124 9.69747
R112 drain_left.n99 drain_left.n84 9.69747
R113 drain_left.n64 drain_left.n63 9.45567
R114 drain_left.n131 drain_left.n130 9.45567
R115 drain_left.n63 drain_left.n62 9.3005
R116 drain_left.n2 drain_left.n1 9.3005
R117 drain_left.n57 drain_left.n56 9.3005
R118 drain_left.n55 drain_left.n54 9.3005
R119 drain_left.n6 drain_left.n5 9.3005
R120 drain_left.n49 drain_left.n48 9.3005
R121 drain_left.n47 drain_left.n46 9.3005
R122 drain_left.n23 drain_left.n22 9.3005
R123 drain_left.n18 drain_left.n17 9.3005
R124 drain_left.n29 drain_left.n28 9.3005
R125 drain_left.n31 drain_left.n30 9.3005
R126 drain_left.n14 drain_left.n13 9.3005
R127 drain_left.n37 drain_left.n36 9.3005
R128 drain_left.n39 drain_left.n38 9.3005
R129 drain_left.n40 drain_left.n9 9.3005
R130 drain_left.n91 drain_left.n90 9.3005
R131 drain_left.n86 drain_left.n85 9.3005
R132 drain_left.n97 drain_left.n96 9.3005
R133 drain_left.n99 drain_left.n98 9.3005
R134 drain_left.n82 drain_left.n81 9.3005
R135 drain_left.n105 drain_left.n104 9.3005
R136 drain_left.n107 drain_left.n106 9.3005
R137 drain_left.n79 drain_left.n76 9.3005
R138 drain_left.n130 drain_left.n129 9.3005
R139 drain_left.n69 drain_left.n68 9.3005
R140 drain_left.n124 drain_left.n123 9.3005
R141 drain_left.n122 drain_left.n121 9.3005
R142 drain_left.n73 drain_left.n72 9.3005
R143 drain_left.n116 drain_left.n115 9.3005
R144 drain_left.n114 drain_left.n113 9.3005
R145 drain_left.n28 drain_left.n27 8.92171
R146 drain_left.n61 drain_left.n2 8.92171
R147 drain_left.n128 drain_left.n69 8.92171
R148 drain_left.n96 drain_left.n95 8.92171
R149 drain_left.n24 drain_left.n18 8.14595
R150 drain_left.n62 drain_left.n0 8.14595
R151 drain_left.n129 drain_left.n67 8.14595
R152 drain_left.n92 drain_left.n86 8.14595
R153 drain_left.n23 drain_left.n20 7.3702
R154 drain_left.n91 drain_left.n88 7.3702
R155 drain_left drain_left.n133 6.15322
R156 drain_left.n24 drain_left.n23 5.81868
R157 drain_left.n64 drain_left.n0 5.81868
R158 drain_left.n131 drain_left.n67 5.81868
R159 drain_left.n92 drain_left.n91 5.81868
R160 drain_left.n27 drain_left.n18 5.04292
R161 drain_left.n62 drain_left.n61 5.04292
R162 drain_left.n129 drain_left.n128 5.04292
R163 drain_left.n95 drain_left.n86 5.04292
R164 drain_left.n28 drain_left.n16 4.26717
R165 drain_left.n58 drain_left.n2 4.26717
R166 drain_left.n125 drain_left.n69 4.26717
R167 drain_left.n96 drain_left.n84 4.26717
R168 drain_left.n32 drain_left.n31 3.49141
R169 drain_left.n57 drain_left.n4 3.49141
R170 drain_left.n124 drain_left.n71 3.49141
R171 drain_left.n100 drain_left.n99 3.49141
R172 drain_left.n22 drain_left.n21 2.84303
R173 drain_left.n90 drain_left.n89 2.84303
R174 drain_left.n35 drain_left.n14 2.71565
R175 drain_left.n54 drain_left.n53 2.71565
R176 drain_left.n121 drain_left.n120 2.71565
R177 drain_left.n103 drain_left.n82 2.71565
R178 drain_left.n36 drain_left.n12 1.93989
R179 drain_left.n50 drain_left.n6 1.93989
R180 drain_left.n117 drain_left.n73 1.93989
R181 drain_left.n104 drain_left.n80 1.93989
R182 drain_left.n65 drain_left.t0 1.6505
R183 drain_left.n65 drain_left.t5 1.6505
R184 drain_left.n132 drain_left.t2 1.6505
R185 drain_left.n132 drain_left.t4 1.6505
R186 drain_left.n41 drain_left.n39 1.16414
R187 drain_left.n49 drain_left.n8 1.16414
R188 drain_left.n116 drain_left.n75 1.16414
R189 drain_left.n108 drain_left.n107 1.16414
R190 drain_left.n40 drain_left.n10 0.388379
R191 drain_left.n46 drain_left.n45 0.388379
R192 drain_left.n113 drain_left.n112 0.388379
R193 drain_left.n79 drain_left.n77 0.388379
R194 drain_left.n22 drain_left.n17 0.155672
R195 drain_left.n29 drain_left.n17 0.155672
R196 drain_left.n30 drain_left.n29 0.155672
R197 drain_left.n30 drain_left.n13 0.155672
R198 drain_left.n37 drain_left.n13 0.155672
R199 drain_left.n38 drain_left.n37 0.155672
R200 drain_left.n38 drain_left.n9 0.155672
R201 drain_left.n47 drain_left.n9 0.155672
R202 drain_left.n48 drain_left.n47 0.155672
R203 drain_left.n48 drain_left.n5 0.155672
R204 drain_left.n55 drain_left.n5 0.155672
R205 drain_left.n56 drain_left.n55 0.155672
R206 drain_left.n56 drain_left.n1 0.155672
R207 drain_left.n63 drain_left.n1 0.155672
R208 drain_left.n130 drain_left.n68 0.155672
R209 drain_left.n123 drain_left.n68 0.155672
R210 drain_left.n123 drain_left.n122 0.155672
R211 drain_left.n122 drain_left.n72 0.155672
R212 drain_left.n115 drain_left.n72 0.155672
R213 drain_left.n115 drain_left.n114 0.155672
R214 drain_left.n114 drain_left.n76 0.155672
R215 drain_left.n106 drain_left.n76 0.155672
R216 drain_left.n106 drain_left.n105 0.155672
R217 drain_left.n105 drain_left.n81 0.155672
R218 drain_left.n98 drain_left.n81 0.155672
R219 drain_left.n98 drain_left.n97 0.155672
R220 drain_left.n97 drain_left.n85 0.155672
R221 drain_left.n90 drain_left.n85 0.155672
R222 source.n266 source.n206 289.615
R223 source.n198 source.n138 289.615
R224 source.n60 source.n0 289.615
R225 source.n128 source.n68 289.615
R226 source.n226 source.n225 185
R227 source.n231 source.n230 185
R228 source.n233 source.n232 185
R229 source.n222 source.n221 185
R230 source.n239 source.n238 185
R231 source.n241 source.n240 185
R232 source.n218 source.n217 185
R233 source.n248 source.n247 185
R234 source.n249 source.n216 185
R235 source.n251 source.n250 185
R236 source.n214 source.n213 185
R237 source.n257 source.n256 185
R238 source.n259 source.n258 185
R239 source.n210 source.n209 185
R240 source.n265 source.n264 185
R241 source.n267 source.n266 185
R242 source.n158 source.n157 185
R243 source.n163 source.n162 185
R244 source.n165 source.n164 185
R245 source.n154 source.n153 185
R246 source.n171 source.n170 185
R247 source.n173 source.n172 185
R248 source.n150 source.n149 185
R249 source.n180 source.n179 185
R250 source.n181 source.n148 185
R251 source.n183 source.n182 185
R252 source.n146 source.n145 185
R253 source.n189 source.n188 185
R254 source.n191 source.n190 185
R255 source.n142 source.n141 185
R256 source.n197 source.n196 185
R257 source.n199 source.n198 185
R258 source.n61 source.n60 185
R259 source.n59 source.n58 185
R260 source.n4 source.n3 185
R261 source.n53 source.n52 185
R262 source.n51 source.n50 185
R263 source.n8 source.n7 185
R264 source.n45 source.n44 185
R265 source.n43 source.n10 185
R266 source.n42 source.n41 185
R267 source.n13 source.n11 185
R268 source.n36 source.n35 185
R269 source.n34 source.n33 185
R270 source.n17 source.n16 185
R271 source.n28 source.n27 185
R272 source.n26 source.n25 185
R273 source.n21 source.n20 185
R274 source.n129 source.n128 185
R275 source.n127 source.n126 185
R276 source.n72 source.n71 185
R277 source.n121 source.n120 185
R278 source.n119 source.n118 185
R279 source.n76 source.n75 185
R280 source.n113 source.n112 185
R281 source.n111 source.n78 185
R282 source.n110 source.n109 185
R283 source.n81 source.n79 185
R284 source.n104 source.n103 185
R285 source.n102 source.n101 185
R286 source.n85 source.n84 185
R287 source.n96 source.n95 185
R288 source.n94 source.n93 185
R289 source.n89 source.n88 185
R290 source.n227 source.t2 149.524
R291 source.n159 source.t6 149.524
R292 source.n22 source.t8 149.524
R293 source.n90 source.t5 149.524
R294 source.n231 source.n225 104.615
R295 source.n232 source.n231 104.615
R296 source.n232 source.n221 104.615
R297 source.n239 source.n221 104.615
R298 source.n240 source.n239 104.615
R299 source.n240 source.n217 104.615
R300 source.n248 source.n217 104.615
R301 source.n249 source.n248 104.615
R302 source.n250 source.n249 104.615
R303 source.n250 source.n213 104.615
R304 source.n257 source.n213 104.615
R305 source.n258 source.n257 104.615
R306 source.n258 source.n209 104.615
R307 source.n265 source.n209 104.615
R308 source.n266 source.n265 104.615
R309 source.n163 source.n157 104.615
R310 source.n164 source.n163 104.615
R311 source.n164 source.n153 104.615
R312 source.n171 source.n153 104.615
R313 source.n172 source.n171 104.615
R314 source.n172 source.n149 104.615
R315 source.n180 source.n149 104.615
R316 source.n181 source.n180 104.615
R317 source.n182 source.n181 104.615
R318 source.n182 source.n145 104.615
R319 source.n189 source.n145 104.615
R320 source.n190 source.n189 104.615
R321 source.n190 source.n141 104.615
R322 source.n197 source.n141 104.615
R323 source.n198 source.n197 104.615
R324 source.n60 source.n59 104.615
R325 source.n59 source.n3 104.615
R326 source.n52 source.n3 104.615
R327 source.n52 source.n51 104.615
R328 source.n51 source.n7 104.615
R329 source.n44 source.n7 104.615
R330 source.n44 source.n43 104.615
R331 source.n43 source.n42 104.615
R332 source.n42 source.n11 104.615
R333 source.n35 source.n11 104.615
R334 source.n35 source.n34 104.615
R335 source.n34 source.n16 104.615
R336 source.n27 source.n16 104.615
R337 source.n27 source.n26 104.615
R338 source.n26 source.n20 104.615
R339 source.n128 source.n127 104.615
R340 source.n127 source.n71 104.615
R341 source.n120 source.n71 104.615
R342 source.n120 source.n119 104.615
R343 source.n119 source.n75 104.615
R344 source.n112 source.n75 104.615
R345 source.n112 source.n111 104.615
R346 source.n111 source.n110 104.615
R347 source.n110 source.n79 104.615
R348 source.n103 source.n79 104.615
R349 source.n103 source.n102 104.615
R350 source.n102 source.n84 104.615
R351 source.n95 source.n84 104.615
R352 source.n95 source.n94 104.615
R353 source.n94 source.n88 104.615
R354 source.t2 source.n225 52.3082
R355 source.t6 source.n157 52.3082
R356 source.t8 source.n20 52.3082
R357 source.t5 source.n88 52.3082
R358 source.n67 source.n66 42.8739
R359 source.n135 source.n134 42.8739
R360 source.n205 source.n204 42.8737
R361 source.n137 source.n136 42.8737
R362 source.n271 source.n270 29.8581
R363 source.n203 source.n202 29.8581
R364 source.n65 source.n64 29.8581
R365 source.n133 source.n132 29.8581
R366 source.n137 source.n135 22.2877
R367 source.n272 source.n65 16.2748
R368 source.n251 source.n216 13.1884
R369 source.n183 source.n148 13.1884
R370 source.n45 source.n10 13.1884
R371 source.n113 source.n78 13.1884
R372 source.n247 source.n246 12.8005
R373 source.n252 source.n214 12.8005
R374 source.n179 source.n178 12.8005
R375 source.n184 source.n146 12.8005
R376 source.n46 source.n8 12.8005
R377 source.n41 source.n12 12.8005
R378 source.n114 source.n76 12.8005
R379 source.n109 source.n80 12.8005
R380 source.n245 source.n218 12.0247
R381 source.n256 source.n255 12.0247
R382 source.n177 source.n150 12.0247
R383 source.n188 source.n187 12.0247
R384 source.n50 source.n49 12.0247
R385 source.n40 source.n13 12.0247
R386 source.n118 source.n117 12.0247
R387 source.n108 source.n81 12.0247
R388 source.n242 source.n241 11.249
R389 source.n259 source.n212 11.249
R390 source.n174 source.n173 11.249
R391 source.n191 source.n144 11.249
R392 source.n53 source.n6 11.249
R393 source.n37 source.n36 11.249
R394 source.n121 source.n74 11.249
R395 source.n105 source.n104 11.249
R396 source.n238 source.n220 10.4732
R397 source.n260 source.n210 10.4732
R398 source.n170 source.n152 10.4732
R399 source.n192 source.n142 10.4732
R400 source.n54 source.n4 10.4732
R401 source.n33 source.n15 10.4732
R402 source.n122 source.n72 10.4732
R403 source.n101 source.n83 10.4732
R404 source.n227 source.n226 10.2747
R405 source.n159 source.n158 10.2747
R406 source.n22 source.n21 10.2747
R407 source.n90 source.n89 10.2747
R408 source.n237 source.n222 9.69747
R409 source.n264 source.n263 9.69747
R410 source.n169 source.n154 9.69747
R411 source.n196 source.n195 9.69747
R412 source.n58 source.n57 9.69747
R413 source.n32 source.n17 9.69747
R414 source.n126 source.n125 9.69747
R415 source.n100 source.n85 9.69747
R416 source.n270 source.n269 9.45567
R417 source.n202 source.n201 9.45567
R418 source.n64 source.n63 9.45567
R419 source.n132 source.n131 9.45567
R420 source.n269 source.n268 9.3005
R421 source.n208 source.n207 9.3005
R422 source.n263 source.n262 9.3005
R423 source.n261 source.n260 9.3005
R424 source.n212 source.n211 9.3005
R425 source.n255 source.n254 9.3005
R426 source.n253 source.n252 9.3005
R427 source.n229 source.n228 9.3005
R428 source.n224 source.n223 9.3005
R429 source.n235 source.n234 9.3005
R430 source.n237 source.n236 9.3005
R431 source.n220 source.n219 9.3005
R432 source.n243 source.n242 9.3005
R433 source.n245 source.n244 9.3005
R434 source.n246 source.n215 9.3005
R435 source.n201 source.n200 9.3005
R436 source.n140 source.n139 9.3005
R437 source.n195 source.n194 9.3005
R438 source.n193 source.n192 9.3005
R439 source.n144 source.n143 9.3005
R440 source.n187 source.n186 9.3005
R441 source.n185 source.n184 9.3005
R442 source.n161 source.n160 9.3005
R443 source.n156 source.n155 9.3005
R444 source.n167 source.n166 9.3005
R445 source.n169 source.n168 9.3005
R446 source.n152 source.n151 9.3005
R447 source.n175 source.n174 9.3005
R448 source.n177 source.n176 9.3005
R449 source.n178 source.n147 9.3005
R450 source.n24 source.n23 9.3005
R451 source.n19 source.n18 9.3005
R452 source.n30 source.n29 9.3005
R453 source.n32 source.n31 9.3005
R454 source.n15 source.n14 9.3005
R455 source.n38 source.n37 9.3005
R456 source.n40 source.n39 9.3005
R457 source.n12 source.n9 9.3005
R458 source.n63 source.n62 9.3005
R459 source.n2 source.n1 9.3005
R460 source.n57 source.n56 9.3005
R461 source.n55 source.n54 9.3005
R462 source.n6 source.n5 9.3005
R463 source.n49 source.n48 9.3005
R464 source.n47 source.n46 9.3005
R465 source.n92 source.n91 9.3005
R466 source.n87 source.n86 9.3005
R467 source.n98 source.n97 9.3005
R468 source.n100 source.n99 9.3005
R469 source.n83 source.n82 9.3005
R470 source.n106 source.n105 9.3005
R471 source.n108 source.n107 9.3005
R472 source.n80 source.n77 9.3005
R473 source.n131 source.n130 9.3005
R474 source.n70 source.n69 9.3005
R475 source.n125 source.n124 9.3005
R476 source.n123 source.n122 9.3005
R477 source.n74 source.n73 9.3005
R478 source.n117 source.n116 9.3005
R479 source.n115 source.n114 9.3005
R480 source.n234 source.n233 8.92171
R481 source.n267 source.n208 8.92171
R482 source.n166 source.n165 8.92171
R483 source.n199 source.n140 8.92171
R484 source.n61 source.n2 8.92171
R485 source.n29 source.n28 8.92171
R486 source.n129 source.n70 8.92171
R487 source.n97 source.n96 8.92171
R488 source.n230 source.n224 8.14595
R489 source.n268 source.n206 8.14595
R490 source.n162 source.n156 8.14595
R491 source.n200 source.n138 8.14595
R492 source.n62 source.n0 8.14595
R493 source.n25 source.n19 8.14595
R494 source.n130 source.n68 8.14595
R495 source.n93 source.n87 8.14595
R496 source.n229 source.n226 7.3702
R497 source.n161 source.n158 7.3702
R498 source.n24 source.n21 7.3702
R499 source.n92 source.n89 7.3702
R500 source.n230 source.n229 5.81868
R501 source.n270 source.n206 5.81868
R502 source.n162 source.n161 5.81868
R503 source.n202 source.n138 5.81868
R504 source.n64 source.n0 5.81868
R505 source.n25 source.n24 5.81868
R506 source.n132 source.n68 5.81868
R507 source.n93 source.n92 5.81868
R508 source.n272 source.n271 5.51343
R509 source.n233 source.n224 5.04292
R510 source.n268 source.n267 5.04292
R511 source.n165 source.n156 5.04292
R512 source.n200 source.n199 5.04292
R513 source.n62 source.n61 5.04292
R514 source.n28 source.n19 5.04292
R515 source.n130 source.n129 5.04292
R516 source.n96 source.n87 5.04292
R517 source.n234 source.n222 4.26717
R518 source.n264 source.n208 4.26717
R519 source.n166 source.n154 4.26717
R520 source.n196 source.n140 4.26717
R521 source.n58 source.n2 4.26717
R522 source.n29 source.n17 4.26717
R523 source.n126 source.n70 4.26717
R524 source.n97 source.n85 4.26717
R525 source.n238 source.n237 3.49141
R526 source.n263 source.n210 3.49141
R527 source.n170 source.n169 3.49141
R528 source.n195 source.n142 3.49141
R529 source.n57 source.n4 3.49141
R530 source.n33 source.n32 3.49141
R531 source.n125 source.n72 3.49141
R532 source.n101 source.n100 3.49141
R533 source.n228 source.n227 2.84303
R534 source.n160 source.n159 2.84303
R535 source.n23 source.n22 2.84303
R536 source.n91 source.n90 2.84303
R537 source.n241 source.n220 2.71565
R538 source.n260 source.n259 2.71565
R539 source.n173 source.n152 2.71565
R540 source.n192 source.n191 2.71565
R541 source.n54 source.n53 2.71565
R542 source.n36 source.n15 2.71565
R543 source.n122 source.n121 2.71565
R544 source.n104 source.n83 2.71565
R545 source.n242 source.n218 1.93989
R546 source.n256 source.n212 1.93989
R547 source.n174 source.n150 1.93989
R548 source.n188 source.n144 1.93989
R549 source.n50 source.n6 1.93989
R550 source.n37 source.n13 1.93989
R551 source.n118 source.n74 1.93989
R552 source.n105 source.n81 1.93989
R553 source.n204 source.t0 1.6505
R554 source.n204 source.t4 1.6505
R555 source.n136 source.t9 1.6505
R556 source.n136 source.t7 1.6505
R557 source.n66 source.t10 1.6505
R558 source.n66 source.t11 1.6505
R559 source.n134 source.t3 1.6505
R560 source.n134 source.t1 1.6505
R561 source.n247 source.n245 1.16414
R562 source.n255 source.n214 1.16414
R563 source.n179 source.n177 1.16414
R564 source.n187 source.n146 1.16414
R565 source.n49 source.n8 1.16414
R566 source.n41 source.n40 1.16414
R567 source.n117 source.n76 1.16414
R568 source.n109 source.n108 1.16414
R569 source.n133 source.n67 0.720328
R570 source.n205 source.n203 0.720328
R571 source.n135 source.n133 0.5005
R572 source.n67 source.n65 0.5005
R573 source.n203 source.n137 0.5005
R574 source.n271 source.n205 0.5005
R575 source.n246 source.n216 0.388379
R576 source.n252 source.n251 0.388379
R577 source.n178 source.n148 0.388379
R578 source.n184 source.n183 0.388379
R579 source.n46 source.n45 0.388379
R580 source.n12 source.n10 0.388379
R581 source.n114 source.n113 0.388379
R582 source.n80 source.n78 0.388379
R583 source source.n272 0.188
R584 source.n228 source.n223 0.155672
R585 source.n235 source.n223 0.155672
R586 source.n236 source.n235 0.155672
R587 source.n236 source.n219 0.155672
R588 source.n243 source.n219 0.155672
R589 source.n244 source.n243 0.155672
R590 source.n244 source.n215 0.155672
R591 source.n253 source.n215 0.155672
R592 source.n254 source.n253 0.155672
R593 source.n254 source.n211 0.155672
R594 source.n261 source.n211 0.155672
R595 source.n262 source.n261 0.155672
R596 source.n262 source.n207 0.155672
R597 source.n269 source.n207 0.155672
R598 source.n160 source.n155 0.155672
R599 source.n167 source.n155 0.155672
R600 source.n168 source.n167 0.155672
R601 source.n168 source.n151 0.155672
R602 source.n175 source.n151 0.155672
R603 source.n176 source.n175 0.155672
R604 source.n176 source.n147 0.155672
R605 source.n185 source.n147 0.155672
R606 source.n186 source.n185 0.155672
R607 source.n186 source.n143 0.155672
R608 source.n193 source.n143 0.155672
R609 source.n194 source.n193 0.155672
R610 source.n194 source.n139 0.155672
R611 source.n201 source.n139 0.155672
R612 source.n63 source.n1 0.155672
R613 source.n56 source.n1 0.155672
R614 source.n56 source.n55 0.155672
R615 source.n55 source.n5 0.155672
R616 source.n48 source.n5 0.155672
R617 source.n48 source.n47 0.155672
R618 source.n47 source.n9 0.155672
R619 source.n39 source.n9 0.155672
R620 source.n39 source.n38 0.155672
R621 source.n38 source.n14 0.155672
R622 source.n31 source.n14 0.155672
R623 source.n31 source.n30 0.155672
R624 source.n30 source.n18 0.155672
R625 source.n23 source.n18 0.155672
R626 source.n131 source.n69 0.155672
R627 source.n124 source.n69 0.155672
R628 source.n124 source.n123 0.155672
R629 source.n123 source.n73 0.155672
R630 source.n116 source.n73 0.155672
R631 source.n116 source.n115 0.155672
R632 source.n115 source.n77 0.155672
R633 source.n107 source.n77 0.155672
R634 source.n107 source.n106 0.155672
R635 source.n106 source.n82 0.155672
R636 source.n99 source.n82 0.155672
R637 source.n99 source.n98 0.155672
R638 source.n98 source.n86 0.155672
R639 source.n91 source.n86 0.155672
R640 minus.n2 minus.t2 1330.32
R641 minus.n0 minus.t3 1330.32
R642 minus.n6 minus.t4 1330.32
R643 minus.n4 minus.t5 1330.32
R644 minus.n1 minus.t0 1282.12
R645 minus.n5 minus.t1 1282.12
R646 minus.n3 minus.n0 161.489
R647 minus.n7 minus.n4 161.489
R648 minus.n3 minus.n2 161.3
R649 minus.n7 minus.n6 161.3
R650 minus.n2 minus.n1 36.5157
R651 minus.n1 minus.n0 36.5157
R652 minus.n5 minus.n4 36.5157
R653 minus.n6 minus.n5 36.5157
R654 minus.n8 minus.n3 33.5763
R655 minus.n8 minus.n7 6.48535
R656 minus minus.n8 0.188
R657 drain_right.n60 drain_right.n0 289.615
R658 drain_right.n128 drain_right.n68 289.615
R659 drain_right.n20 drain_right.n19 185
R660 drain_right.n25 drain_right.n24 185
R661 drain_right.n27 drain_right.n26 185
R662 drain_right.n16 drain_right.n15 185
R663 drain_right.n33 drain_right.n32 185
R664 drain_right.n35 drain_right.n34 185
R665 drain_right.n12 drain_right.n11 185
R666 drain_right.n42 drain_right.n41 185
R667 drain_right.n43 drain_right.n10 185
R668 drain_right.n45 drain_right.n44 185
R669 drain_right.n8 drain_right.n7 185
R670 drain_right.n51 drain_right.n50 185
R671 drain_right.n53 drain_right.n52 185
R672 drain_right.n4 drain_right.n3 185
R673 drain_right.n59 drain_right.n58 185
R674 drain_right.n61 drain_right.n60 185
R675 drain_right.n129 drain_right.n128 185
R676 drain_right.n127 drain_right.n126 185
R677 drain_right.n72 drain_right.n71 185
R678 drain_right.n121 drain_right.n120 185
R679 drain_right.n119 drain_right.n118 185
R680 drain_right.n76 drain_right.n75 185
R681 drain_right.n113 drain_right.n112 185
R682 drain_right.n111 drain_right.n78 185
R683 drain_right.n110 drain_right.n109 185
R684 drain_right.n81 drain_right.n79 185
R685 drain_right.n104 drain_right.n103 185
R686 drain_right.n102 drain_right.n101 185
R687 drain_right.n85 drain_right.n84 185
R688 drain_right.n96 drain_right.n95 185
R689 drain_right.n94 drain_right.n93 185
R690 drain_right.n89 drain_right.n88 185
R691 drain_right.n21 drain_right.t0 149.524
R692 drain_right.n90 drain_right.t3 149.524
R693 drain_right.n25 drain_right.n19 104.615
R694 drain_right.n26 drain_right.n25 104.615
R695 drain_right.n26 drain_right.n15 104.615
R696 drain_right.n33 drain_right.n15 104.615
R697 drain_right.n34 drain_right.n33 104.615
R698 drain_right.n34 drain_right.n11 104.615
R699 drain_right.n42 drain_right.n11 104.615
R700 drain_right.n43 drain_right.n42 104.615
R701 drain_right.n44 drain_right.n43 104.615
R702 drain_right.n44 drain_right.n7 104.615
R703 drain_right.n51 drain_right.n7 104.615
R704 drain_right.n52 drain_right.n51 104.615
R705 drain_right.n52 drain_right.n3 104.615
R706 drain_right.n59 drain_right.n3 104.615
R707 drain_right.n60 drain_right.n59 104.615
R708 drain_right.n128 drain_right.n127 104.615
R709 drain_right.n127 drain_right.n71 104.615
R710 drain_right.n120 drain_right.n71 104.615
R711 drain_right.n120 drain_right.n119 104.615
R712 drain_right.n119 drain_right.n75 104.615
R713 drain_right.n112 drain_right.n75 104.615
R714 drain_right.n112 drain_right.n111 104.615
R715 drain_right.n111 drain_right.n110 104.615
R716 drain_right.n110 drain_right.n79 104.615
R717 drain_right.n103 drain_right.n79 104.615
R718 drain_right.n103 drain_right.n102 104.615
R719 drain_right.n102 drain_right.n84 104.615
R720 drain_right.n95 drain_right.n84 104.615
R721 drain_right.n95 drain_right.n94 104.615
R722 drain_right.n94 drain_right.n88 104.615
R723 drain_right.n133 drain_right.n67 60.0525
R724 drain_right.n66 drain_right.n65 59.6222
R725 drain_right.t0 drain_right.n19 52.3082
R726 drain_right.t3 drain_right.n88 52.3082
R727 drain_right.n66 drain_right.n64 46.8565
R728 drain_right.n133 drain_right.n132 46.5369
R729 drain_right drain_right.n66 28.1888
R730 drain_right.n45 drain_right.n10 13.1884
R731 drain_right.n113 drain_right.n78 13.1884
R732 drain_right.n41 drain_right.n40 12.8005
R733 drain_right.n46 drain_right.n8 12.8005
R734 drain_right.n114 drain_right.n76 12.8005
R735 drain_right.n109 drain_right.n80 12.8005
R736 drain_right.n39 drain_right.n12 12.0247
R737 drain_right.n50 drain_right.n49 12.0247
R738 drain_right.n118 drain_right.n117 12.0247
R739 drain_right.n108 drain_right.n81 12.0247
R740 drain_right.n36 drain_right.n35 11.249
R741 drain_right.n53 drain_right.n6 11.249
R742 drain_right.n121 drain_right.n74 11.249
R743 drain_right.n105 drain_right.n104 11.249
R744 drain_right.n32 drain_right.n14 10.4732
R745 drain_right.n54 drain_right.n4 10.4732
R746 drain_right.n122 drain_right.n72 10.4732
R747 drain_right.n101 drain_right.n83 10.4732
R748 drain_right.n21 drain_right.n20 10.2747
R749 drain_right.n90 drain_right.n89 10.2747
R750 drain_right.n31 drain_right.n16 9.69747
R751 drain_right.n58 drain_right.n57 9.69747
R752 drain_right.n126 drain_right.n125 9.69747
R753 drain_right.n100 drain_right.n85 9.69747
R754 drain_right.n64 drain_right.n63 9.45567
R755 drain_right.n132 drain_right.n131 9.45567
R756 drain_right.n63 drain_right.n62 9.3005
R757 drain_right.n2 drain_right.n1 9.3005
R758 drain_right.n57 drain_right.n56 9.3005
R759 drain_right.n55 drain_right.n54 9.3005
R760 drain_right.n6 drain_right.n5 9.3005
R761 drain_right.n49 drain_right.n48 9.3005
R762 drain_right.n47 drain_right.n46 9.3005
R763 drain_right.n23 drain_right.n22 9.3005
R764 drain_right.n18 drain_right.n17 9.3005
R765 drain_right.n29 drain_right.n28 9.3005
R766 drain_right.n31 drain_right.n30 9.3005
R767 drain_right.n14 drain_right.n13 9.3005
R768 drain_right.n37 drain_right.n36 9.3005
R769 drain_right.n39 drain_right.n38 9.3005
R770 drain_right.n40 drain_right.n9 9.3005
R771 drain_right.n92 drain_right.n91 9.3005
R772 drain_right.n87 drain_right.n86 9.3005
R773 drain_right.n98 drain_right.n97 9.3005
R774 drain_right.n100 drain_right.n99 9.3005
R775 drain_right.n83 drain_right.n82 9.3005
R776 drain_right.n106 drain_right.n105 9.3005
R777 drain_right.n108 drain_right.n107 9.3005
R778 drain_right.n80 drain_right.n77 9.3005
R779 drain_right.n131 drain_right.n130 9.3005
R780 drain_right.n70 drain_right.n69 9.3005
R781 drain_right.n125 drain_right.n124 9.3005
R782 drain_right.n123 drain_right.n122 9.3005
R783 drain_right.n74 drain_right.n73 9.3005
R784 drain_right.n117 drain_right.n116 9.3005
R785 drain_right.n115 drain_right.n114 9.3005
R786 drain_right.n28 drain_right.n27 8.92171
R787 drain_right.n61 drain_right.n2 8.92171
R788 drain_right.n129 drain_right.n70 8.92171
R789 drain_right.n97 drain_right.n96 8.92171
R790 drain_right.n24 drain_right.n18 8.14595
R791 drain_right.n62 drain_right.n0 8.14595
R792 drain_right.n130 drain_right.n68 8.14595
R793 drain_right.n93 drain_right.n87 8.14595
R794 drain_right.n23 drain_right.n20 7.3702
R795 drain_right.n92 drain_right.n89 7.3702
R796 drain_right drain_right.n133 5.90322
R797 drain_right.n24 drain_right.n23 5.81868
R798 drain_right.n64 drain_right.n0 5.81868
R799 drain_right.n132 drain_right.n68 5.81868
R800 drain_right.n93 drain_right.n92 5.81868
R801 drain_right.n27 drain_right.n18 5.04292
R802 drain_right.n62 drain_right.n61 5.04292
R803 drain_right.n130 drain_right.n129 5.04292
R804 drain_right.n96 drain_right.n87 5.04292
R805 drain_right.n28 drain_right.n16 4.26717
R806 drain_right.n58 drain_right.n2 4.26717
R807 drain_right.n126 drain_right.n70 4.26717
R808 drain_right.n97 drain_right.n85 4.26717
R809 drain_right.n32 drain_right.n31 3.49141
R810 drain_right.n57 drain_right.n4 3.49141
R811 drain_right.n125 drain_right.n72 3.49141
R812 drain_right.n101 drain_right.n100 3.49141
R813 drain_right.n22 drain_right.n21 2.84303
R814 drain_right.n91 drain_right.n90 2.84303
R815 drain_right.n35 drain_right.n14 2.71565
R816 drain_right.n54 drain_right.n53 2.71565
R817 drain_right.n122 drain_right.n121 2.71565
R818 drain_right.n104 drain_right.n83 2.71565
R819 drain_right.n36 drain_right.n12 1.93989
R820 drain_right.n50 drain_right.n6 1.93989
R821 drain_right.n118 drain_right.n74 1.93989
R822 drain_right.n105 drain_right.n81 1.93989
R823 drain_right.n65 drain_right.t4 1.6505
R824 drain_right.n65 drain_right.t1 1.6505
R825 drain_right.n67 drain_right.t5 1.6505
R826 drain_right.n67 drain_right.t2 1.6505
R827 drain_right.n41 drain_right.n39 1.16414
R828 drain_right.n49 drain_right.n8 1.16414
R829 drain_right.n117 drain_right.n76 1.16414
R830 drain_right.n109 drain_right.n108 1.16414
R831 drain_right.n40 drain_right.n10 0.388379
R832 drain_right.n46 drain_right.n45 0.388379
R833 drain_right.n114 drain_right.n113 0.388379
R834 drain_right.n80 drain_right.n78 0.388379
R835 drain_right.n22 drain_right.n17 0.155672
R836 drain_right.n29 drain_right.n17 0.155672
R837 drain_right.n30 drain_right.n29 0.155672
R838 drain_right.n30 drain_right.n13 0.155672
R839 drain_right.n37 drain_right.n13 0.155672
R840 drain_right.n38 drain_right.n37 0.155672
R841 drain_right.n38 drain_right.n9 0.155672
R842 drain_right.n47 drain_right.n9 0.155672
R843 drain_right.n48 drain_right.n47 0.155672
R844 drain_right.n48 drain_right.n5 0.155672
R845 drain_right.n55 drain_right.n5 0.155672
R846 drain_right.n56 drain_right.n55 0.155672
R847 drain_right.n56 drain_right.n1 0.155672
R848 drain_right.n63 drain_right.n1 0.155672
R849 drain_right.n131 drain_right.n69 0.155672
R850 drain_right.n124 drain_right.n69 0.155672
R851 drain_right.n124 drain_right.n123 0.155672
R852 drain_right.n123 drain_right.n73 0.155672
R853 drain_right.n116 drain_right.n73 0.155672
R854 drain_right.n116 drain_right.n115 0.155672
R855 drain_right.n115 drain_right.n77 0.155672
R856 drain_right.n107 drain_right.n77 0.155672
R857 drain_right.n107 drain_right.n106 0.155672
R858 drain_right.n106 drain_right.n82 0.155672
R859 drain_right.n99 drain_right.n82 0.155672
R860 drain_right.n99 drain_right.n98 0.155672
R861 drain_right.n98 drain_right.n86 0.155672
R862 drain_right.n91 drain_right.n86 0.155672
C0 source drain_right 15.099599f
C1 plus drain_right 0.26552f
C2 plus source 1.97593f
C3 minus drain_left 0.170597f
C4 drain_left drain_right 0.551872f
C5 drain_left source 15.111899f
C6 plus drain_left 2.5667f
C7 minus drain_right 2.45959f
C8 minus source 1.96122f
C9 plus minus 4.62222f
C10 drain_right a_n1180_n3288# 6.42256f
C11 drain_left a_n1180_n3288# 6.60579f
C12 source a_n1180_n3288# 6.023682f
C13 minus a_n1180_n3288# 4.508079f
C14 plus a_n1180_n3288# 6.13455f
C15 drain_right.n0 a_n1180_n3288# 0.03836f
C16 drain_right.n1 a_n1180_n3288# 0.028959f
C17 drain_right.n2 a_n1180_n3288# 0.015561f
C18 drain_right.n3 a_n1180_n3288# 0.036781f
C19 drain_right.n4 a_n1180_n3288# 0.016477f
C20 drain_right.n5 a_n1180_n3288# 0.028959f
C21 drain_right.n6 a_n1180_n3288# 0.015561f
C22 drain_right.n7 a_n1180_n3288# 0.036781f
C23 drain_right.n8 a_n1180_n3288# 0.016477f
C24 drain_right.n9 a_n1180_n3288# 0.028959f
C25 drain_right.n10 a_n1180_n3288# 0.016019f
C26 drain_right.n11 a_n1180_n3288# 0.036781f
C27 drain_right.n12 a_n1180_n3288# 0.016477f
C28 drain_right.n13 a_n1180_n3288# 0.028959f
C29 drain_right.n14 a_n1180_n3288# 0.015561f
C30 drain_right.n15 a_n1180_n3288# 0.036781f
C31 drain_right.n16 a_n1180_n3288# 0.016477f
C32 drain_right.n17 a_n1180_n3288# 0.028959f
C33 drain_right.n18 a_n1180_n3288# 0.015561f
C34 drain_right.n19 a_n1180_n3288# 0.027586f
C35 drain_right.n20 a_n1180_n3288# 0.026001f
C36 drain_right.t0 a_n1180_n3288# 0.062121f
C37 drain_right.n21 a_n1180_n3288# 0.20879f
C38 drain_right.n22 a_n1180_n3288# 1.46092f
C39 drain_right.n23 a_n1180_n3288# 0.015561f
C40 drain_right.n24 a_n1180_n3288# 0.016477f
C41 drain_right.n25 a_n1180_n3288# 0.036781f
C42 drain_right.n26 a_n1180_n3288# 0.036781f
C43 drain_right.n27 a_n1180_n3288# 0.016477f
C44 drain_right.n28 a_n1180_n3288# 0.015561f
C45 drain_right.n29 a_n1180_n3288# 0.028959f
C46 drain_right.n30 a_n1180_n3288# 0.028959f
C47 drain_right.n31 a_n1180_n3288# 0.015561f
C48 drain_right.n32 a_n1180_n3288# 0.016477f
C49 drain_right.n33 a_n1180_n3288# 0.036781f
C50 drain_right.n34 a_n1180_n3288# 0.036781f
C51 drain_right.n35 a_n1180_n3288# 0.016477f
C52 drain_right.n36 a_n1180_n3288# 0.015561f
C53 drain_right.n37 a_n1180_n3288# 0.028959f
C54 drain_right.n38 a_n1180_n3288# 0.028959f
C55 drain_right.n39 a_n1180_n3288# 0.015561f
C56 drain_right.n40 a_n1180_n3288# 0.015561f
C57 drain_right.n41 a_n1180_n3288# 0.016477f
C58 drain_right.n42 a_n1180_n3288# 0.036781f
C59 drain_right.n43 a_n1180_n3288# 0.036781f
C60 drain_right.n44 a_n1180_n3288# 0.036781f
C61 drain_right.n45 a_n1180_n3288# 0.016019f
C62 drain_right.n46 a_n1180_n3288# 0.015561f
C63 drain_right.n47 a_n1180_n3288# 0.028959f
C64 drain_right.n48 a_n1180_n3288# 0.028959f
C65 drain_right.n49 a_n1180_n3288# 0.015561f
C66 drain_right.n50 a_n1180_n3288# 0.016477f
C67 drain_right.n51 a_n1180_n3288# 0.036781f
C68 drain_right.n52 a_n1180_n3288# 0.036781f
C69 drain_right.n53 a_n1180_n3288# 0.016477f
C70 drain_right.n54 a_n1180_n3288# 0.015561f
C71 drain_right.n55 a_n1180_n3288# 0.028959f
C72 drain_right.n56 a_n1180_n3288# 0.028959f
C73 drain_right.n57 a_n1180_n3288# 0.015561f
C74 drain_right.n58 a_n1180_n3288# 0.016477f
C75 drain_right.n59 a_n1180_n3288# 0.036781f
C76 drain_right.n60 a_n1180_n3288# 0.075478f
C77 drain_right.n61 a_n1180_n3288# 0.016477f
C78 drain_right.n62 a_n1180_n3288# 0.015561f
C79 drain_right.n63 a_n1180_n3288# 0.06219f
C80 drain_right.n64 a_n1180_n3288# 0.062273f
C81 drain_right.t4 a_n1180_n3288# 0.274609f
C82 drain_right.t1 a_n1180_n3288# 0.274609f
C83 drain_right.n65 a_n1180_n3288# 2.44397f
C84 drain_right.n66 a_n1180_n3288# 1.55005f
C85 drain_right.t5 a_n1180_n3288# 0.274609f
C86 drain_right.t2 a_n1180_n3288# 0.274609f
C87 drain_right.n67 a_n1180_n3288# 2.4465f
C88 drain_right.n68 a_n1180_n3288# 0.03836f
C89 drain_right.n69 a_n1180_n3288# 0.028959f
C90 drain_right.n70 a_n1180_n3288# 0.015561f
C91 drain_right.n71 a_n1180_n3288# 0.036781f
C92 drain_right.n72 a_n1180_n3288# 0.016477f
C93 drain_right.n73 a_n1180_n3288# 0.028959f
C94 drain_right.n74 a_n1180_n3288# 0.015561f
C95 drain_right.n75 a_n1180_n3288# 0.036781f
C96 drain_right.n76 a_n1180_n3288# 0.016477f
C97 drain_right.n77 a_n1180_n3288# 0.028959f
C98 drain_right.n78 a_n1180_n3288# 0.016019f
C99 drain_right.n79 a_n1180_n3288# 0.036781f
C100 drain_right.n80 a_n1180_n3288# 0.015561f
C101 drain_right.n81 a_n1180_n3288# 0.016477f
C102 drain_right.n82 a_n1180_n3288# 0.028959f
C103 drain_right.n83 a_n1180_n3288# 0.015561f
C104 drain_right.n84 a_n1180_n3288# 0.036781f
C105 drain_right.n85 a_n1180_n3288# 0.016477f
C106 drain_right.n86 a_n1180_n3288# 0.028959f
C107 drain_right.n87 a_n1180_n3288# 0.015561f
C108 drain_right.n88 a_n1180_n3288# 0.027586f
C109 drain_right.n89 a_n1180_n3288# 0.026001f
C110 drain_right.t3 a_n1180_n3288# 0.062121f
C111 drain_right.n90 a_n1180_n3288# 0.20879f
C112 drain_right.n91 a_n1180_n3288# 1.46092f
C113 drain_right.n92 a_n1180_n3288# 0.015561f
C114 drain_right.n93 a_n1180_n3288# 0.016477f
C115 drain_right.n94 a_n1180_n3288# 0.036781f
C116 drain_right.n95 a_n1180_n3288# 0.036781f
C117 drain_right.n96 a_n1180_n3288# 0.016477f
C118 drain_right.n97 a_n1180_n3288# 0.015561f
C119 drain_right.n98 a_n1180_n3288# 0.028959f
C120 drain_right.n99 a_n1180_n3288# 0.028959f
C121 drain_right.n100 a_n1180_n3288# 0.015561f
C122 drain_right.n101 a_n1180_n3288# 0.016477f
C123 drain_right.n102 a_n1180_n3288# 0.036781f
C124 drain_right.n103 a_n1180_n3288# 0.036781f
C125 drain_right.n104 a_n1180_n3288# 0.016477f
C126 drain_right.n105 a_n1180_n3288# 0.015561f
C127 drain_right.n106 a_n1180_n3288# 0.028959f
C128 drain_right.n107 a_n1180_n3288# 0.028959f
C129 drain_right.n108 a_n1180_n3288# 0.015561f
C130 drain_right.n109 a_n1180_n3288# 0.016477f
C131 drain_right.n110 a_n1180_n3288# 0.036781f
C132 drain_right.n111 a_n1180_n3288# 0.036781f
C133 drain_right.n112 a_n1180_n3288# 0.036781f
C134 drain_right.n113 a_n1180_n3288# 0.016019f
C135 drain_right.n114 a_n1180_n3288# 0.015561f
C136 drain_right.n115 a_n1180_n3288# 0.028959f
C137 drain_right.n116 a_n1180_n3288# 0.028959f
C138 drain_right.n117 a_n1180_n3288# 0.015561f
C139 drain_right.n118 a_n1180_n3288# 0.016477f
C140 drain_right.n119 a_n1180_n3288# 0.036781f
C141 drain_right.n120 a_n1180_n3288# 0.036781f
C142 drain_right.n121 a_n1180_n3288# 0.016477f
C143 drain_right.n122 a_n1180_n3288# 0.015561f
C144 drain_right.n123 a_n1180_n3288# 0.028959f
C145 drain_right.n124 a_n1180_n3288# 0.028959f
C146 drain_right.n125 a_n1180_n3288# 0.015561f
C147 drain_right.n126 a_n1180_n3288# 0.016477f
C148 drain_right.n127 a_n1180_n3288# 0.036781f
C149 drain_right.n128 a_n1180_n3288# 0.075478f
C150 drain_right.n129 a_n1180_n3288# 0.016477f
C151 drain_right.n130 a_n1180_n3288# 0.015561f
C152 drain_right.n131 a_n1180_n3288# 0.06219f
C153 drain_right.n132 a_n1180_n3288# 0.061693f
C154 drain_right.n133 a_n1180_n3288# 0.683302f
C155 minus.t3 a_n1180_n3288# 0.400599f
C156 minus.n0 a_n1180_n3288# 0.173255f
C157 minus.t2 a_n1180_n3288# 0.400599f
C158 minus.t0 a_n1180_n3288# 0.394756f
C159 minus.n1 a_n1180_n3288# 0.15899f
C160 minus.n2 a_n1180_n3288# 0.173187f
C161 minus.n3 a_n1180_n3288# 1.51825f
C162 minus.t5 a_n1180_n3288# 0.400599f
C163 minus.n4 a_n1180_n3288# 0.173255f
C164 minus.t1 a_n1180_n3288# 0.394756f
C165 minus.n5 a_n1180_n3288# 0.15899f
C166 minus.t4 a_n1180_n3288# 0.400599f
C167 minus.n6 a_n1180_n3288# 0.173187f
C168 minus.n7 a_n1180_n3288# 0.361091f
C169 minus.n8 a_n1180_n3288# 1.78731f
C170 source.n0 a_n1180_n3288# 0.034735f
C171 source.n1 a_n1180_n3288# 0.026222f
C172 source.n2 a_n1180_n3288# 0.014091f
C173 source.n3 a_n1180_n3288# 0.033305f
C174 source.n4 a_n1180_n3288# 0.01492f
C175 source.n5 a_n1180_n3288# 0.026222f
C176 source.n6 a_n1180_n3288# 0.014091f
C177 source.n7 a_n1180_n3288# 0.033305f
C178 source.n8 a_n1180_n3288# 0.01492f
C179 source.n9 a_n1180_n3288# 0.026222f
C180 source.n10 a_n1180_n3288# 0.014505f
C181 source.n11 a_n1180_n3288# 0.033305f
C182 source.n12 a_n1180_n3288# 0.014091f
C183 source.n13 a_n1180_n3288# 0.01492f
C184 source.n14 a_n1180_n3288# 0.026222f
C185 source.n15 a_n1180_n3288# 0.014091f
C186 source.n16 a_n1180_n3288# 0.033305f
C187 source.n17 a_n1180_n3288# 0.01492f
C188 source.n18 a_n1180_n3288# 0.026222f
C189 source.n19 a_n1180_n3288# 0.014091f
C190 source.n20 a_n1180_n3288# 0.024979f
C191 source.n21 a_n1180_n3288# 0.023544f
C192 source.t8 a_n1180_n3288# 0.056251f
C193 source.n22 a_n1180_n3288# 0.18906f
C194 source.n23 a_n1180_n3288# 1.32287f
C195 source.n24 a_n1180_n3288# 0.014091f
C196 source.n25 a_n1180_n3288# 0.01492f
C197 source.n26 a_n1180_n3288# 0.033305f
C198 source.n27 a_n1180_n3288# 0.033305f
C199 source.n28 a_n1180_n3288# 0.01492f
C200 source.n29 a_n1180_n3288# 0.014091f
C201 source.n30 a_n1180_n3288# 0.026222f
C202 source.n31 a_n1180_n3288# 0.026222f
C203 source.n32 a_n1180_n3288# 0.014091f
C204 source.n33 a_n1180_n3288# 0.01492f
C205 source.n34 a_n1180_n3288# 0.033305f
C206 source.n35 a_n1180_n3288# 0.033305f
C207 source.n36 a_n1180_n3288# 0.01492f
C208 source.n37 a_n1180_n3288# 0.014091f
C209 source.n38 a_n1180_n3288# 0.026222f
C210 source.n39 a_n1180_n3288# 0.026222f
C211 source.n40 a_n1180_n3288# 0.014091f
C212 source.n41 a_n1180_n3288# 0.01492f
C213 source.n42 a_n1180_n3288# 0.033305f
C214 source.n43 a_n1180_n3288# 0.033305f
C215 source.n44 a_n1180_n3288# 0.033305f
C216 source.n45 a_n1180_n3288# 0.014505f
C217 source.n46 a_n1180_n3288# 0.014091f
C218 source.n47 a_n1180_n3288# 0.026222f
C219 source.n48 a_n1180_n3288# 0.026222f
C220 source.n49 a_n1180_n3288# 0.014091f
C221 source.n50 a_n1180_n3288# 0.01492f
C222 source.n51 a_n1180_n3288# 0.033305f
C223 source.n52 a_n1180_n3288# 0.033305f
C224 source.n53 a_n1180_n3288# 0.01492f
C225 source.n54 a_n1180_n3288# 0.014091f
C226 source.n55 a_n1180_n3288# 0.026222f
C227 source.n56 a_n1180_n3288# 0.026222f
C228 source.n57 a_n1180_n3288# 0.014091f
C229 source.n58 a_n1180_n3288# 0.01492f
C230 source.n59 a_n1180_n3288# 0.033305f
C231 source.n60 a_n1180_n3288# 0.068346f
C232 source.n61 a_n1180_n3288# 0.01492f
C233 source.n62 a_n1180_n3288# 0.014091f
C234 source.n63 a_n1180_n3288# 0.056313f
C235 source.n64 a_n1180_n3288# 0.03772f
C236 source.n65 a_n1180_n3288# 1.04934f
C237 source.t10 a_n1180_n3288# 0.24866f
C238 source.t11 a_n1180_n3288# 0.24866f
C239 source.n66 a_n1180_n3288# 2.12903f
C240 source.n67 a_n1180_n3288# 0.371158f
C241 source.n68 a_n1180_n3288# 0.034735f
C242 source.n69 a_n1180_n3288# 0.026222f
C243 source.n70 a_n1180_n3288# 0.014091f
C244 source.n71 a_n1180_n3288# 0.033305f
C245 source.n72 a_n1180_n3288# 0.01492f
C246 source.n73 a_n1180_n3288# 0.026222f
C247 source.n74 a_n1180_n3288# 0.014091f
C248 source.n75 a_n1180_n3288# 0.033305f
C249 source.n76 a_n1180_n3288# 0.01492f
C250 source.n77 a_n1180_n3288# 0.026222f
C251 source.n78 a_n1180_n3288# 0.014505f
C252 source.n79 a_n1180_n3288# 0.033305f
C253 source.n80 a_n1180_n3288# 0.014091f
C254 source.n81 a_n1180_n3288# 0.01492f
C255 source.n82 a_n1180_n3288# 0.026222f
C256 source.n83 a_n1180_n3288# 0.014091f
C257 source.n84 a_n1180_n3288# 0.033305f
C258 source.n85 a_n1180_n3288# 0.01492f
C259 source.n86 a_n1180_n3288# 0.026222f
C260 source.n87 a_n1180_n3288# 0.014091f
C261 source.n88 a_n1180_n3288# 0.024979f
C262 source.n89 a_n1180_n3288# 0.023544f
C263 source.t5 a_n1180_n3288# 0.056251f
C264 source.n90 a_n1180_n3288# 0.18906f
C265 source.n91 a_n1180_n3288# 1.32287f
C266 source.n92 a_n1180_n3288# 0.014091f
C267 source.n93 a_n1180_n3288# 0.01492f
C268 source.n94 a_n1180_n3288# 0.033305f
C269 source.n95 a_n1180_n3288# 0.033305f
C270 source.n96 a_n1180_n3288# 0.01492f
C271 source.n97 a_n1180_n3288# 0.014091f
C272 source.n98 a_n1180_n3288# 0.026222f
C273 source.n99 a_n1180_n3288# 0.026222f
C274 source.n100 a_n1180_n3288# 0.014091f
C275 source.n101 a_n1180_n3288# 0.01492f
C276 source.n102 a_n1180_n3288# 0.033305f
C277 source.n103 a_n1180_n3288# 0.033305f
C278 source.n104 a_n1180_n3288# 0.01492f
C279 source.n105 a_n1180_n3288# 0.014091f
C280 source.n106 a_n1180_n3288# 0.026222f
C281 source.n107 a_n1180_n3288# 0.026222f
C282 source.n108 a_n1180_n3288# 0.014091f
C283 source.n109 a_n1180_n3288# 0.01492f
C284 source.n110 a_n1180_n3288# 0.033305f
C285 source.n111 a_n1180_n3288# 0.033305f
C286 source.n112 a_n1180_n3288# 0.033305f
C287 source.n113 a_n1180_n3288# 0.014505f
C288 source.n114 a_n1180_n3288# 0.014091f
C289 source.n115 a_n1180_n3288# 0.026222f
C290 source.n116 a_n1180_n3288# 0.026222f
C291 source.n117 a_n1180_n3288# 0.014091f
C292 source.n118 a_n1180_n3288# 0.01492f
C293 source.n119 a_n1180_n3288# 0.033305f
C294 source.n120 a_n1180_n3288# 0.033305f
C295 source.n121 a_n1180_n3288# 0.01492f
C296 source.n122 a_n1180_n3288# 0.014091f
C297 source.n123 a_n1180_n3288# 0.026222f
C298 source.n124 a_n1180_n3288# 0.026222f
C299 source.n125 a_n1180_n3288# 0.014091f
C300 source.n126 a_n1180_n3288# 0.01492f
C301 source.n127 a_n1180_n3288# 0.033305f
C302 source.n128 a_n1180_n3288# 0.068346f
C303 source.n129 a_n1180_n3288# 0.01492f
C304 source.n130 a_n1180_n3288# 0.014091f
C305 source.n131 a_n1180_n3288# 0.056313f
C306 source.n132 a_n1180_n3288# 0.03772f
C307 source.n133 a_n1180_n3288# 0.123043f
C308 source.t3 a_n1180_n3288# 0.24866f
C309 source.t1 a_n1180_n3288# 0.24866f
C310 source.n134 a_n1180_n3288# 2.12903f
C311 source.n135 a_n1180_n3288# 1.75072f
C312 source.t9 a_n1180_n3288# 0.24866f
C313 source.t7 a_n1180_n3288# 0.24866f
C314 source.n136 a_n1180_n3288# 2.12902f
C315 source.n137 a_n1180_n3288# 1.75073f
C316 source.n138 a_n1180_n3288# 0.034735f
C317 source.n139 a_n1180_n3288# 0.026222f
C318 source.n140 a_n1180_n3288# 0.014091f
C319 source.n141 a_n1180_n3288# 0.033305f
C320 source.n142 a_n1180_n3288# 0.01492f
C321 source.n143 a_n1180_n3288# 0.026222f
C322 source.n144 a_n1180_n3288# 0.014091f
C323 source.n145 a_n1180_n3288# 0.033305f
C324 source.n146 a_n1180_n3288# 0.01492f
C325 source.n147 a_n1180_n3288# 0.026222f
C326 source.n148 a_n1180_n3288# 0.014505f
C327 source.n149 a_n1180_n3288# 0.033305f
C328 source.n150 a_n1180_n3288# 0.01492f
C329 source.n151 a_n1180_n3288# 0.026222f
C330 source.n152 a_n1180_n3288# 0.014091f
C331 source.n153 a_n1180_n3288# 0.033305f
C332 source.n154 a_n1180_n3288# 0.01492f
C333 source.n155 a_n1180_n3288# 0.026222f
C334 source.n156 a_n1180_n3288# 0.014091f
C335 source.n157 a_n1180_n3288# 0.024979f
C336 source.n158 a_n1180_n3288# 0.023544f
C337 source.t6 a_n1180_n3288# 0.056251f
C338 source.n159 a_n1180_n3288# 0.18906f
C339 source.n160 a_n1180_n3288# 1.32287f
C340 source.n161 a_n1180_n3288# 0.014091f
C341 source.n162 a_n1180_n3288# 0.01492f
C342 source.n163 a_n1180_n3288# 0.033305f
C343 source.n164 a_n1180_n3288# 0.033305f
C344 source.n165 a_n1180_n3288# 0.01492f
C345 source.n166 a_n1180_n3288# 0.014091f
C346 source.n167 a_n1180_n3288# 0.026222f
C347 source.n168 a_n1180_n3288# 0.026222f
C348 source.n169 a_n1180_n3288# 0.014091f
C349 source.n170 a_n1180_n3288# 0.01492f
C350 source.n171 a_n1180_n3288# 0.033305f
C351 source.n172 a_n1180_n3288# 0.033305f
C352 source.n173 a_n1180_n3288# 0.01492f
C353 source.n174 a_n1180_n3288# 0.014091f
C354 source.n175 a_n1180_n3288# 0.026222f
C355 source.n176 a_n1180_n3288# 0.026222f
C356 source.n177 a_n1180_n3288# 0.014091f
C357 source.n178 a_n1180_n3288# 0.014091f
C358 source.n179 a_n1180_n3288# 0.01492f
C359 source.n180 a_n1180_n3288# 0.033305f
C360 source.n181 a_n1180_n3288# 0.033305f
C361 source.n182 a_n1180_n3288# 0.033305f
C362 source.n183 a_n1180_n3288# 0.014505f
C363 source.n184 a_n1180_n3288# 0.014091f
C364 source.n185 a_n1180_n3288# 0.026222f
C365 source.n186 a_n1180_n3288# 0.026222f
C366 source.n187 a_n1180_n3288# 0.014091f
C367 source.n188 a_n1180_n3288# 0.01492f
C368 source.n189 a_n1180_n3288# 0.033305f
C369 source.n190 a_n1180_n3288# 0.033305f
C370 source.n191 a_n1180_n3288# 0.01492f
C371 source.n192 a_n1180_n3288# 0.014091f
C372 source.n193 a_n1180_n3288# 0.026222f
C373 source.n194 a_n1180_n3288# 0.026222f
C374 source.n195 a_n1180_n3288# 0.014091f
C375 source.n196 a_n1180_n3288# 0.01492f
C376 source.n197 a_n1180_n3288# 0.033305f
C377 source.n198 a_n1180_n3288# 0.068346f
C378 source.n199 a_n1180_n3288# 0.01492f
C379 source.n200 a_n1180_n3288# 0.014091f
C380 source.n201 a_n1180_n3288# 0.056313f
C381 source.n202 a_n1180_n3288# 0.03772f
C382 source.n203 a_n1180_n3288# 0.123043f
C383 source.t0 a_n1180_n3288# 0.24866f
C384 source.t4 a_n1180_n3288# 0.24866f
C385 source.n204 a_n1180_n3288# 2.12902f
C386 source.n205 a_n1180_n3288# 0.371171f
C387 source.n206 a_n1180_n3288# 0.034735f
C388 source.n207 a_n1180_n3288# 0.026222f
C389 source.n208 a_n1180_n3288# 0.014091f
C390 source.n209 a_n1180_n3288# 0.033305f
C391 source.n210 a_n1180_n3288# 0.01492f
C392 source.n211 a_n1180_n3288# 0.026222f
C393 source.n212 a_n1180_n3288# 0.014091f
C394 source.n213 a_n1180_n3288# 0.033305f
C395 source.n214 a_n1180_n3288# 0.01492f
C396 source.n215 a_n1180_n3288# 0.026222f
C397 source.n216 a_n1180_n3288# 0.014505f
C398 source.n217 a_n1180_n3288# 0.033305f
C399 source.n218 a_n1180_n3288# 0.01492f
C400 source.n219 a_n1180_n3288# 0.026222f
C401 source.n220 a_n1180_n3288# 0.014091f
C402 source.n221 a_n1180_n3288# 0.033305f
C403 source.n222 a_n1180_n3288# 0.01492f
C404 source.n223 a_n1180_n3288# 0.026222f
C405 source.n224 a_n1180_n3288# 0.014091f
C406 source.n225 a_n1180_n3288# 0.024979f
C407 source.n226 a_n1180_n3288# 0.023544f
C408 source.t2 a_n1180_n3288# 0.056251f
C409 source.n227 a_n1180_n3288# 0.18906f
C410 source.n228 a_n1180_n3288# 1.32287f
C411 source.n229 a_n1180_n3288# 0.014091f
C412 source.n230 a_n1180_n3288# 0.01492f
C413 source.n231 a_n1180_n3288# 0.033305f
C414 source.n232 a_n1180_n3288# 0.033305f
C415 source.n233 a_n1180_n3288# 0.01492f
C416 source.n234 a_n1180_n3288# 0.014091f
C417 source.n235 a_n1180_n3288# 0.026222f
C418 source.n236 a_n1180_n3288# 0.026222f
C419 source.n237 a_n1180_n3288# 0.014091f
C420 source.n238 a_n1180_n3288# 0.01492f
C421 source.n239 a_n1180_n3288# 0.033305f
C422 source.n240 a_n1180_n3288# 0.033305f
C423 source.n241 a_n1180_n3288# 0.01492f
C424 source.n242 a_n1180_n3288# 0.014091f
C425 source.n243 a_n1180_n3288# 0.026222f
C426 source.n244 a_n1180_n3288# 0.026222f
C427 source.n245 a_n1180_n3288# 0.014091f
C428 source.n246 a_n1180_n3288# 0.014091f
C429 source.n247 a_n1180_n3288# 0.01492f
C430 source.n248 a_n1180_n3288# 0.033305f
C431 source.n249 a_n1180_n3288# 0.033305f
C432 source.n250 a_n1180_n3288# 0.033305f
C433 source.n251 a_n1180_n3288# 0.014505f
C434 source.n252 a_n1180_n3288# 0.014091f
C435 source.n253 a_n1180_n3288# 0.026222f
C436 source.n254 a_n1180_n3288# 0.026222f
C437 source.n255 a_n1180_n3288# 0.014091f
C438 source.n256 a_n1180_n3288# 0.01492f
C439 source.n257 a_n1180_n3288# 0.033305f
C440 source.n258 a_n1180_n3288# 0.033305f
C441 source.n259 a_n1180_n3288# 0.01492f
C442 source.n260 a_n1180_n3288# 0.014091f
C443 source.n261 a_n1180_n3288# 0.026222f
C444 source.n262 a_n1180_n3288# 0.026222f
C445 source.n263 a_n1180_n3288# 0.014091f
C446 source.n264 a_n1180_n3288# 0.01492f
C447 source.n265 a_n1180_n3288# 0.033305f
C448 source.n266 a_n1180_n3288# 0.068346f
C449 source.n267 a_n1180_n3288# 0.01492f
C450 source.n268 a_n1180_n3288# 0.014091f
C451 source.n269 a_n1180_n3288# 0.056313f
C452 source.n270 a_n1180_n3288# 0.03772f
C453 source.n271 a_n1180_n3288# 0.247029f
C454 source.n272 a_n1180_n3288# 1.643f
C455 drain_left.n0 a_n1180_n3288# 0.038331f
C456 drain_left.n1 a_n1180_n3288# 0.028937f
C457 drain_left.n2 a_n1180_n3288# 0.015549f
C458 drain_left.n3 a_n1180_n3288# 0.036753f
C459 drain_left.n4 a_n1180_n3288# 0.016464f
C460 drain_left.n5 a_n1180_n3288# 0.028937f
C461 drain_left.n6 a_n1180_n3288# 0.015549f
C462 drain_left.n7 a_n1180_n3288# 0.036753f
C463 drain_left.n8 a_n1180_n3288# 0.016464f
C464 drain_left.n9 a_n1180_n3288# 0.028937f
C465 drain_left.n10 a_n1180_n3288# 0.016007f
C466 drain_left.n11 a_n1180_n3288# 0.036753f
C467 drain_left.n12 a_n1180_n3288# 0.016464f
C468 drain_left.n13 a_n1180_n3288# 0.028937f
C469 drain_left.n14 a_n1180_n3288# 0.015549f
C470 drain_left.n15 a_n1180_n3288# 0.036753f
C471 drain_left.n16 a_n1180_n3288# 0.016464f
C472 drain_left.n17 a_n1180_n3288# 0.028937f
C473 drain_left.n18 a_n1180_n3288# 0.015549f
C474 drain_left.n19 a_n1180_n3288# 0.027565f
C475 drain_left.n20 a_n1180_n3288# 0.025982f
C476 drain_left.t3 a_n1180_n3288# 0.062074f
C477 drain_left.n21 a_n1180_n3288# 0.208633f
C478 drain_left.n22 a_n1180_n3288# 1.45983f
C479 drain_left.n23 a_n1180_n3288# 0.015549f
C480 drain_left.n24 a_n1180_n3288# 0.016464f
C481 drain_left.n25 a_n1180_n3288# 0.036753f
C482 drain_left.n26 a_n1180_n3288# 0.036753f
C483 drain_left.n27 a_n1180_n3288# 0.016464f
C484 drain_left.n28 a_n1180_n3288# 0.015549f
C485 drain_left.n29 a_n1180_n3288# 0.028937f
C486 drain_left.n30 a_n1180_n3288# 0.028937f
C487 drain_left.n31 a_n1180_n3288# 0.015549f
C488 drain_left.n32 a_n1180_n3288# 0.016464f
C489 drain_left.n33 a_n1180_n3288# 0.036753f
C490 drain_left.n34 a_n1180_n3288# 0.036753f
C491 drain_left.n35 a_n1180_n3288# 0.016464f
C492 drain_left.n36 a_n1180_n3288# 0.015549f
C493 drain_left.n37 a_n1180_n3288# 0.028937f
C494 drain_left.n38 a_n1180_n3288# 0.028937f
C495 drain_left.n39 a_n1180_n3288# 0.015549f
C496 drain_left.n40 a_n1180_n3288# 0.015549f
C497 drain_left.n41 a_n1180_n3288# 0.016464f
C498 drain_left.n42 a_n1180_n3288# 0.036753f
C499 drain_left.n43 a_n1180_n3288# 0.036753f
C500 drain_left.n44 a_n1180_n3288# 0.036753f
C501 drain_left.n45 a_n1180_n3288# 0.016007f
C502 drain_left.n46 a_n1180_n3288# 0.015549f
C503 drain_left.n47 a_n1180_n3288# 0.028937f
C504 drain_left.n48 a_n1180_n3288# 0.028937f
C505 drain_left.n49 a_n1180_n3288# 0.015549f
C506 drain_left.n50 a_n1180_n3288# 0.016464f
C507 drain_left.n51 a_n1180_n3288# 0.036753f
C508 drain_left.n52 a_n1180_n3288# 0.036753f
C509 drain_left.n53 a_n1180_n3288# 0.016464f
C510 drain_left.n54 a_n1180_n3288# 0.015549f
C511 drain_left.n55 a_n1180_n3288# 0.028937f
C512 drain_left.n56 a_n1180_n3288# 0.028937f
C513 drain_left.n57 a_n1180_n3288# 0.015549f
C514 drain_left.n58 a_n1180_n3288# 0.016464f
C515 drain_left.n59 a_n1180_n3288# 0.036753f
C516 drain_left.n60 a_n1180_n3288# 0.075422f
C517 drain_left.n61 a_n1180_n3288# 0.016464f
C518 drain_left.n62 a_n1180_n3288# 0.015549f
C519 drain_left.n63 a_n1180_n3288# 0.062143f
C520 drain_left.n64 a_n1180_n3288# 0.062226f
C521 drain_left.t0 a_n1180_n3288# 0.274404f
C522 drain_left.t5 a_n1180_n3288# 0.274404f
C523 drain_left.n65 a_n1180_n3288# 2.44214f
C524 drain_left.n66 a_n1180_n3288# 1.60967f
C525 drain_left.n67 a_n1180_n3288# 0.038331f
C526 drain_left.n68 a_n1180_n3288# 0.028937f
C527 drain_left.n69 a_n1180_n3288# 0.015549f
C528 drain_left.n70 a_n1180_n3288# 0.036753f
C529 drain_left.n71 a_n1180_n3288# 0.016464f
C530 drain_left.n72 a_n1180_n3288# 0.028937f
C531 drain_left.n73 a_n1180_n3288# 0.015549f
C532 drain_left.n74 a_n1180_n3288# 0.036753f
C533 drain_left.n75 a_n1180_n3288# 0.016464f
C534 drain_left.n76 a_n1180_n3288# 0.028937f
C535 drain_left.n77 a_n1180_n3288# 0.016007f
C536 drain_left.n78 a_n1180_n3288# 0.036753f
C537 drain_left.n79 a_n1180_n3288# 0.015549f
C538 drain_left.n80 a_n1180_n3288# 0.016464f
C539 drain_left.n81 a_n1180_n3288# 0.028937f
C540 drain_left.n82 a_n1180_n3288# 0.015549f
C541 drain_left.n83 a_n1180_n3288# 0.036753f
C542 drain_left.n84 a_n1180_n3288# 0.016464f
C543 drain_left.n85 a_n1180_n3288# 0.028937f
C544 drain_left.n86 a_n1180_n3288# 0.015549f
C545 drain_left.n87 a_n1180_n3288# 0.027565f
C546 drain_left.n88 a_n1180_n3288# 0.025982f
C547 drain_left.t1 a_n1180_n3288# 0.062074f
C548 drain_left.n89 a_n1180_n3288# 0.208633f
C549 drain_left.n90 a_n1180_n3288# 1.45983f
C550 drain_left.n91 a_n1180_n3288# 0.015549f
C551 drain_left.n92 a_n1180_n3288# 0.016464f
C552 drain_left.n93 a_n1180_n3288# 0.036753f
C553 drain_left.n94 a_n1180_n3288# 0.036753f
C554 drain_left.n95 a_n1180_n3288# 0.016464f
C555 drain_left.n96 a_n1180_n3288# 0.015549f
C556 drain_left.n97 a_n1180_n3288# 0.028937f
C557 drain_left.n98 a_n1180_n3288# 0.028937f
C558 drain_left.n99 a_n1180_n3288# 0.015549f
C559 drain_left.n100 a_n1180_n3288# 0.016464f
C560 drain_left.n101 a_n1180_n3288# 0.036753f
C561 drain_left.n102 a_n1180_n3288# 0.036753f
C562 drain_left.n103 a_n1180_n3288# 0.016464f
C563 drain_left.n104 a_n1180_n3288# 0.015549f
C564 drain_left.n105 a_n1180_n3288# 0.028937f
C565 drain_left.n106 a_n1180_n3288# 0.028937f
C566 drain_left.n107 a_n1180_n3288# 0.015549f
C567 drain_left.n108 a_n1180_n3288# 0.016464f
C568 drain_left.n109 a_n1180_n3288# 0.036753f
C569 drain_left.n110 a_n1180_n3288# 0.036753f
C570 drain_left.n111 a_n1180_n3288# 0.036753f
C571 drain_left.n112 a_n1180_n3288# 0.016007f
C572 drain_left.n113 a_n1180_n3288# 0.015549f
C573 drain_left.n114 a_n1180_n3288# 0.028937f
C574 drain_left.n115 a_n1180_n3288# 0.028937f
C575 drain_left.n116 a_n1180_n3288# 0.015549f
C576 drain_left.n117 a_n1180_n3288# 0.016464f
C577 drain_left.n118 a_n1180_n3288# 0.036753f
C578 drain_left.n119 a_n1180_n3288# 0.036753f
C579 drain_left.n120 a_n1180_n3288# 0.016464f
C580 drain_left.n121 a_n1180_n3288# 0.015549f
C581 drain_left.n122 a_n1180_n3288# 0.028937f
C582 drain_left.n123 a_n1180_n3288# 0.028937f
C583 drain_left.n124 a_n1180_n3288# 0.015549f
C584 drain_left.n125 a_n1180_n3288# 0.016464f
C585 drain_left.n126 a_n1180_n3288# 0.036753f
C586 drain_left.n127 a_n1180_n3288# 0.075422f
C587 drain_left.n128 a_n1180_n3288# 0.016464f
C588 drain_left.n129 a_n1180_n3288# 0.015549f
C589 drain_left.n130 a_n1180_n3288# 0.062143f
C590 drain_left.n131 a_n1180_n3288# 0.062706f
C591 drain_left.t2 a_n1180_n3288# 0.274404f
C592 drain_left.t4 a_n1180_n3288# 0.274404f
C593 drain_left.n132 a_n1180_n3288# 2.44177f
C594 drain_left.n133 a_n1180_n3288# 0.673523f
C595 plus.t1 a_n1180_n3288# 0.411702f
C596 plus.n0 a_n1180_n3288# 0.178057f
C597 plus.t0 a_n1180_n3288# 0.405696f
C598 plus.n1 a_n1180_n3288# 0.163396f
C599 plus.t3 a_n1180_n3288# 0.411702f
C600 plus.n2 a_n1180_n3288# 0.177987f
C601 plus.n3 a_n1180_n3288# 0.59364f
C602 plus.t5 a_n1180_n3288# 0.411702f
C603 plus.n4 a_n1180_n3288# 0.178057f
C604 plus.t2 a_n1180_n3288# 0.411702f
C605 plus.t4 a_n1180_n3288# 0.405696f
C606 plus.n5 a_n1180_n3288# 0.163396f
C607 plus.n6 a_n1180_n3288# 0.177987f
C608 plus.n7 a_n1180_n3288# 1.32287f
.ends

