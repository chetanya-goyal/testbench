* NGSPICE file created from diffpair59.ext - technology: sky130A

.subckt diffpair59 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t40 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X1 a_n3134_n1088# a_n3134_n1088# a_n3134_n1088# a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.6
X2 drain_left.t22 plus.t1 source.t41 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X3 source.t42 plus.t2 drain_left.t21 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X4 drain_left.t20 plus.t3 source.t39 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X5 source.t18 minus.t0 drain_right.t23 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X6 source.t31 plus.t4 drain_left.t19 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X7 source.t25 plus.t5 drain_left.t18 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X8 drain_right.t22 minus.t1 source.t22 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X9 a_n3134_n1088# a_n3134_n1088# a_n3134_n1088# a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X10 drain_left.t17 plus.t6 source.t45 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X11 source.t5 minus.t2 drain_right.t21 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X12 drain_right.t20 minus.t3 source.t21 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X13 drain_right.t19 minus.t4 source.t7 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X14 drain_right.t18 minus.t5 source.t13 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X15 source.t17 minus.t6 drain_right.t17 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X16 source.t4 minus.t7 drain_right.t16 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X17 source.t29 plus.t7 drain_left.t16 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X18 source.t47 plus.t8 drain_left.t15 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X19 drain_right.t15 minus.t8 source.t1 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X20 source.t3 minus.t9 drain_right.t14 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X21 drain_right.t13 minus.t10 source.t6 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X22 source.t46 plus.t9 drain_left.t14 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X23 drain_left.t13 plus.t10 source.t34 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X24 source.t35 plus.t11 drain_left.t12 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X25 source.t12 minus.t11 drain_right.t12 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X26 source.t16 minus.t12 drain_right.t11 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X27 a_n3134_n1088# a_n3134_n1088# a_n3134_n1088# a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X28 drain_right.t10 minus.t13 source.t0 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X29 drain_left.t11 plus.t12 source.t43 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X30 drain_left.t10 plus.t13 source.t32 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X31 source.t20 minus.t14 drain_right.t9 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X32 drain_left.t9 plus.t14 source.t24 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X33 source.t33 plus.t15 drain_left.t8 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X34 drain_right.t8 minus.t15 source.t2 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X35 a_n3134_n1088# a_n3134_n1088# a_n3134_n1088# a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.6
X36 drain_right.t7 minus.t16 source.t11 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X37 drain_left.t7 plus.t16 source.t27 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X38 drain_left.t6 plus.t17 source.t30 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.6
X39 drain_left.t5 plus.t18 source.t44 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X40 source.t37 plus.t19 drain_left.t4 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X41 source.t38 plus.t20 drain_left.t3 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X42 source.t15 minus.t17 drain_right.t6 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X43 drain_right.t5 minus.t18 source.t9 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X44 source.t28 plus.t21 drain_left.t2 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X45 source.t10 minus.t19 drain_right.t4 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X46 source.t14 minus.t20 drain_right.t3 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X47 drain_right.t2 minus.t21 source.t8 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X48 source.t26 plus.t22 drain_left.t1 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X49 drain_right.t1 minus.t22 source.t23 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
X50 source.t19 minus.t23 drain_right.t0 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.6
X51 drain_left.t0 plus.t23 source.t36 a_n3134_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.6
R0 plus.n13 plus.n8 161.3
R1 plus.n15 plus.n14 161.3
R2 plus.n16 plus.n7 161.3
R3 plus.n18 plus.n17 161.3
R4 plus.n19 plus.n6 161.3
R5 plus.n21 plus.n20 161.3
R6 plus.n22 plus.n5 161.3
R7 plus.n24 plus.n23 161.3
R8 plus.n25 plus.n4 161.3
R9 plus.n27 plus.n26 161.3
R10 plus.n28 plus.n3 161.3
R11 plus.n30 plus.n1 161.3
R12 plus.n31 plus.n0 161.3
R13 plus.n33 plus.n32 161.3
R14 plus.n47 plus.n42 161.3
R15 plus.n49 plus.n48 161.3
R16 plus.n50 plus.n41 161.3
R17 plus.n52 plus.n51 161.3
R18 plus.n53 plus.n40 161.3
R19 plus.n55 plus.n54 161.3
R20 plus.n56 plus.n39 161.3
R21 plus.n58 plus.n57 161.3
R22 plus.n59 plus.n38 161.3
R23 plus.n61 plus.n60 161.3
R24 plus.n62 plus.n37 161.3
R25 plus.n64 plus.n35 161.3
R26 plus.n65 plus.n34 161.3
R27 plus.n67 plus.n66 161.3
R28 plus.n9 plus.t19 131.998
R29 plus.n43 plus.t12 131.998
R30 plus.n32 plus.t17 105.638
R31 plus.n30 plus.t20 105.638
R32 plus.n29 plus.t0 105.638
R33 plus.n28 plus.t2 105.638
R34 plus.n4 plus.t3 105.638
R35 plus.n22 plus.t5 105.638
R36 plus.n6 plus.t6 105.638
R37 plus.n16 plus.t11 105.638
R38 plus.n8 plus.t13 105.638
R39 plus.n11 plus.t15 105.638
R40 plus.n10 plus.t18 105.638
R41 plus.n66 plus.t8 105.638
R42 plus.n64 plus.t10 105.638
R43 plus.n63 plus.t7 105.638
R44 plus.n62 plus.t16 105.638
R45 plus.n38 plus.t22 105.638
R46 plus.n56 plus.t1 105.638
R47 plus.n40 plus.t9 105.638
R48 plus.n50 plus.t14 105.638
R49 plus.n42 plus.t21 105.638
R50 plus.n45 plus.t23 105.638
R51 plus.n44 plus.t4 105.638
R52 plus.n12 plus.n11 80.6037
R53 plus.n29 plus.n2 80.6037
R54 plus.n46 plus.n45 80.6037
R55 plus.n63 plus.n36 80.6037
R56 plus.n30 plus.n29 48.2005
R57 plus.n29 plus.n28 48.2005
R58 plus.n11 plus.n8 48.2005
R59 plus.n11 plus.n10 48.2005
R60 plus.n64 plus.n63 48.2005
R61 plus.n63 plus.n62 48.2005
R62 plus.n45 plus.n42 48.2005
R63 plus.n45 plus.n44 48.2005
R64 plus.n32 plus.n31 46.0096
R65 plus.n66 plus.n65 46.0096
R66 plus.n12 plus.n9 45.1822
R67 plus.n46 plus.n43 45.1822
R68 plus.n27 plus.n4 44.549
R69 plus.n16 plus.n15 44.549
R70 plus.n61 plus.n38 44.549
R71 plus.n50 plus.n49 44.549
R72 plus.n23 plus.n22 34.3247
R73 plus.n17 plus.n6 34.3247
R74 plus.n57 plus.n56 34.3247
R75 plus.n51 plus.n40 34.3247
R76 plus plus.n67 30.8096
R77 plus.n21 plus.n6 24.1005
R78 plus.n22 plus.n21 24.1005
R79 plus.n56 plus.n55 24.1005
R80 plus.n55 plus.n40 24.1005
R81 plus.n10 plus.n9 14.1472
R82 plus.n44 plus.n43 14.1472
R83 plus.n23 plus.n4 13.8763
R84 plus.n17 plus.n16 13.8763
R85 plus.n57 plus.n38 13.8763
R86 plus.n51 plus.n50 13.8763
R87 plus plus.n33 8.08005
R88 plus.n28 plus.n27 3.65202
R89 plus.n15 plus.n8 3.65202
R90 plus.n62 plus.n61 3.65202
R91 plus.n49 plus.n42 3.65202
R92 plus.n31 plus.n30 2.19141
R93 plus.n65 plus.n64 2.19141
R94 plus.n13 plus.n12 0.285035
R95 plus.n3 plus.n2 0.285035
R96 plus.n2 plus.n1 0.285035
R97 plus.n36 plus.n35 0.285035
R98 plus.n37 plus.n36 0.285035
R99 plus.n47 plus.n46 0.285035
R100 plus.n14 plus.n13 0.189894
R101 plus.n14 plus.n7 0.189894
R102 plus.n18 plus.n7 0.189894
R103 plus.n19 plus.n18 0.189894
R104 plus.n20 plus.n19 0.189894
R105 plus.n20 plus.n5 0.189894
R106 plus.n24 plus.n5 0.189894
R107 plus.n25 plus.n24 0.189894
R108 plus.n26 plus.n25 0.189894
R109 plus.n26 plus.n3 0.189894
R110 plus.n1 plus.n0 0.189894
R111 plus.n33 plus.n0 0.189894
R112 plus.n67 plus.n34 0.189894
R113 plus.n35 plus.n34 0.189894
R114 plus.n60 plus.n37 0.189894
R115 plus.n60 plus.n59 0.189894
R116 plus.n59 plus.n58 0.189894
R117 plus.n58 plus.n39 0.189894
R118 plus.n54 plus.n39 0.189894
R119 plus.n54 plus.n53 0.189894
R120 plus.n53 plus.n52 0.189894
R121 plus.n52 plus.n41 0.189894
R122 plus.n48 plus.n41 0.189894
R123 plus.n48 plus.n47 0.189894
R124 source.n0 source.t30 243.255
R125 source.n11 source.t37 243.255
R126 source.n12 source.t2 243.255
R127 source.n23 source.t16 243.255
R128 source.n47 source.t1 243.254
R129 source.n36 source.t19 243.254
R130 source.n35 source.t43 243.254
R131 source.n24 source.t47 243.254
R132 source.n2 source.n1 223.454
R133 source.n4 source.n3 223.454
R134 source.n6 source.n5 223.454
R135 source.n8 source.n7 223.454
R136 source.n10 source.n9 223.454
R137 source.n14 source.n13 223.454
R138 source.n16 source.n15 223.454
R139 source.n18 source.n17 223.454
R140 source.n20 source.n19 223.454
R141 source.n22 source.n21 223.454
R142 source.n46 source.n45 223.453
R143 source.n44 source.n43 223.453
R144 source.n42 source.n41 223.453
R145 source.n40 source.n39 223.453
R146 source.n38 source.n37 223.453
R147 source.n34 source.n33 223.453
R148 source.n32 source.n31 223.453
R149 source.n30 source.n29 223.453
R150 source.n28 source.n27 223.453
R151 source.n26 source.n25 223.453
R152 source.n45 source.t11 19.8005
R153 source.n45 source.t10 19.8005
R154 source.n43 source.t13 19.8005
R155 source.n43 source.t14 19.8005
R156 source.n41 source.t8 19.8005
R157 source.n41 source.t3 19.8005
R158 source.n39 source.t23 19.8005
R159 source.n39 source.t15 19.8005
R160 source.n37 source.t6 19.8005
R161 source.n37 source.t4 19.8005
R162 source.n33 source.t36 19.8005
R163 source.n33 source.t31 19.8005
R164 source.n31 source.t24 19.8005
R165 source.n31 source.t28 19.8005
R166 source.n29 source.t41 19.8005
R167 source.n29 source.t46 19.8005
R168 source.n27 source.t27 19.8005
R169 source.n27 source.t26 19.8005
R170 source.n25 source.t34 19.8005
R171 source.n25 source.t29 19.8005
R172 source.n1 source.t40 19.8005
R173 source.n1 source.t38 19.8005
R174 source.n3 source.t39 19.8005
R175 source.n3 source.t42 19.8005
R176 source.n5 source.t45 19.8005
R177 source.n5 source.t25 19.8005
R178 source.n7 source.t32 19.8005
R179 source.n7 source.t35 19.8005
R180 source.n9 source.t44 19.8005
R181 source.n9 source.t33 19.8005
R182 source.n13 source.t0 19.8005
R183 source.n13 source.t20 19.8005
R184 source.n15 source.t21 19.8005
R185 source.n15 source.t12 19.8005
R186 source.n17 source.t7 19.8005
R187 source.n17 source.t17 19.8005
R188 source.n19 source.t22 19.8005
R189 source.n19 source.t5 19.8005
R190 source.n21 source.t9 19.8005
R191 source.n21 source.t18 19.8005
R192 source.n24 source.n23 13.7561
R193 source.n48 source.n0 8.09232
R194 source.n48 source.n47 5.66429
R195 source.n23 source.n22 0.802224
R196 source.n22 source.n20 0.802224
R197 source.n20 source.n18 0.802224
R198 source.n18 source.n16 0.802224
R199 source.n16 source.n14 0.802224
R200 source.n14 source.n12 0.802224
R201 source.n11 source.n10 0.802224
R202 source.n10 source.n8 0.802224
R203 source.n8 source.n6 0.802224
R204 source.n6 source.n4 0.802224
R205 source.n4 source.n2 0.802224
R206 source.n2 source.n0 0.802224
R207 source.n26 source.n24 0.802224
R208 source.n28 source.n26 0.802224
R209 source.n30 source.n28 0.802224
R210 source.n32 source.n30 0.802224
R211 source.n34 source.n32 0.802224
R212 source.n35 source.n34 0.802224
R213 source.n38 source.n36 0.802224
R214 source.n40 source.n38 0.802224
R215 source.n42 source.n40 0.802224
R216 source.n44 source.n42 0.802224
R217 source.n46 source.n44 0.802224
R218 source.n47 source.n46 0.802224
R219 source.n12 source.n11 0.470328
R220 source.n36 source.n35 0.470328
R221 source source.n48 0.188
R222 drain_left.n13 drain_left.n11 240.935
R223 drain_left.n7 drain_left.n5 240.934
R224 drain_left.n2 drain_left.n0 240.934
R225 drain_left.n21 drain_left.n20 240.132
R226 drain_left.n19 drain_left.n18 240.132
R227 drain_left.n17 drain_left.n16 240.132
R228 drain_left.n15 drain_left.n14 240.132
R229 drain_left.n13 drain_left.n12 240.132
R230 drain_left.n7 drain_left.n6 240.131
R231 drain_left.n9 drain_left.n8 240.131
R232 drain_left.n4 drain_left.n3 240.131
R233 drain_left.n2 drain_left.n1 240.131
R234 drain_left drain_left.n10 26.6501
R235 drain_left.n5 drain_left.t19 19.8005
R236 drain_left.n5 drain_left.t11 19.8005
R237 drain_left.n6 drain_left.t2 19.8005
R238 drain_left.n6 drain_left.t0 19.8005
R239 drain_left.n8 drain_left.t14 19.8005
R240 drain_left.n8 drain_left.t9 19.8005
R241 drain_left.n3 drain_left.t1 19.8005
R242 drain_left.n3 drain_left.t22 19.8005
R243 drain_left.n1 drain_left.t16 19.8005
R244 drain_left.n1 drain_left.t7 19.8005
R245 drain_left.n0 drain_left.t15 19.8005
R246 drain_left.n0 drain_left.t13 19.8005
R247 drain_left.n20 drain_left.t3 19.8005
R248 drain_left.n20 drain_left.t6 19.8005
R249 drain_left.n18 drain_left.t21 19.8005
R250 drain_left.n18 drain_left.t23 19.8005
R251 drain_left.n16 drain_left.t18 19.8005
R252 drain_left.n16 drain_left.t20 19.8005
R253 drain_left.n14 drain_left.t12 19.8005
R254 drain_left.n14 drain_left.t17 19.8005
R255 drain_left.n12 drain_left.t8 19.8005
R256 drain_left.n12 drain_left.t10 19.8005
R257 drain_left.n11 drain_left.t4 19.8005
R258 drain_left.n11 drain_left.t5 19.8005
R259 drain_left drain_left.n21 6.45494
R260 drain_left.n9 drain_left.n7 0.802224
R261 drain_left.n4 drain_left.n2 0.802224
R262 drain_left.n15 drain_left.n13 0.802224
R263 drain_left.n17 drain_left.n15 0.802224
R264 drain_left.n19 drain_left.n17 0.802224
R265 drain_left.n21 drain_left.n19 0.802224
R266 drain_left.n10 drain_left.n9 0.346016
R267 drain_left.n10 drain_left.n4 0.346016
R268 minus.n33 minus.n32 161.3
R269 minus.n31 minus.n0 161.3
R270 minus.n30 minus.n29 161.3
R271 minus.n27 minus.n26 161.3
R272 minus.n25 minus.n2 161.3
R273 minus.n24 minus.n23 161.3
R274 minus.n22 minus.n3 161.3
R275 minus.n21 minus.n20 161.3
R276 minus.n19 minus.n4 161.3
R277 minus.n18 minus.n17 161.3
R278 minus.n16 minus.n5 161.3
R279 minus.n15 minus.n14 161.3
R280 minus.n13 minus.n6 161.3
R281 minus.n12 minus.n11 161.3
R282 minus.n67 minus.n66 161.3
R283 minus.n65 minus.n34 161.3
R284 minus.n64 minus.n63 161.3
R285 minus.n61 minus.n60 161.3
R286 minus.n59 minus.n36 161.3
R287 minus.n58 minus.n57 161.3
R288 minus.n56 minus.n37 161.3
R289 minus.n55 minus.n54 161.3
R290 minus.n53 minus.n38 161.3
R291 minus.n52 minus.n51 161.3
R292 minus.n50 minus.n39 161.3
R293 minus.n49 minus.n48 161.3
R294 minus.n47 minus.n40 161.3
R295 minus.n46 minus.n45 161.3
R296 minus.n9 minus.t15 131.998
R297 minus.n43 minus.t23 131.998
R298 minus.n8 minus.t14 105.638
R299 minus.n7 minus.t13 105.638
R300 minus.n12 minus.t11 105.638
R301 minus.n14 minus.t3 105.638
R302 minus.n18 minus.t6 105.638
R303 minus.n20 minus.t4 105.638
R304 minus.n24 minus.t2 105.638
R305 minus.n26 minus.t1 105.638
R306 minus.n1 minus.t0 105.638
R307 minus.n30 minus.t18 105.638
R308 minus.n32 minus.t12 105.638
R309 minus.n42 minus.t10 105.638
R310 minus.n41 minus.t7 105.638
R311 minus.n46 minus.t22 105.638
R312 minus.n48 minus.t17 105.638
R313 minus.n52 minus.t21 105.638
R314 minus.n54 minus.t9 105.638
R315 minus.n58 minus.t5 105.638
R316 minus.n60 minus.t20 105.638
R317 minus.n35 minus.t16 105.638
R318 minus.n64 minus.t19 105.638
R319 minus.n66 minus.t8 105.638
R320 minus.n28 minus.n1 80.6037
R321 minus.n10 minus.n7 80.6037
R322 minus.n62 minus.n35 80.6037
R323 minus.n44 minus.n41 80.6037
R324 minus.n8 minus.n7 48.2005
R325 minus.n12 minus.n7 48.2005
R326 minus.n26 minus.n1 48.2005
R327 minus.n30 minus.n1 48.2005
R328 minus.n42 minus.n41 48.2005
R329 minus.n46 minus.n41 48.2005
R330 minus.n60 minus.n35 48.2005
R331 minus.n64 minus.n35 48.2005
R332 minus.n32 minus.n31 46.0096
R333 minus.n66 minus.n65 46.0096
R334 minus.n10 minus.n9 45.1822
R335 minus.n44 minus.n43 45.1822
R336 minus.n14 minus.n13 44.549
R337 minus.n25 minus.n24 44.549
R338 minus.n48 minus.n47 44.549
R339 minus.n59 minus.n58 44.549
R340 minus.n18 minus.n5 34.3247
R341 minus.n20 minus.n3 34.3247
R342 minus.n52 minus.n39 34.3247
R343 minus.n54 minus.n37 34.3247
R344 minus.n68 minus.n33 32.7619
R345 minus.n20 minus.n19 24.1005
R346 minus.n19 minus.n18 24.1005
R347 minus.n53 minus.n52 24.1005
R348 minus.n54 minus.n53 24.1005
R349 minus.n9 minus.n8 14.1472
R350 minus.n43 minus.n42 14.1472
R351 minus.n14 minus.n5 13.8763
R352 minus.n24 minus.n3 13.8763
R353 minus.n48 minus.n39 13.8763
R354 minus.n58 minus.n37 13.8763
R355 minus.n68 minus.n67 6.60277
R356 minus.n13 minus.n12 3.65202
R357 minus.n26 minus.n25 3.65202
R358 minus.n47 minus.n46 3.65202
R359 minus.n60 minus.n59 3.65202
R360 minus.n31 minus.n30 2.19141
R361 minus.n65 minus.n64 2.19141
R362 minus.n29 minus.n28 0.285035
R363 minus.n28 minus.n27 0.285035
R364 minus.n11 minus.n10 0.285035
R365 minus.n45 minus.n44 0.285035
R366 minus.n62 minus.n61 0.285035
R367 minus.n63 minus.n62 0.285035
R368 minus.n33 minus.n0 0.189894
R369 minus.n29 minus.n0 0.189894
R370 minus.n27 minus.n2 0.189894
R371 minus.n23 minus.n2 0.189894
R372 minus.n23 minus.n22 0.189894
R373 minus.n22 minus.n21 0.189894
R374 minus.n21 minus.n4 0.189894
R375 minus.n17 minus.n4 0.189894
R376 minus.n17 minus.n16 0.189894
R377 minus.n16 minus.n15 0.189894
R378 minus.n15 minus.n6 0.189894
R379 minus.n11 minus.n6 0.189894
R380 minus.n45 minus.n40 0.189894
R381 minus.n49 minus.n40 0.189894
R382 minus.n50 minus.n49 0.189894
R383 minus.n51 minus.n50 0.189894
R384 minus.n51 minus.n38 0.189894
R385 minus.n55 minus.n38 0.189894
R386 minus.n56 minus.n55 0.189894
R387 minus.n57 minus.n56 0.189894
R388 minus.n57 minus.n36 0.189894
R389 minus.n61 minus.n36 0.189894
R390 minus.n63 minus.n34 0.189894
R391 minus.n67 minus.n34 0.189894
R392 minus minus.n68 0.188
R393 drain_right.n13 drain_right.n11 240.935
R394 drain_right.n7 drain_right.n5 240.934
R395 drain_right.n2 drain_right.n0 240.934
R396 drain_right.n13 drain_right.n12 240.132
R397 drain_right.n15 drain_right.n14 240.132
R398 drain_right.n17 drain_right.n16 240.132
R399 drain_right.n19 drain_right.n18 240.132
R400 drain_right.n21 drain_right.n20 240.132
R401 drain_right.n7 drain_right.n6 240.131
R402 drain_right.n9 drain_right.n8 240.131
R403 drain_right.n4 drain_right.n3 240.131
R404 drain_right.n2 drain_right.n1 240.131
R405 drain_right drain_right.n10 26.0969
R406 drain_right.n5 drain_right.t4 19.8005
R407 drain_right.n5 drain_right.t15 19.8005
R408 drain_right.n6 drain_right.t3 19.8005
R409 drain_right.n6 drain_right.t7 19.8005
R410 drain_right.n8 drain_right.t14 19.8005
R411 drain_right.n8 drain_right.t18 19.8005
R412 drain_right.n3 drain_right.t6 19.8005
R413 drain_right.n3 drain_right.t2 19.8005
R414 drain_right.n1 drain_right.t16 19.8005
R415 drain_right.n1 drain_right.t1 19.8005
R416 drain_right.n0 drain_right.t0 19.8005
R417 drain_right.n0 drain_right.t13 19.8005
R418 drain_right.n11 drain_right.t9 19.8005
R419 drain_right.n11 drain_right.t8 19.8005
R420 drain_right.n12 drain_right.t12 19.8005
R421 drain_right.n12 drain_right.t10 19.8005
R422 drain_right.n14 drain_right.t17 19.8005
R423 drain_right.n14 drain_right.t20 19.8005
R424 drain_right.n16 drain_right.t21 19.8005
R425 drain_right.n16 drain_right.t19 19.8005
R426 drain_right.n18 drain_right.t23 19.8005
R427 drain_right.n18 drain_right.t22 19.8005
R428 drain_right.n20 drain_right.t11 19.8005
R429 drain_right.n20 drain_right.t5 19.8005
R430 drain_right drain_right.n21 6.45494
R431 drain_right.n9 drain_right.n7 0.802224
R432 drain_right.n4 drain_right.n2 0.802224
R433 drain_right.n21 drain_right.n19 0.802224
R434 drain_right.n19 drain_right.n17 0.802224
R435 drain_right.n17 drain_right.n15 0.802224
R436 drain_right.n15 drain_right.n13 0.802224
R437 drain_right.n10 drain_right.n9 0.346016
R438 drain_right.n10 drain_right.n4 0.346016
C0 minus drain_left 0.181851f
C1 source drain_left 6.68584f
C2 minus source 2.69406f
C3 plus drain_right 0.480445f
C4 drain_left drain_right 1.71735f
C5 minus drain_right 1.83148f
C6 source drain_right 6.68787f
C7 plus drain_left 2.14456f
C8 minus plus 5.03424f
C9 plus source 2.70792f
C10 drain_right a_n3134_n1088# 5.12661f
C11 drain_left a_n3134_n1088# 5.963059f
C12 source a_n3134_n1088# 3.004243f
C13 minus a_n3134_n1088# 11.708188f
C14 plus a_n3134_n1088# 13.123679f
C15 drain_right.t0 a_n3134_n1088# 0.017039f
C16 drain_right.t13 a_n3134_n1088# 0.017039f
C17 drain_right.n0 a_n3134_n1088# 0.067111f
C18 drain_right.t16 a_n3134_n1088# 0.017039f
C19 drain_right.t1 a_n3134_n1088# 0.017039f
C20 drain_right.n1 a_n3134_n1088# 0.06621f
C21 drain_right.n2 a_n3134_n1088# 0.532174f
C22 drain_right.t6 a_n3134_n1088# 0.017039f
C23 drain_right.t2 a_n3134_n1088# 0.017039f
C24 drain_right.n3 a_n3134_n1088# 0.06621f
C25 drain_right.n4 a_n3134_n1088# 0.231945f
C26 drain_right.t4 a_n3134_n1088# 0.017039f
C27 drain_right.t15 a_n3134_n1088# 0.017039f
C28 drain_right.n5 a_n3134_n1088# 0.067111f
C29 drain_right.t3 a_n3134_n1088# 0.017039f
C30 drain_right.t7 a_n3134_n1088# 0.017039f
C31 drain_right.n6 a_n3134_n1088# 0.06621f
C32 drain_right.n7 a_n3134_n1088# 0.532174f
C33 drain_right.t14 a_n3134_n1088# 0.017039f
C34 drain_right.t18 a_n3134_n1088# 0.017039f
C35 drain_right.n8 a_n3134_n1088# 0.06621f
C36 drain_right.n9 a_n3134_n1088# 0.231945f
C37 drain_right.n10 a_n3134_n1088# 0.826518f
C38 drain_right.t9 a_n3134_n1088# 0.017039f
C39 drain_right.t8 a_n3134_n1088# 0.017039f
C40 drain_right.n11 a_n3134_n1088# 0.067111f
C41 drain_right.t12 a_n3134_n1088# 0.017039f
C42 drain_right.t10 a_n3134_n1088# 0.017039f
C43 drain_right.n12 a_n3134_n1088# 0.06621f
C44 drain_right.n13 a_n3134_n1088# 0.532174f
C45 drain_right.t17 a_n3134_n1088# 0.017039f
C46 drain_right.t20 a_n3134_n1088# 0.017039f
C47 drain_right.n14 a_n3134_n1088# 0.06621f
C48 drain_right.n15 a_n3134_n1088# 0.262195f
C49 drain_right.t21 a_n3134_n1088# 0.017039f
C50 drain_right.t19 a_n3134_n1088# 0.017039f
C51 drain_right.n16 a_n3134_n1088# 0.06621f
C52 drain_right.n17 a_n3134_n1088# 0.262195f
C53 drain_right.t23 a_n3134_n1088# 0.017039f
C54 drain_right.t22 a_n3134_n1088# 0.017039f
C55 drain_right.n18 a_n3134_n1088# 0.06621f
C56 drain_right.n19 a_n3134_n1088# 0.262195f
C57 drain_right.t11 a_n3134_n1088# 0.017039f
C58 drain_right.t5 a_n3134_n1088# 0.017039f
C59 drain_right.n20 a_n3134_n1088# 0.06621f
C60 drain_right.n21 a_n3134_n1088# 0.450219f
C61 minus.n0 a_n3134_n1088# 0.035312f
C62 minus.t0 a_n3134_n1088# 0.071845f
C63 minus.n1 a_n3134_n1088# 0.081141f
C64 minus.t18 a_n3134_n1088# 0.071845f
C65 minus.n2 a_n3134_n1088# 0.035312f
C66 minus.n3 a_n3134_n1088# 0.008013f
C67 minus.t2 a_n3134_n1088# 0.071845f
C68 minus.n4 a_n3134_n1088# 0.035312f
C69 minus.n5 a_n3134_n1088# 0.008013f
C70 minus.t6 a_n3134_n1088# 0.071845f
C71 minus.n6 a_n3134_n1088# 0.035312f
C72 minus.t13 a_n3134_n1088# 0.071845f
C73 minus.n7 a_n3134_n1088# 0.081141f
C74 minus.t11 a_n3134_n1088# 0.071845f
C75 minus.t15 a_n3134_n1088# 0.086439f
C76 minus.t14 a_n3134_n1088# 0.071845f
C77 minus.n8 a_n3134_n1088# 0.080681f
C78 minus.n9 a_n3134_n1088# 0.060037f
C79 minus.n10 a_n3134_n1088# 0.170892f
C80 minus.n11 a_n3134_n1088# 0.047119f
C81 minus.n12 a_n3134_n1088# 0.073673f
C82 minus.n13 a_n3134_n1088# 0.008013f
C83 minus.t3 a_n3134_n1088# 0.071845f
C84 minus.n14 a_n3134_n1088# 0.074652f
C85 minus.n15 a_n3134_n1088# 0.035312f
C86 minus.n16 a_n3134_n1088# 0.035312f
C87 minus.n17 a_n3134_n1088# 0.035312f
C88 minus.n18 a_n3134_n1088# 0.074652f
C89 minus.n19 a_n3134_n1088# 0.008013f
C90 minus.t4 a_n3134_n1088# 0.071845f
C91 minus.n20 a_n3134_n1088# 0.074652f
C92 minus.n21 a_n3134_n1088# 0.035312f
C93 minus.n22 a_n3134_n1088# 0.035312f
C94 minus.n23 a_n3134_n1088# 0.035312f
C95 minus.n24 a_n3134_n1088# 0.074652f
C96 minus.n25 a_n3134_n1088# 0.008013f
C97 minus.t1 a_n3134_n1088# 0.071845f
C98 minus.n26 a_n3134_n1088# 0.073673f
C99 minus.n27 a_n3134_n1088# 0.047119f
C100 minus.n28 a_n3134_n1088# 0.047009f
C101 minus.n29 a_n3134_n1088# 0.047119f
C102 minus.n30 a_n3134_n1088# 0.073455f
C103 minus.n31 a_n3134_n1088# 0.008013f
C104 minus.t12 a_n3134_n1088# 0.071845f
C105 minus.n32 a_n3134_n1088# 0.072802f
C106 minus.n33 a_n3134_n1088# 1.06731f
C107 minus.n34 a_n3134_n1088# 0.035312f
C108 minus.t16 a_n3134_n1088# 0.071845f
C109 minus.n35 a_n3134_n1088# 0.081141f
C110 minus.n36 a_n3134_n1088# 0.035312f
C111 minus.n37 a_n3134_n1088# 0.008013f
C112 minus.n38 a_n3134_n1088# 0.035312f
C113 minus.n39 a_n3134_n1088# 0.008013f
C114 minus.n40 a_n3134_n1088# 0.035312f
C115 minus.t7 a_n3134_n1088# 0.071845f
C116 minus.n41 a_n3134_n1088# 0.081141f
C117 minus.t23 a_n3134_n1088# 0.086439f
C118 minus.t10 a_n3134_n1088# 0.071845f
C119 minus.n42 a_n3134_n1088# 0.080681f
C120 minus.n43 a_n3134_n1088# 0.060037f
C121 minus.n44 a_n3134_n1088# 0.170892f
C122 minus.n45 a_n3134_n1088# 0.047119f
C123 minus.t22 a_n3134_n1088# 0.071845f
C124 minus.n46 a_n3134_n1088# 0.073673f
C125 minus.n47 a_n3134_n1088# 0.008013f
C126 minus.t17 a_n3134_n1088# 0.071845f
C127 minus.n48 a_n3134_n1088# 0.074652f
C128 minus.n49 a_n3134_n1088# 0.035312f
C129 minus.n50 a_n3134_n1088# 0.035312f
C130 minus.n51 a_n3134_n1088# 0.035312f
C131 minus.t21 a_n3134_n1088# 0.071845f
C132 minus.n52 a_n3134_n1088# 0.074652f
C133 minus.n53 a_n3134_n1088# 0.008013f
C134 minus.t9 a_n3134_n1088# 0.071845f
C135 minus.n54 a_n3134_n1088# 0.074652f
C136 minus.n55 a_n3134_n1088# 0.035312f
C137 minus.n56 a_n3134_n1088# 0.035312f
C138 minus.n57 a_n3134_n1088# 0.035312f
C139 minus.t5 a_n3134_n1088# 0.071845f
C140 minus.n58 a_n3134_n1088# 0.074652f
C141 minus.n59 a_n3134_n1088# 0.008013f
C142 minus.t20 a_n3134_n1088# 0.071845f
C143 minus.n60 a_n3134_n1088# 0.073673f
C144 minus.n61 a_n3134_n1088# 0.047119f
C145 minus.n62 a_n3134_n1088# 0.047009f
C146 minus.n63 a_n3134_n1088# 0.047119f
C147 minus.t19 a_n3134_n1088# 0.071845f
C148 minus.n64 a_n3134_n1088# 0.073455f
C149 minus.n65 a_n3134_n1088# 0.008013f
C150 minus.t8 a_n3134_n1088# 0.071845f
C151 minus.n66 a_n3134_n1088# 0.072802f
C152 minus.n67 a_n3134_n1088# 0.239367f
C153 minus.n68 a_n3134_n1088# 1.30534f
C154 drain_left.t15 a_n3134_n1088# 0.022102f
C155 drain_left.t13 a_n3134_n1088# 0.022102f
C156 drain_left.n0 a_n3134_n1088# 0.08705f
C157 drain_left.t16 a_n3134_n1088# 0.022102f
C158 drain_left.t7 a_n3134_n1088# 0.022102f
C159 drain_left.n1 a_n3134_n1088# 0.085881f
C160 drain_left.n2 a_n3134_n1088# 0.690285f
C161 drain_left.t1 a_n3134_n1088# 0.022102f
C162 drain_left.t22 a_n3134_n1088# 0.022102f
C163 drain_left.n3 a_n3134_n1088# 0.085881f
C164 drain_left.n4 a_n3134_n1088# 0.300857f
C165 drain_left.t19 a_n3134_n1088# 0.022102f
C166 drain_left.t11 a_n3134_n1088# 0.022102f
C167 drain_left.n5 a_n3134_n1088# 0.08705f
C168 drain_left.t2 a_n3134_n1088# 0.022102f
C169 drain_left.t0 a_n3134_n1088# 0.022102f
C170 drain_left.n6 a_n3134_n1088# 0.085881f
C171 drain_left.n7 a_n3134_n1088# 0.690285f
C172 drain_left.t14 a_n3134_n1088# 0.022102f
C173 drain_left.t9 a_n3134_n1088# 0.022102f
C174 drain_left.n8 a_n3134_n1088# 0.085881f
C175 drain_left.n9 a_n3134_n1088# 0.300857f
C176 drain_left.n10 a_n3134_n1088# 1.12565f
C177 drain_left.t4 a_n3134_n1088# 0.022102f
C178 drain_left.t5 a_n3134_n1088# 0.022102f
C179 drain_left.n11 a_n3134_n1088# 0.08705f
C180 drain_left.t8 a_n3134_n1088# 0.022102f
C181 drain_left.t10 a_n3134_n1088# 0.022102f
C182 drain_left.n12 a_n3134_n1088# 0.085881f
C183 drain_left.n13 a_n3134_n1088# 0.690284f
C184 drain_left.t12 a_n3134_n1088# 0.022102f
C185 drain_left.t17 a_n3134_n1088# 0.022102f
C186 drain_left.n14 a_n3134_n1088# 0.085881f
C187 drain_left.n15 a_n3134_n1088# 0.340094f
C188 drain_left.t18 a_n3134_n1088# 0.022102f
C189 drain_left.t20 a_n3134_n1088# 0.022102f
C190 drain_left.n16 a_n3134_n1088# 0.085881f
C191 drain_left.n17 a_n3134_n1088# 0.340094f
C192 drain_left.t21 a_n3134_n1088# 0.022102f
C193 drain_left.t23 a_n3134_n1088# 0.022102f
C194 drain_left.n18 a_n3134_n1088# 0.085881f
C195 drain_left.n19 a_n3134_n1088# 0.340094f
C196 drain_left.t3 a_n3134_n1088# 0.022102f
C197 drain_left.t6 a_n3134_n1088# 0.022102f
C198 drain_left.n20 a_n3134_n1088# 0.085881f
C199 drain_left.n21 a_n3134_n1088# 0.58398f
C200 source.t30 a_n3134_n1088# 0.164354f
C201 source.n0 a_n3134_n1088# 0.761368f
C202 source.t40 a_n3134_n1088# 0.029529f
C203 source.t38 a_n3134_n1088# 0.029529f
C204 source.n1 a_n3134_n1088# 0.095767f
C205 source.n2 a_n3134_n1088# 0.422565f
C206 source.t39 a_n3134_n1088# 0.029529f
C207 source.t42 a_n3134_n1088# 0.029529f
C208 source.n3 a_n3134_n1088# 0.095767f
C209 source.n4 a_n3134_n1088# 0.422565f
C210 source.t45 a_n3134_n1088# 0.029529f
C211 source.t25 a_n3134_n1088# 0.029529f
C212 source.n5 a_n3134_n1088# 0.095767f
C213 source.n6 a_n3134_n1088# 0.422565f
C214 source.t32 a_n3134_n1088# 0.029529f
C215 source.t35 a_n3134_n1088# 0.029529f
C216 source.n7 a_n3134_n1088# 0.095767f
C217 source.n8 a_n3134_n1088# 0.422565f
C218 source.t44 a_n3134_n1088# 0.029529f
C219 source.t33 a_n3134_n1088# 0.029529f
C220 source.n9 a_n3134_n1088# 0.095767f
C221 source.n10 a_n3134_n1088# 0.422565f
C222 source.t37 a_n3134_n1088# 0.164354f
C223 source.n11 a_n3134_n1088# 0.39455f
C224 source.t2 a_n3134_n1088# 0.164354f
C225 source.n12 a_n3134_n1088# 0.39455f
C226 source.t0 a_n3134_n1088# 0.029529f
C227 source.t20 a_n3134_n1088# 0.029529f
C228 source.n13 a_n3134_n1088# 0.095767f
C229 source.n14 a_n3134_n1088# 0.422565f
C230 source.t21 a_n3134_n1088# 0.029529f
C231 source.t12 a_n3134_n1088# 0.029529f
C232 source.n15 a_n3134_n1088# 0.095767f
C233 source.n16 a_n3134_n1088# 0.422565f
C234 source.t7 a_n3134_n1088# 0.029529f
C235 source.t17 a_n3134_n1088# 0.029529f
C236 source.n17 a_n3134_n1088# 0.095767f
C237 source.n18 a_n3134_n1088# 0.422565f
C238 source.t22 a_n3134_n1088# 0.029529f
C239 source.t5 a_n3134_n1088# 0.029529f
C240 source.n19 a_n3134_n1088# 0.095767f
C241 source.n20 a_n3134_n1088# 0.422565f
C242 source.t9 a_n3134_n1088# 0.029529f
C243 source.t18 a_n3134_n1088# 0.029529f
C244 source.n21 a_n3134_n1088# 0.095767f
C245 source.n22 a_n3134_n1088# 0.422565f
C246 source.t16 a_n3134_n1088# 0.164354f
C247 source.n23 a_n3134_n1088# 1.06742f
C248 source.t47 a_n3134_n1088# 0.164354f
C249 source.n24 a_n3134_n1088# 1.06742f
C250 source.t34 a_n3134_n1088# 0.029529f
C251 source.t29 a_n3134_n1088# 0.029529f
C252 source.n25 a_n3134_n1088# 0.095767f
C253 source.n26 a_n3134_n1088# 0.422566f
C254 source.t27 a_n3134_n1088# 0.029529f
C255 source.t26 a_n3134_n1088# 0.029529f
C256 source.n27 a_n3134_n1088# 0.095767f
C257 source.n28 a_n3134_n1088# 0.422566f
C258 source.t41 a_n3134_n1088# 0.029529f
C259 source.t46 a_n3134_n1088# 0.029529f
C260 source.n29 a_n3134_n1088# 0.095767f
C261 source.n30 a_n3134_n1088# 0.422566f
C262 source.t24 a_n3134_n1088# 0.029529f
C263 source.t28 a_n3134_n1088# 0.029529f
C264 source.n31 a_n3134_n1088# 0.095767f
C265 source.n32 a_n3134_n1088# 0.422566f
C266 source.t36 a_n3134_n1088# 0.029529f
C267 source.t31 a_n3134_n1088# 0.029529f
C268 source.n33 a_n3134_n1088# 0.095767f
C269 source.n34 a_n3134_n1088# 0.422566f
C270 source.t43 a_n3134_n1088# 0.164354f
C271 source.n35 a_n3134_n1088# 0.39455f
C272 source.t19 a_n3134_n1088# 0.164354f
C273 source.n36 a_n3134_n1088# 0.39455f
C274 source.t6 a_n3134_n1088# 0.029529f
C275 source.t4 a_n3134_n1088# 0.029529f
C276 source.n37 a_n3134_n1088# 0.095767f
C277 source.n38 a_n3134_n1088# 0.422566f
C278 source.t23 a_n3134_n1088# 0.029529f
C279 source.t15 a_n3134_n1088# 0.029529f
C280 source.n39 a_n3134_n1088# 0.095767f
C281 source.n40 a_n3134_n1088# 0.422566f
C282 source.t8 a_n3134_n1088# 0.029529f
C283 source.t3 a_n3134_n1088# 0.029529f
C284 source.n41 a_n3134_n1088# 0.095767f
C285 source.n42 a_n3134_n1088# 0.422566f
C286 source.t13 a_n3134_n1088# 0.029529f
C287 source.t14 a_n3134_n1088# 0.029529f
C288 source.n43 a_n3134_n1088# 0.095767f
C289 source.n44 a_n3134_n1088# 0.422566f
C290 source.t11 a_n3134_n1088# 0.029529f
C291 source.t10 a_n3134_n1088# 0.029529f
C292 source.n45 a_n3134_n1088# 0.095767f
C293 source.n46 a_n3134_n1088# 0.422566f
C294 source.t1 a_n3134_n1088# 0.164354f
C295 source.n47 a_n3134_n1088# 0.630166f
C296 source.n48 a_n3134_n1088# 0.76988f
C297 plus.n0 a_n3134_n1088# 0.045363f
C298 plus.t17 a_n3134_n1088# 0.092295f
C299 plus.t20 a_n3134_n1088# 0.092295f
C300 plus.n1 a_n3134_n1088# 0.060531f
C301 plus.t0 a_n3134_n1088# 0.092295f
C302 plus.n2 a_n3134_n1088# 0.060389f
C303 plus.t2 a_n3134_n1088# 0.092295f
C304 plus.n3 a_n3134_n1088# 0.060531f
C305 plus.t3 a_n3134_n1088# 0.092295f
C306 plus.n4 a_n3134_n1088# 0.095901f
C307 plus.n5 a_n3134_n1088# 0.045363f
C308 plus.t5 a_n3134_n1088# 0.092295f
C309 plus.t6 a_n3134_n1088# 0.092295f
C310 plus.n6 a_n3134_n1088# 0.095901f
C311 plus.n7 a_n3134_n1088# 0.045363f
C312 plus.t11 a_n3134_n1088# 0.092295f
C313 plus.t13 a_n3134_n1088# 0.092295f
C314 plus.n8 a_n3134_n1088# 0.094643f
C315 plus.t19 a_n3134_n1088# 0.111043f
C316 plus.n9 a_n3134_n1088# 0.077126f
C317 plus.t15 a_n3134_n1088# 0.092295f
C318 plus.t18 a_n3134_n1088# 0.092295f
C319 plus.n10 a_n3134_n1088# 0.103646f
C320 plus.n11 a_n3134_n1088# 0.104237f
C321 plus.n12 a_n3134_n1088# 0.219535f
C322 plus.n13 a_n3134_n1088# 0.060531f
C323 plus.n14 a_n3134_n1088# 0.045363f
C324 plus.n15 a_n3134_n1088# 0.010294f
C325 plus.n16 a_n3134_n1088# 0.095901f
C326 plus.n17 a_n3134_n1088# 0.010294f
C327 plus.n18 a_n3134_n1088# 0.045363f
C328 plus.n19 a_n3134_n1088# 0.045363f
C329 plus.n20 a_n3134_n1088# 0.045363f
C330 plus.n21 a_n3134_n1088# 0.010294f
C331 plus.n22 a_n3134_n1088# 0.095901f
C332 plus.n23 a_n3134_n1088# 0.010294f
C333 plus.n24 a_n3134_n1088# 0.045363f
C334 plus.n25 a_n3134_n1088# 0.045363f
C335 plus.n26 a_n3134_n1088# 0.045363f
C336 plus.n27 a_n3134_n1088# 0.010294f
C337 plus.n28 a_n3134_n1088# 0.094643f
C338 plus.n29 a_n3134_n1088# 0.104237f
C339 plus.n30 a_n3134_n1088# 0.094363f
C340 plus.n31 a_n3134_n1088# 0.010294f
C341 plus.n32 a_n3134_n1088# 0.093524f
C342 plus.n33 a_n3134_n1088# 0.32253f
C343 plus.n34 a_n3134_n1088# 0.045363f
C344 plus.t8 a_n3134_n1088# 0.092295f
C345 plus.n35 a_n3134_n1088# 0.060531f
C346 plus.t10 a_n3134_n1088# 0.092295f
C347 plus.n36 a_n3134_n1088# 0.060389f
C348 plus.t7 a_n3134_n1088# 0.092295f
C349 plus.n37 a_n3134_n1088# 0.060531f
C350 plus.t16 a_n3134_n1088# 0.092295f
C351 plus.t22 a_n3134_n1088# 0.092295f
C352 plus.n38 a_n3134_n1088# 0.095901f
C353 plus.n39 a_n3134_n1088# 0.045363f
C354 plus.t1 a_n3134_n1088# 0.092295f
C355 plus.t9 a_n3134_n1088# 0.092295f
C356 plus.n40 a_n3134_n1088# 0.095901f
C357 plus.n41 a_n3134_n1088# 0.045363f
C358 plus.t14 a_n3134_n1088# 0.092295f
C359 plus.t21 a_n3134_n1088# 0.092295f
C360 plus.n42 a_n3134_n1088# 0.094643f
C361 plus.t12 a_n3134_n1088# 0.111043f
C362 plus.n43 a_n3134_n1088# 0.077126f
C363 plus.t23 a_n3134_n1088# 0.092295f
C364 plus.t4 a_n3134_n1088# 0.092295f
C365 plus.n44 a_n3134_n1088# 0.103646f
C366 plus.n45 a_n3134_n1088# 0.104237f
C367 plus.n46 a_n3134_n1088# 0.219535f
C368 plus.n47 a_n3134_n1088# 0.060531f
C369 plus.n48 a_n3134_n1088# 0.045363f
C370 plus.n49 a_n3134_n1088# 0.010294f
C371 plus.n50 a_n3134_n1088# 0.095901f
C372 plus.n51 a_n3134_n1088# 0.010294f
C373 plus.n52 a_n3134_n1088# 0.045363f
C374 plus.n53 a_n3134_n1088# 0.045363f
C375 plus.n54 a_n3134_n1088# 0.045363f
C376 plus.n55 a_n3134_n1088# 0.010294f
C377 plus.n56 a_n3134_n1088# 0.095901f
C378 plus.n57 a_n3134_n1088# 0.010294f
C379 plus.n58 a_n3134_n1088# 0.045363f
C380 plus.n59 a_n3134_n1088# 0.045363f
C381 plus.n60 a_n3134_n1088# 0.045363f
C382 plus.n61 a_n3134_n1088# 0.010294f
C383 plus.n62 a_n3134_n1088# 0.094643f
C384 plus.n63 a_n3134_n1088# 0.104237f
C385 plus.n64 a_n3134_n1088# 0.094363f
C386 plus.n65 a_n3134_n1088# 0.010294f
C387 plus.n66 a_n3134_n1088# 0.093524f
C388 plus.n67 a_n3134_n1088# 1.31985f
.ends

