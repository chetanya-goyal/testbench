* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right.t1 minus.t0 source.t3 a_n1128_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.39 ps=2.78 w=1 l=0.7
X1 a_n1128_n1092# a_n1128_n1092# a_n1128_n1092# a_n1128_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.7
X2 a_n1128_n1092# a_n1128_n1092# a_n1128_n1092# a_n1128_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X3 drain_left.t1 plus.t0 source.t0 a_n1128_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.39 ps=2.78 w=1 l=0.7
X4 drain_right.t0 minus.t1 source.t2 a_n1128_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.39 ps=2.78 w=1 l=0.7
X5 a_n1128_n1092# a_n1128_n1092# a_n1128_n1092# a_n1128_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X6 a_n1128_n1092# a_n1128_n1092# a_n1128_n1092# a_n1128_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X7 drain_left.t0 plus.t1 source.t1 a_n1128_n1092# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.39 ps=2.78 w=1 l=0.7
R0 minus.n0 minus.t0 277.038
R1 minus.n0 minus.t1 258.464
R2 minus minus.n0 0.188
R3 source.n0 source.t0 243.255
R4 source.n1 source.t3 243.255
R5 source.n3 source.t2 243.254
R6 source.n2 source.t1 243.254
R7 source.n2 source.n1 14.7454
R8 source.n4 source.n0 8.15058
R9 source.n4 source.n3 5.7074
R10 source.n1 source.n0 0.914293
R11 source.n3 source.n2 0.914293
R12 source source.n4 0.188
R13 drain_right drain_right.t0 279.704
R14 drain_right drain_right.t1 266.029
R15 plus plus.t1 275.087
R16 plus plus.t0 259.94
R17 drain_left drain_left.t0 280.257
R18 drain_left drain_left.t1 266.474
C0 drain_left minus 0.179499f
C1 source plus 0.523143f
C2 drain_right source 1.65551f
C3 drain_left plus 0.49308f
C4 drain_right drain_left 0.458259f
C5 minus plus 2.51401f
C6 drain_right minus 0.388799f
C7 drain_right plus 0.267937f
C8 source drain_left 1.65638f
C9 source minus 0.509238f
C10 drain_right a_n1128_n1092# 1.70022f
C11 drain_left a_n1128_n1092# 1.80529f
C12 source a_n1128_n1092# 1.8893f
C13 minus a_n1128_n1092# 3.249432f
C14 plus a_n1128_n1092# 5.16154f
C15 plus.t0 a_n1128_n1092# 0.17512f
C16 plus.t1 a_n1128_n1092# 0.236801f
C17 minus.t0 a_n1128_n1092# 0.235394f
C18 minus.t1 a_n1128_n1092# 0.166919f
C19 minus.n0 a_n1128_n1092# 2.07003f
.ends

