* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t9 plus.t0 source.t18 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X1 drain_right.t9 minus.t0 source.t9 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X2 a_n1472_n1088# a_n1472_n1088# a_n1472_n1088# a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.3
X3 drain_right.t8 minus.t1 source.t8 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X4 source.t10 plus.t1 drain_left.t8 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X5 drain_left.t7 plus.t2 source.t11 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X6 source.t6 minus.t2 drain_right.t7 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X7 drain_left.t6 plus.t3 source.t13 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X8 drain_right.t6 minus.t3 source.t7 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X9 drain_left.t5 plus.t4 source.t12 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X10 source.t15 plus.t5 drain_left.t4 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X11 a_n1472_n1088# a_n1472_n1088# a_n1472_n1088# a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X12 drain_left.t3 plus.t6 source.t17 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X13 source.t2 minus.t4 drain_right.t5 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X14 a_n1472_n1088# a_n1472_n1088# a_n1472_n1088# a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X15 a_n1472_n1088# a_n1472_n1088# a_n1472_n1088# a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X16 drain_right.t4 minus.t5 source.t3 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X17 drain_right.t3 minus.t6 source.t5 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X18 source.t14 plus.t7 drain_left.t2 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X19 drain_left.t1 plus.t8 source.t16 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X20 source.t0 minus.t7 drain_right.t2 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X21 drain_right.t1 minus.t8 source.t4 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X22 source.t1 minus.t9 drain_right.t0 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X23 source.t19 plus.t9 drain_left.t0 a_n1472_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
R0 plus.n3 plus.t2 222.743
R1 plus.n9 plus.t4 222.743
R2 plus.n14 plus.t6 222.743
R3 plus.n20 plus.t3 222.743
R4 plus.n6 plus.t8 184.768
R5 plus.n2 plus.t5 184.768
R6 plus.n8 plus.t9 184.768
R7 plus.n17 plus.t0 184.768
R8 plus.n13 plus.t1 184.768
R9 plus.n19 plus.t7 184.768
R10 plus.n4 plus.n3 161.489
R11 plus.n15 plus.n14 161.489
R12 plus.n4 plus.n1 161.3
R13 plus.n6 plus.n5 161.3
R14 plus.n7 plus.n0 161.3
R15 plus.n10 plus.n9 161.3
R16 plus.n15 plus.n12 161.3
R17 plus.n17 plus.n16 161.3
R18 plus.n18 plus.n11 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n6 plus.n1 73.0308
R21 plus.n7 plus.n6 73.0308
R22 plus.n18 plus.n17 73.0308
R23 plus.n17 plus.n12 73.0308
R24 plus.n3 plus.n2 54.0429
R25 plus.n9 plus.n8 54.0429
R26 plus.n20 plus.n19 54.0429
R27 plus.n14 plus.n13 54.0429
R28 plus plus.n21 24.3986
R29 plus.n2 plus.n1 18.9884
R30 plus.n8 plus.n7 18.9884
R31 plus.n19 plus.n18 18.9884
R32 plus.n13 plus.n12 18.9884
R33 plus plus.n10 7.96452
R34 plus.n5 plus.n4 0.189894
R35 plus.n5 plus.n0 0.189894
R36 plus.n10 plus.n0 0.189894
R37 plus.n21 plus.n11 0.189894
R38 plus.n16 plus.n11 0.189894
R39 plus.n16 plus.n15 0.189894
R40 source.n0 source.t12 243.255
R41 source.n5 source.t3 243.255
R42 source.n19 source.t7 243.254
R43 source.n14 source.t17 243.254
R44 source.n2 source.n1 223.454
R45 source.n4 source.n3 223.454
R46 source.n7 source.n6 223.454
R47 source.n9 source.n8 223.454
R48 source.n18 source.n17 223.453
R49 source.n16 source.n15 223.453
R50 source.n13 source.n12 223.453
R51 source.n11 source.n10 223.453
R52 source.n17 source.t8 19.8005
R53 source.n17 source.t0 19.8005
R54 source.n15 source.t5 19.8005
R55 source.n15 source.t6 19.8005
R56 source.n12 source.t18 19.8005
R57 source.n12 source.t10 19.8005
R58 source.n10 source.t13 19.8005
R59 source.n10 source.t14 19.8005
R60 source.n1 source.t16 19.8005
R61 source.n1 source.t19 19.8005
R62 source.n3 source.t11 19.8005
R63 source.n3 source.t15 19.8005
R64 source.n6 source.t9 19.8005
R65 source.n6 source.t1 19.8005
R66 source.n8 source.t4 19.8005
R67 source.n8 source.t2 19.8005
R68 source.n11 source.n9 14.0406
R69 source.n20 source.n0 7.96301
R70 source.n20 source.n19 5.53498
R71 source.n5 source.n4 0.741879
R72 source.n16 source.n14 0.741879
R73 source.n9 source.n7 0.543603
R74 source.n7 source.n5 0.543603
R75 source.n4 source.n2 0.543603
R76 source.n2 source.n0 0.543603
R77 source.n13 source.n11 0.543603
R78 source.n14 source.n13 0.543603
R79 source.n18 source.n16 0.543603
R80 source.n19 source.n18 0.543603
R81 source source.n20 0.188
R82 drain_left.n5 drain_left.t7 260.476
R83 drain_left.n1 drain_left.t6 260.474
R84 drain_left.n3 drain_left.n2 240.483
R85 drain_left.n7 drain_left.n6 240.132
R86 drain_left.n5 drain_left.n4 240.132
R87 drain_left.n1 drain_left.n0 240.131
R88 drain_left drain_left.n3 21.3419
R89 drain_left.n2 drain_left.t8 19.8005
R90 drain_left.n2 drain_left.t3 19.8005
R91 drain_left.n0 drain_left.t2 19.8005
R92 drain_left.n0 drain_left.t9 19.8005
R93 drain_left.n6 drain_left.t0 19.8005
R94 drain_left.n6 drain_left.t5 19.8005
R95 drain_left.n4 drain_left.t4 19.8005
R96 drain_left.n4 drain_left.t1 19.8005
R97 drain_left drain_left.n7 6.19632
R98 drain_left.n7 drain_left.n5 0.543603
R99 drain_left.n3 drain_left.n1 0.0809298
R100 minus.n9 minus.t8 222.743
R101 minus.n3 minus.t5 222.743
R102 minus.n20 minus.t3 222.743
R103 minus.n14 minus.t6 222.743
R104 minus.n6 minus.t0 184.768
R105 minus.n8 minus.t4 184.768
R106 minus.n2 minus.t9 184.768
R107 minus.n17 minus.t1 184.768
R108 minus.n19 minus.t7 184.768
R109 minus.n13 minus.t2 184.768
R110 minus.n4 minus.n3 161.489
R111 minus.n15 minus.n14 161.489
R112 minus.n10 minus.n9 161.3
R113 minus.n7 minus.n0 161.3
R114 minus.n6 minus.n5 161.3
R115 minus.n4 minus.n1 161.3
R116 minus.n21 minus.n20 161.3
R117 minus.n18 minus.n11 161.3
R118 minus.n17 minus.n16 161.3
R119 minus.n15 minus.n12 161.3
R120 minus.n7 minus.n6 73.0308
R121 minus.n6 minus.n1 73.0308
R122 minus.n17 minus.n12 73.0308
R123 minus.n18 minus.n17 73.0308
R124 minus.n9 minus.n8 54.0429
R125 minus.n3 minus.n2 54.0429
R126 minus.n14 minus.n13 54.0429
R127 minus.n20 minus.n19 54.0429
R128 minus.n22 minus.n10 26.3509
R129 minus.n8 minus.n7 18.9884
R130 minus.n2 minus.n1 18.9884
R131 minus.n13 minus.n12 18.9884
R132 minus.n19 minus.n18 18.9884
R133 minus.n22 minus.n21 6.48724
R134 minus.n10 minus.n0 0.189894
R135 minus.n5 minus.n0 0.189894
R136 minus.n5 minus.n4 0.189894
R137 minus.n16 minus.n15 0.189894
R138 minus.n16 minus.n11 0.189894
R139 minus.n21 minus.n11 0.189894
R140 minus minus.n22 0.188
R141 drain_right.n1 drain_right.t3 260.474
R142 drain_right.n7 drain_right.t1 259.933
R143 drain_right.n6 drain_right.n4 240.675
R144 drain_right.n3 drain_right.n2 240.483
R145 drain_right.n6 drain_right.n5 240.132
R146 drain_right.n1 drain_right.n0 240.131
R147 drain_right drain_right.n3 20.7887
R148 drain_right.n2 drain_right.t2 19.8005
R149 drain_right.n2 drain_right.t6 19.8005
R150 drain_right.n0 drain_right.t7 19.8005
R151 drain_right.n0 drain_right.t8 19.8005
R152 drain_right.n4 drain_right.t0 19.8005
R153 drain_right.n4 drain_right.t4 19.8005
R154 drain_right.n5 drain_right.t5 19.8005
R155 drain_right.n5 drain_right.t9 19.8005
R156 drain_right drain_right.n7 5.92477
R157 drain_right.n7 drain_right.n6 0.543603
R158 drain_right.n3 drain_right.n1 0.0809298
C0 drain_right minus 0.693317f
C1 source plus 0.912033f
C2 plus minus 2.96011f
C3 drain_right plus 0.303523f
C4 source drain_left 3.72007f
C5 minus drain_left 0.179062f
C6 drain_right drain_left 0.720388f
C7 source minus 0.898115f
C8 drain_right source 3.71795f
C9 plus drain_left 0.833428f
C10 drain_right a_n1472_n1088# 3.1787f
C11 drain_left a_n1472_n1088# 3.38267f
C12 source a_n1472_n1088# 2.03066f
C13 minus a_n1472_n1088# 4.79854f
C14 plus a_n1472_n1088# 5.501058f
C15 drain_right.t3 a_n1472_n1088# 0.111767f
C16 drain_right.t7 a_n1472_n1088# 0.017997f
C17 drain_right.t8 a_n1472_n1088# 0.017997f
C18 drain_right.n0 a_n1472_n1088# 0.069929f
C19 drain_right.n1 a_n1472_n1088# 0.427112f
C20 drain_right.t2 a_n1472_n1088# 0.017997f
C21 drain_right.t6 a_n1472_n1088# 0.017997f
C22 drain_right.n2 a_n1472_n1088# 0.070274f
C23 drain_right.n3 a_n1472_n1088# 0.718362f
C24 drain_right.t0 a_n1472_n1088# 0.017997f
C25 drain_right.t4 a_n1472_n1088# 0.017997f
C26 drain_right.n4 a_n1472_n1088# 0.070489f
C27 drain_right.t5 a_n1472_n1088# 0.017997f
C28 drain_right.t9 a_n1472_n1088# 0.017997f
C29 drain_right.n5 a_n1472_n1088# 0.069929f
C30 drain_right.n6 a_n1472_n1088# 0.486549f
C31 drain_right.t1 a_n1472_n1088# 0.111316f
C32 drain_right.n7 a_n1472_n1088# 0.405972f
C33 minus.n0 a_n1472_n1088# 0.035436f
C34 minus.t8 a_n1472_n1088# 0.038752f
C35 minus.t4 a_n1472_n1088# 0.032772f
C36 minus.t0 a_n1472_n1088# 0.032772f
C37 minus.n1 a_n1472_n1088# 0.014596f
C38 minus.t9 a_n1472_n1088# 0.032772f
C39 minus.n2 a_n1472_n1088# 0.033765f
C40 minus.t5 a_n1472_n1088# 0.038752f
C41 minus.n3 a_n1472_n1088# 0.043741f
C42 minus.n4 a_n1472_n1088# 0.077814f
C43 minus.n5 a_n1472_n1088# 0.035436f
C44 minus.n6 a_n1472_n1088# 0.045521f
C45 minus.n7 a_n1472_n1088# 0.014596f
C46 minus.n8 a_n1472_n1088# 0.033765f
C47 minus.n9 a_n1472_n1088# 0.043692f
C48 minus.n10 a_n1472_n1088# 0.732532f
C49 minus.n11 a_n1472_n1088# 0.035436f
C50 minus.t7 a_n1472_n1088# 0.032772f
C51 minus.t1 a_n1472_n1088# 0.032772f
C52 minus.n12 a_n1472_n1088# 0.014596f
C53 minus.t6 a_n1472_n1088# 0.038752f
C54 minus.t2 a_n1472_n1088# 0.032772f
C55 minus.n13 a_n1472_n1088# 0.033765f
C56 minus.n14 a_n1472_n1088# 0.043741f
C57 minus.n15 a_n1472_n1088# 0.077814f
C58 minus.n16 a_n1472_n1088# 0.035436f
C59 minus.n17 a_n1472_n1088# 0.045521f
C60 minus.n18 a_n1472_n1088# 0.014596f
C61 minus.n19 a_n1472_n1088# 0.033765f
C62 minus.t3 a_n1472_n1088# 0.038752f
C63 minus.n20 a_n1472_n1088# 0.043692f
C64 minus.n21 a_n1472_n1088# 0.230608f
C65 minus.n22 a_n1472_n1088# 0.905225f
C66 drain_left.t6 a_n1472_n1088# 0.109139f
C67 drain_left.t2 a_n1472_n1088# 0.017574f
C68 drain_left.t9 a_n1472_n1088# 0.017574f
C69 drain_left.n0 a_n1472_n1088# 0.068285f
C70 drain_left.n1 a_n1472_n1088# 0.41707f
C71 drain_left.t8 a_n1472_n1088# 0.017574f
C72 drain_left.t3 a_n1472_n1088# 0.017574f
C73 drain_left.n2 a_n1472_n1088# 0.068622f
C74 drain_left.n3 a_n1472_n1088# 0.74456f
C75 drain_left.t7 a_n1472_n1088# 0.109139f
C76 drain_left.t4 a_n1472_n1088# 0.017574f
C77 drain_left.t1 a_n1472_n1088# 0.017574f
C78 drain_left.n4 a_n1472_n1088# 0.068285f
C79 drain_left.n5 a_n1472_n1088# 0.443813f
C80 drain_left.t0 a_n1472_n1088# 0.017574f
C81 drain_left.t5 a_n1472_n1088# 0.017574f
C82 drain_left.n6 a_n1472_n1088# 0.068285f
C83 drain_left.n7 a_n1472_n1088# 0.418453f
C84 source.t12 a_n1472_n1088# 0.133436f
C85 source.n0 a_n1472_n1088# 0.572954f
C86 source.t16 a_n1472_n1088# 0.023974f
C87 source.t19 a_n1472_n1088# 0.023974f
C88 source.n1 a_n1472_n1088# 0.077752f
C89 source.n2 a_n1472_n1088# 0.29251f
C90 source.t11 a_n1472_n1088# 0.023974f
C91 source.t15 a_n1472_n1088# 0.023974f
C92 source.n3 a_n1472_n1088# 0.077752f
C93 source.n4 a_n1472_n1088# 0.311892f
C94 source.t3 a_n1472_n1088# 0.133436f
C95 source.n5 a_n1472_n1088# 0.321592f
C96 source.t9 a_n1472_n1088# 0.023974f
C97 source.t1 a_n1472_n1088# 0.023974f
C98 source.n6 a_n1472_n1088# 0.077752f
C99 source.n7 a_n1472_n1088# 0.29251f
C100 source.t4 a_n1472_n1088# 0.023974f
C101 source.t2 a_n1472_n1088# 0.023974f
C102 source.n8 a_n1472_n1088# 0.077752f
C103 source.n9 a_n1472_n1088# 0.859446f
C104 source.t13 a_n1472_n1088# 0.023974f
C105 source.t14 a_n1472_n1088# 0.023974f
C106 source.n10 a_n1472_n1088# 0.077752f
C107 source.n11 a_n1472_n1088# 0.859446f
C108 source.t18 a_n1472_n1088# 0.023974f
C109 source.t10 a_n1472_n1088# 0.023974f
C110 source.n12 a_n1472_n1088# 0.077752f
C111 source.n13 a_n1472_n1088# 0.29251f
C112 source.t17 a_n1472_n1088# 0.133436f
C113 source.n14 a_n1472_n1088# 0.321592f
C114 source.t5 a_n1472_n1088# 0.023974f
C115 source.t6 a_n1472_n1088# 0.023974f
C116 source.n15 a_n1472_n1088# 0.077752f
C117 source.n16 a_n1472_n1088# 0.311893f
C118 source.t8 a_n1472_n1088# 0.023974f
C119 source.t0 a_n1472_n1088# 0.023974f
C120 source.n17 a_n1472_n1088# 0.077752f
C121 source.n18 a_n1472_n1088# 0.29251f
C122 source.t7 a_n1472_n1088# 0.133436f
C123 source.n19 a_n1472_n1088# 0.466304f
C124 source.n20 a_n1472_n1088# 0.614428f
C125 plus.n0 a_n1472_n1088# 0.036304f
C126 plus.t9 a_n1472_n1088# 0.033574f
C127 plus.t8 a_n1472_n1088# 0.033574f
C128 plus.n1 a_n1472_n1088# 0.014953f
C129 plus.t2 a_n1472_n1088# 0.039701f
C130 plus.t5 a_n1472_n1088# 0.033574f
C131 plus.n2 a_n1472_n1088# 0.034591f
C132 plus.n3 a_n1472_n1088# 0.044812f
C133 plus.n4 a_n1472_n1088# 0.079719f
C134 plus.n5 a_n1472_n1088# 0.036304f
C135 plus.n6 a_n1472_n1088# 0.046634f
C136 plus.n7 a_n1472_n1088# 0.014953f
C137 plus.n8 a_n1472_n1088# 0.034591f
C138 plus.t4 a_n1472_n1088# 0.039701f
C139 plus.n9 a_n1472_n1088# 0.044761f
C140 plus.n10 a_n1472_n1088# 0.247746f
C141 plus.n11 a_n1472_n1088# 0.036304f
C142 plus.t3 a_n1472_n1088# 0.039701f
C143 plus.t7 a_n1472_n1088# 0.033574f
C144 plus.t0 a_n1472_n1088# 0.033574f
C145 plus.n12 a_n1472_n1088# 0.014953f
C146 plus.t1 a_n1472_n1088# 0.033574f
C147 plus.n13 a_n1472_n1088# 0.034591f
C148 plus.t6 a_n1472_n1088# 0.039701f
C149 plus.n14 a_n1472_n1088# 0.044812f
C150 plus.n15 a_n1472_n1088# 0.079719f
C151 plus.n16 a_n1472_n1088# 0.036304f
C152 plus.n17 a_n1472_n1088# 0.046634f
C153 plus.n18 a_n1472_n1088# 0.014953f
C154 plus.n19 a_n1472_n1088# 0.034591f
C155 plus.n20 a_n1472_n1088# 0.044761f
C156 plus.n21 a_n1472_n1088# 0.731527f
.ends

