* NGSPICE file created from diffpair325.ext - technology: sky130A

.subckt diffpair325 minus drain_right drain_left source plus
X0 drain_left.t11 plus.t0 source.t20 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X1 source.t16 plus.t1 drain_left.t10 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X2 a_n1626_n2688# a_n1626_n2688# a_n1626_n2688# a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=34.2 ps=151.6 w=9 l=0.15
X3 source.t8 minus.t0 drain_right.t11 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X4 a_n1626_n2688# a_n1626_n2688# a_n1626_n2688# a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X5 drain_left.t9 plus.t2 source.t19 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X6 drain_right.t10 minus.t1 source.t6 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X7 drain_left.t8 plus.t3 source.t12 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X8 drain_right.t9 minus.t2 source.t11 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X9 source.t1 minus.t3 drain_right.t8 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X10 source.t21 plus.t4 drain_left.t7 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X11 drain_right.t7 minus.t4 source.t7 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X12 drain_right.t6 minus.t5 source.t10 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X13 a_n1626_n2688# a_n1626_n2688# a_n1626_n2688# a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X14 source.t9 minus.t6 drain_right.t5 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X15 source.t0 minus.t7 drain_right.t4 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X16 source.t22 plus.t5 drain_left.t6 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X17 drain_right.t3 minus.t8 source.t5 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X18 drain_left.t5 plus.t6 source.t14 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X19 source.t2 minus.t9 drain_right.t2 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X20 drain_right.t1 minus.t10 source.t4 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X21 source.t13 plus.t7 drain_left.t4 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X22 a_n1626_n2688# a_n1626_n2688# a_n1626_n2688# a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X23 drain_left.t3 plus.t8 source.t23 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X24 drain_left.t2 plus.t9 source.t17 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X25 source.t3 minus.t11 drain_right.t0 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X26 source.t15 plus.t10 drain_left.t1 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X27 source.t18 plus.t11 drain_left.t0 a_n1626_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
R0 plus.n2 plus.t5 1709.64
R1 plus.n13 plus.t8 1709.64
R2 plus.n17 plus.t2 1709.64
R3 plus.n28 plus.t10 1709.64
R4 plus.n3 plus.t9 1654.87
R5 plus.n4 plus.t7 1654.87
R6 plus.n10 plus.t6 1654.87
R7 plus.n12 plus.t11 1654.87
R8 plus.n19 plus.t4 1654.87
R9 plus.n18 plus.t0 1654.87
R10 plus.n25 plus.t1 1654.87
R11 plus.n27 plus.t3 1654.87
R12 plus.n6 plus.n2 161.489
R13 plus.n21 plus.n17 161.489
R14 plus.n6 plus.n5 161.3
R15 plus.n7 plus.n1 161.3
R16 plus.n9 plus.n8 161.3
R17 plus.n11 plus.n0 161.3
R18 plus.n14 plus.n13 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n22 plus.n16 161.3
R21 plus.n24 plus.n23 161.3
R22 plus.n26 plus.n15 161.3
R23 plus.n29 plus.n28 161.3
R24 plus.n9 plus.n1 73.0308
R25 plus.n24 plus.n16 73.0308
R26 plus.n5 plus.n4 62.0763
R27 plus.n11 plus.n10 62.0763
R28 plus.n26 plus.n25 62.0763
R29 plus.n20 plus.n18 62.0763
R30 plus.n3 plus.n2 40.1672
R31 plus.n13 plus.n12 40.1672
R32 plus.n28 plus.n27 40.1672
R33 plus.n19 plus.n17 40.1672
R34 plus.n5 plus.n3 32.8641
R35 plus.n12 plus.n11 32.8641
R36 plus.n27 plus.n26 32.8641
R37 plus.n20 plus.n19 32.8641
R38 plus plus.n29 28.0672
R39 plus plus.n14 11.0497
R40 plus.n4 plus.n1 10.955
R41 plus.n10 plus.n9 10.955
R42 plus.n25 plus.n24 10.955
R43 plus.n18 plus.n16 10.955
R44 plus.n7 plus.n6 0.189894
R45 plus.n8 plus.n7 0.189894
R46 plus.n8 plus.n0 0.189894
R47 plus.n14 plus.n0 0.189894
R48 plus.n29 plus.n15 0.189894
R49 plus.n23 plus.n15 0.189894
R50 plus.n23 plus.n22 0.189894
R51 plus.n22 plus.n21 0.189894
R52 source.n5 source.t22 52.1921
R53 source.n6 source.t7 52.1921
R54 source.n11 source.t2 52.1921
R55 source.n23 source.t11 52.1919
R56 source.n18 source.t3 52.1919
R57 source.n17 source.t19 52.1919
R58 source.n12 source.t15 52.1919
R59 source.n0 source.t23 52.1919
R60 source.n2 source.n1 48.8588
R61 source.n4 source.n3 48.8588
R62 source.n8 source.n7 48.8588
R63 source.n10 source.n9 48.8588
R64 source.n22 source.n21 48.8586
R65 source.n20 source.n19 48.8586
R66 source.n16 source.n15 48.8586
R67 source.n14 source.n13 48.8586
R68 source.n12 source.n11 19.5753
R69 source.n24 source.n0 14.0322
R70 source.n24 source.n23 5.5436
R71 source.n21 source.t4 3.33383
R72 source.n21 source.t8 3.33383
R73 source.n19 source.t6 3.33383
R74 source.n19 source.t9 3.33383
R75 source.n15 source.t20 3.33383
R76 source.n15 source.t21 3.33383
R77 source.n13 source.t12 3.33383
R78 source.n13 source.t16 3.33383
R79 source.n1 source.t14 3.33383
R80 source.n1 source.t18 3.33383
R81 source.n3 source.t17 3.33383
R82 source.n3 source.t13 3.33383
R83 source.n7 source.t5 3.33383
R84 source.n7 source.t1 3.33383
R85 source.n9 source.t10 3.33383
R86 source.n9 source.t0 3.33383
R87 source.n11 source.n10 0.560845
R88 source.n10 source.n8 0.560845
R89 source.n8 source.n6 0.560845
R90 source.n5 source.n4 0.560845
R91 source.n4 source.n2 0.560845
R92 source.n2 source.n0 0.560845
R93 source.n14 source.n12 0.560845
R94 source.n16 source.n14 0.560845
R95 source.n17 source.n16 0.560845
R96 source.n20 source.n18 0.560845
R97 source.n22 source.n20 0.560845
R98 source.n23 source.n22 0.560845
R99 source.n6 source.n5 0.470328
R100 source.n18 source.n17 0.470328
R101 source source.n24 0.188
R102 drain_left.n6 drain_left.n4 66.0979
R103 drain_left.n3 drain_left.n2 66.0423
R104 drain_left.n3 drain_left.n0 66.0423
R105 drain_left.n6 drain_left.n5 65.5376
R106 drain_left.n8 drain_left.n7 65.5374
R107 drain_left.n3 drain_left.n1 65.5373
R108 drain_left drain_left.n3 27.8961
R109 drain_left drain_left.n8 6.21356
R110 drain_left.n1 drain_left.t10 3.33383
R111 drain_left.n1 drain_left.t11 3.33383
R112 drain_left.n2 drain_left.t7 3.33383
R113 drain_left.n2 drain_left.t9 3.33383
R114 drain_left.n0 drain_left.t1 3.33383
R115 drain_left.n0 drain_left.t8 3.33383
R116 drain_left.n7 drain_left.t0 3.33383
R117 drain_left.n7 drain_left.t3 3.33383
R118 drain_left.n5 drain_left.t4 3.33383
R119 drain_left.n5 drain_left.t5 3.33383
R120 drain_left.n4 drain_left.t6 3.33383
R121 drain_left.n4 drain_left.t2 3.33383
R122 drain_left.n8 drain_left.n6 0.560845
R123 minus.n13 minus.t9 1709.64
R124 minus.n2 minus.t4 1709.64
R125 minus.n28 minus.t2 1709.64
R126 minus.n17 minus.t11 1709.64
R127 minus.n12 minus.t5 1654.87
R128 minus.n10 minus.t7 1654.87
R129 minus.n3 minus.t8 1654.87
R130 minus.n4 minus.t3 1654.87
R131 minus.n27 minus.t0 1654.87
R132 minus.n25 minus.t10 1654.87
R133 minus.n19 minus.t6 1654.87
R134 minus.n18 minus.t1 1654.87
R135 minus.n6 minus.n2 161.489
R136 minus.n21 minus.n17 161.489
R137 minus.n14 minus.n13 161.3
R138 minus.n11 minus.n0 161.3
R139 minus.n9 minus.n8 161.3
R140 minus.n7 minus.n1 161.3
R141 minus.n6 minus.n5 161.3
R142 minus.n29 minus.n28 161.3
R143 minus.n26 minus.n15 161.3
R144 minus.n24 minus.n23 161.3
R145 minus.n22 minus.n16 161.3
R146 minus.n21 minus.n20 161.3
R147 minus.n9 minus.n1 73.0308
R148 minus.n24 minus.n16 73.0308
R149 minus.n11 minus.n10 62.0763
R150 minus.n5 minus.n3 62.0763
R151 minus.n20 minus.n19 62.0763
R152 minus.n26 minus.n25 62.0763
R153 minus.n13 minus.n12 40.1672
R154 minus.n4 minus.n2 40.1672
R155 minus.n18 minus.n17 40.1672
R156 minus.n28 minus.n27 40.1672
R157 minus.n30 minus.n14 33.0497
R158 minus.n12 minus.n11 32.8641
R159 minus.n5 minus.n4 32.8641
R160 minus.n20 minus.n18 32.8641
R161 minus.n27 minus.n26 32.8641
R162 minus.n10 minus.n9 10.955
R163 minus.n3 minus.n1 10.955
R164 minus.n19 minus.n16 10.955
R165 minus.n25 minus.n24 10.955
R166 minus.n30 minus.n29 6.54217
R167 minus.n14 minus.n0 0.189894
R168 minus.n8 minus.n0 0.189894
R169 minus.n8 minus.n7 0.189894
R170 minus.n7 minus.n6 0.189894
R171 minus.n22 minus.n21 0.189894
R172 minus.n23 minus.n22 0.189894
R173 minus.n23 minus.n15 0.189894
R174 minus.n29 minus.n15 0.189894
R175 minus minus.n30 0.188
R176 drain_right.n6 drain_right.n4 66.0978
R177 drain_right.n3 drain_right.n2 66.0423
R178 drain_right.n3 drain_right.n0 66.0423
R179 drain_right.n6 drain_right.n5 65.5376
R180 drain_right.n8 drain_right.n7 65.5376
R181 drain_right.n3 drain_right.n1 65.5373
R182 drain_right drain_right.n3 27.3428
R183 drain_right drain_right.n8 6.21356
R184 drain_right.n1 drain_right.t5 3.33383
R185 drain_right.n1 drain_right.t1 3.33383
R186 drain_right.n2 drain_right.t11 3.33383
R187 drain_right.n2 drain_right.t9 3.33383
R188 drain_right.n0 drain_right.t0 3.33383
R189 drain_right.n0 drain_right.t10 3.33383
R190 drain_right.n4 drain_right.t8 3.33383
R191 drain_right.n4 drain_right.t7 3.33383
R192 drain_right.n5 drain_right.t4 3.33383
R193 drain_right.n5 drain_right.t3 3.33383
R194 drain_right.n7 drain_right.t2 3.33383
R195 drain_right.n7 drain_right.t6 3.33383
R196 drain_right.n8 drain_right.n6 0.560845
C0 minus plus 4.60818f
C1 source drain_right 18.605501f
C2 source minus 1.86883f
C3 source plus 1.88287f
C4 drain_right drain_left 0.801529f
C5 minus drain_left 0.170585f
C6 plus drain_left 2.4131f
C7 minus drain_right 2.25661f
C8 plus drain_right 0.309819f
C9 source drain_left 18.6057f
C10 drain_right a_n1626_n2688# 5.11734f
C11 drain_left a_n1626_n2688# 5.359651f
C12 source a_n1626_n2688# 7.04864f
C13 minus a_n1626_n2688# 5.770333f
C14 plus a_n1626_n2688# 7.249371f
C15 drain_right.t0 a_n1626_n2688# 0.302706f
C16 drain_right.t10 a_n1626_n2688# 0.302706f
C17 drain_right.n0 a_n1626_n2688# 1.95585f
C18 drain_right.t5 a_n1626_n2688# 0.302706f
C19 drain_right.t1 a_n1626_n2688# 0.302706f
C20 drain_right.n1 a_n1626_n2688# 1.9533f
C21 drain_right.t11 a_n1626_n2688# 0.302706f
C22 drain_right.t9 a_n1626_n2688# 0.302706f
C23 drain_right.n2 a_n1626_n2688# 1.95585f
C24 drain_right.n3 a_n1626_n2688# 2.00753f
C25 drain_right.t8 a_n1626_n2688# 0.302706f
C26 drain_right.t7 a_n1626_n2688# 0.302706f
C27 drain_right.n4 a_n1626_n2688# 1.95616f
C28 drain_right.t4 a_n1626_n2688# 0.302706f
C29 drain_right.t3 a_n1626_n2688# 0.302706f
C30 drain_right.n5 a_n1626_n2688# 1.9533f
C31 drain_right.n6 a_n1626_n2688# 0.661357f
C32 drain_right.t2 a_n1626_n2688# 0.302706f
C33 drain_right.t6 a_n1626_n2688# 0.302706f
C34 drain_right.n7 a_n1626_n2688# 1.9533f
C35 drain_right.n8 a_n1626_n2688# 0.56104f
C36 minus.n0 a_n1626_n2688# 0.04374f
C37 minus.t9 a_n1626_n2688# 0.169797f
C38 minus.t5 a_n1626_n2688# 0.167321f
C39 minus.t7 a_n1626_n2688# 0.167321f
C40 minus.n1 a_n1626_n2688# 0.016532f
C41 minus.t4 a_n1626_n2688# 0.169797f
C42 minus.n2 a_n1626_n2688# 0.093429f
C43 minus.t8 a_n1626_n2688# 0.167321f
C44 minus.n3 a_n1626_n2688# 0.076612f
C45 minus.t3 a_n1626_n2688# 0.167321f
C46 minus.n4 a_n1626_n2688# 0.076612f
C47 minus.n5 a_n1626_n2688# 0.018555f
C48 minus.n6 a_n1626_n2688# 0.098203f
C49 minus.n7 a_n1626_n2688# 0.04374f
C50 minus.n8 a_n1626_n2688# 0.04374f
C51 minus.n9 a_n1626_n2688# 0.016532f
C52 minus.n10 a_n1626_n2688# 0.076612f
C53 minus.n11 a_n1626_n2688# 0.018555f
C54 minus.n12 a_n1626_n2688# 0.076612f
C55 minus.n13 a_n1626_n2688# 0.093366f
C56 minus.n14 a_n1626_n2688# 1.33874f
C57 minus.n15 a_n1626_n2688# 0.04374f
C58 minus.t0 a_n1626_n2688# 0.167321f
C59 minus.t10 a_n1626_n2688# 0.167321f
C60 minus.n16 a_n1626_n2688# 0.016532f
C61 minus.t11 a_n1626_n2688# 0.169797f
C62 minus.n17 a_n1626_n2688# 0.093429f
C63 minus.t1 a_n1626_n2688# 0.167321f
C64 minus.n18 a_n1626_n2688# 0.076612f
C65 minus.t6 a_n1626_n2688# 0.167321f
C66 minus.n19 a_n1626_n2688# 0.076612f
C67 minus.n20 a_n1626_n2688# 0.018555f
C68 minus.n21 a_n1626_n2688# 0.098203f
C69 minus.n22 a_n1626_n2688# 0.04374f
C70 minus.n23 a_n1626_n2688# 0.04374f
C71 minus.n24 a_n1626_n2688# 0.016532f
C72 minus.n25 a_n1626_n2688# 0.076612f
C73 minus.n26 a_n1626_n2688# 0.018555f
C74 minus.n27 a_n1626_n2688# 0.076612f
C75 minus.t2 a_n1626_n2688# 0.169797f
C76 minus.n28 a_n1626_n2688# 0.093366f
C77 minus.n29 a_n1626_n2688# 0.290297f
C78 minus.n30 a_n1626_n2688# 1.63879f
C79 drain_left.t1 a_n1626_n2688# 0.302563f
C80 drain_left.t8 a_n1626_n2688# 0.302563f
C81 drain_left.n0 a_n1626_n2688# 1.95493f
C82 drain_left.t10 a_n1626_n2688# 0.302563f
C83 drain_left.t11 a_n1626_n2688# 0.302563f
C84 drain_left.n1 a_n1626_n2688# 1.95238f
C85 drain_left.t7 a_n1626_n2688# 0.302563f
C86 drain_left.t9 a_n1626_n2688# 0.302563f
C87 drain_left.n2 a_n1626_n2688# 1.95493f
C88 drain_left.n3 a_n1626_n2688# 2.06461f
C89 drain_left.t6 a_n1626_n2688# 0.302563f
C90 drain_left.t2 a_n1626_n2688# 0.302563f
C91 drain_left.n4 a_n1626_n2688# 1.95525f
C92 drain_left.t4 a_n1626_n2688# 0.302563f
C93 drain_left.t5 a_n1626_n2688# 0.302563f
C94 drain_left.n5 a_n1626_n2688# 1.95238f
C95 drain_left.n6 a_n1626_n2688# 0.661039f
C96 drain_left.t0 a_n1626_n2688# 0.302563f
C97 drain_left.t3 a_n1626_n2688# 0.302563f
C98 drain_left.n7 a_n1626_n2688# 1.95238f
C99 drain_left.n8 a_n1626_n2688# 0.560783f
C100 source.t23 a_n1626_n2688# 1.70733f
C101 source.n0 a_n1626_n2688# 0.952382f
C102 source.t14 a_n1626_n2688# 0.225907f
C103 source.t18 a_n1626_n2688# 0.225907f
C104 source.n1 a_n1626_n2688# 1.40177f
C105 source.n2 a_n1626_n2688# 0.271094f
C106 source.t17 a_n1626_n2688# 0.225907f
C107 source.t13 a_n1626_n2688# 0.225907f
C108 source.n3 a_n1626_n2688# 1.40177f
C109 source.n4 a_n1626_n2688# 0.271094f
C110 source.t22 a_n1626_n2688# 1.70734f
C111 source.n5 a_n1626_n2688# 0.366049f
C112 source.t7 a_n1626_n2688# 1.70734f
C113 source.n6 a_n1626_n2688# 0.366049f
C114 source.t5 a_n1626_n2688# 0.225907f
C115 source.t1 a_n1626_n2688# 0.225907f
C116 source.n7 a_n1626_n2688# 1.40177f
C117 source.n8 a_n1626_n2688# 0.271094f
C118 source.t10 a_n1626_n2688# 0.225907f
C119 source.t0 a_n1626_n2688# 0.225907f
C120 source.n9 a_n1626_n2688# 1.40177f
C121 source.n10 a_n1626_n2688# 0.271094f
C122 source.t2 a_n1626_n2688# 1.70734f
C123 source.n11 a_n1626_n2688# 1.25737f
C124 source.t15 a_n1626_n2688# 1.70733f
C125 source.n12 a_n1626_n2688# 1.25737f
C126 source.t12 a_n1626_n2688# 0.225907f
C127 source.t16 a_n1626_n2688# 0.225907f
C128 source.n13 a_n1626_n2688# 1.40177f
C129 source.n14 a_n1626_n2688# 0.271097f
C130 source.t20 a_n1626_n2688# 0.225907f
C131 source.t21 a_n1626_n2688# 0.225907f
C132 source.n15 a_n1626_n2688# 1.40177f
C133 source.n16 a_n1626_n2688# 0.271097f
C134 source.t19 a_n1626_n2688# 1.70733f
C135 source.n17 a_n1626_n2688# 0.366053f
C136 source.t3 a_n1626_n2688# 1.70733f
C137 source.n18 a_n1626_n2688# 0.366053f
C138 source.t6 a_n1626_n2688# 0.225907f
C139 source.t9 a_n1626_n2688# 0.225907f
C140 source.n19 a_n1626_n2688# 1.40177f
C141 source.n20 a_n1626_n2688# 0.271097f
C142 source.t4 a_n1626_n2688# 0.225907f
C143 source.t8 a_n1626_n2688# 0.225907f
C144 source.n21 a_n1626_n2688# 1.40177f
C145 source.n22 a_n1626_n2688# 0.271097f
C146 source.t11 a_n1626_n2688# 1.70733f
C147 source.n23 a_n1626_n2688# 0.485326f
C148 source.n24 a_n1626_n2688# 1.09195f
C149 plus.n0 a_n1626_n2688# 0.04495f
C150 plus.t11 a_n1626_n2688# 0.171951f
C151 plus.t6 a_n1626_n2688# 0.171951f
C152 plus.n1 a_n1626_n2688# 0.01699f
C153 plus.t5 a_n1626_n2688# 0.174495f
C154 plus.n2 a_n1626_n2688# 0.096014f
C155 plus.t9 a_n1626_n2688# 0.171951f
C156 plus.n3 a_n1626_n2688# 0.078732f
C157 plus.t7 a_n1626_n2688# 0.171951f
C158 plus.n4 a_n1626_n2688# 0.078732f
C159 plus.n5 a_n1626_n2688# 0.019069f
C160 plus.n6 a_n1626_n2688# 0.10092f
C161 plus.n7 a_n1626_n2688# 0.04495f
C162 plus.n8 a_n1626_n2688# 0.04495f
C163 plus.n9 a_n1626_n2688# 0.01699f
C164 plus.n10 a_n1626_n2688# 0.078732f
C165 plus.n11 a_n1626_n2688# 0.019069f
C166 plus.n12 a_n1626_n2688# 0.078732f
C167 plus.t8 a_n1626_n2688# 0.174495f
C168 plus.n13 a_n1626_n2688# 0.095949f
C169 plus.n14 a_n1626_n2688# 0.446136f
C170 plus.n15 a_n1626_n2688# 0.04495f
C171 plus.t10 a_n1626_n2688# 0.174495f
C172 plus.t3 a_n1626_n2688# 0.171951f
C173 plus.t1 a_n1626_n2688# 0.171951f
C174 plus.n16 a_n1626_n2688# 0.01699f
C175 plus.t2 a_n1626_n2688# 0.174495f
C176 plus.n17 a_n1626_n2688# 0.096014f
C177 plus.t0 a_n1626_n2688# 0.171951f
C178 plus.n18 a_n1626_n2688# 0.078732f
C179 plus.t4 a_n1626_n2688# 0.171951f
C180 plus.n19 a_n1626_n2688# 0.078732f
C181 plus.n20 a_n1626_n2688# 0.019069f
C182 plus.n21 a_n1626_n2688# 0.10092f
C183 plus.n22 a_n1626_n2688# 0.04495f
C184 plus.n23 a_n1626_n2688# 0.04495f
C185 plus.n24 a_n1626_n2688# 0.01699f
C186 plus.n25 a_n1626_n2688# 0.078732f
C187 plus.n26 a_n1626_n2688# 0.019069f
C188 plus.n27 a_n1626_n2688# 0.078732f
C189 plus.n28 a_n1626_n2688# 0.095949f
C190 plus.n29 a_n1626_n2688# 1.19934f
.ends

