* NGSPICE file created from diffpair592.ext - technology: sky130A

.subckt diffpair592 minus drain_right drain_left source plus
X0 drain_left.t5 plus.t0 source.t9 a_n1220_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X1 drain_left.t4 plus.t1 source.t8 a_n1220_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X2 drain_right.t5 minus.t0 source.t4 a_n1220_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X3 a_n1220_n4888# a_n1220_n4888# a_n1220_n4888# a_n1220_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.3
X4 drain_right.t4 minus.t1 source.t5 a_n1220_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X5 drain_right.t3 minus.t2 source.t3 a_n1220_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X6 drain_left.t3 plus.t2 source.t11 a_n1220_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X7 a_n1220_n4888# a_n1220_n4888# a_n1220_n4888# a_n1220_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X8 source.t6 plus.t3 drain_left.t2 a_n1220_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X9 drain_right.t2 minus.t3 source.t2 a_n1220_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X10 source.t7 plus.t4 drain_left.t1 a_n1220_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X11 drain_left.t0 plus.t5 source.t10 a_n1220_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X12 a_n1220_n4888# a_n1220_n4888# a_n1220_n4888# a_n1220_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X13 source.t1 minus.t4 drain_right.t1 a_n1220_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X14 source.t0 minus.t5 drain_right.t0 a_n1220_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X15 a_n1220_n4888# a_n1220_n4888# a_n1220_n4888# a_n1220_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
R0 plus.n0 plus.t2 1766.6
R1 plus.n2 plus.t5 1766.6
R2 plus.n4 plus.t0 1766.6
R3 plus.n6 plus.t1 1766.6
R4 plus.n1 plus.t3 1711.1
R5 plus.n5 plus.t4 1711.1
R6 plus.n3 plus.n0 161.489
R7 plus.n7 plus.n4 161.489
R8 plus.n3 plus.n2 161.3
R9 plus.n7 plus.n6 161.3
R10 plus.n1 plus.n0 36.5157
R11 plus.n2 plus.n1 36.5157
R12 plus.n6 plus.n5 36.5157
R13 plus.n5 plus.n4 36.5157
R14 plus plus.n7 30.6865
R15 plus plus.n3 15.2069
R16 source.n0 source.t10 44.1297
R17 source.n3 source.t2 44.1296
R18 source.n11 source.t5 44.1295
R19 source.n8 source.t9 44.1295
R20 source.n2 source.n1 43.1397
R21 source.n5 source.n4 43.1397
R22 source.n10 source.n9 43.1396
R23 source.n7 source.n6 43.1396
R24 source.n7 source.n5 28.4345
R25 source.n12 source.n0 22.357
R26 source.n12 source.n11 5.53498
R27 source.n9 source.t3 0.9905
R28 source.n9 source.t1 0.9905
R29 source.n6 source.t8 0.9905
R30 source.n6 source.t7 0.9905
R31 source.n1 source.t11 0.9905
R32 source.n1 source.t6 0.9905
R33 source.n4 source.t4 0.9905
R34 source.n4 source.t0 0.9905
R35 source.n3 source.n2 0.741879
R36 source.n10 source.n8 0.741879
R37 source.n5 source.n3 0.543603
R38 source.n2 source.n0 0.543603
R39 source.n8 source.n7 0.543603
R40 source.n11 source.n10 0.543603
R41 source source.n12 0.188
R42 drain_left.n3 drain_left.t3 61.3515
R43 drain_left.n1 drain_left.t4 61.1603
R44 drain_left.n1 drain_left.n0 59.8988
R45 drain_left.n3 drain_left.n2 59.8185
R46 drain_left drain_left.n1 34.9212
R47 drain_left drain_left.n3 6.19632
R48 drain_left.n0 drain_left.t1 0.9905
R49 drain_left.n0 drain_left.t5 0.9905
R50 drain_left.n2 drain_left.t2 0.9905
R51 drain_left.n2 drain_left.t0 0.9905
R52 minus.n2 minus.t0 1766.6
R53 minus.n0 minus.t3 1766.6
R54 minus.n6 minus.t1 1766.6
R55 minus.n4 minus.t2 1766.6
R56 minus.n1 minus.t5 1711.1
R57 minus.n5 minus.t4 1711.1
R58 minus.n3 minus.n0 161.489
R59 minus.n7 minus.n4 161.489
R60 minus.n3 minus.n2 161.3
R61 minus.n7 minus.n6 161.3
R62 minus.n8 minus.n3 39.8357
R63 minus.n2 minus.n1 36.5157
R64 minus.n1 minus.n0 36.5157
R65 minus.n5 minus.n4 36.5157
R66 minus.n6 minus.n5 36.5157
R67 minus.n8 minus.n7 6.5327
R68 minus minus.n8 0.188
R69 drain_right.n1 drain_right.t3 61.1603
R70 drain_right.n3 drain_right.t5 60.8084
R71 drain_right.n3 drain_right.n2 60.3616
R72 drain_right.n1 drain_right.n0 59.8988
R73 drain_right drain_right.n1 34.368
R74 drain_right drain_right.n3 5.92477
R75 drain_right.n0 drain_right.t1 0.9905
R76 drain_right.n0 drain_right.t4 0.9905
R77 drain_right.n2 drain_right.t0 0.9905
R78 drain_right.n2 drain_right.t2 0.9905
C0 drain_left source 22.3715f
C1 drain_right plus 0.271207f
C2 minus drain_left 0.17071f
C3 source plus 3.5352f
C4 minus plus 6.14977f
C5 source drain_right 22.353302f
C6 minus drain_right 4.34574f
C7 minus source 3.52007f
C8 drain_left plus 4.4552f
C9 drain_left drain_right 0.572212f
C10 drain_right a_n1220_n4888# 8.672029f
C11 drain_left a_n1220_n4888# 8.871571f
C12 source a_n1220_n4888# 8.919166f
C13 minus a_n1220_n4888# 5.199373f
C14 plus a_n1220_n4888# 7.86072f
C15 drain_right.t3 a_n1220_n4888# 5.13924f
C16 drain_right.t1 a_n1220_n4888# 0.439358f
C17 drain_right.t4 a_n1220_n4888# 0.439358f
C18 drain_right.n0 a_n1220_n4888# 4.01712f
C19 drain_right.n1 a_n1220_n4888# 2.32886f
C20 drain_right.t0 a_n1220_n4888# 0.439358f
C21 drain_right.t2 a_n1220_n4888# 0.439358f
C22 drain_right.n2 a_n1220_n4888# 4.01979f
C23 drain_right.t5 a_n1220_n4888# 5.13721f
C24 drain_right.n3 a_n1220_n4888# 0.944096f
C25 minus.t3 a_n1220_n4888# 0.985149f
C26 minus.n0 a_n1220_n4888# 0.380314f
C27 minus.t0 a_n1220_n4888# 0.985149f
C28 minus.t5 a_n1220_n4888# 0.973585f
C29 minus.n1 a_n1220_n4888# 0.361664f
C30 minus.n2 a_n1220_n4888# 0.380223f
C31 minus.n3 a_n1220_n4888# 2.43709f
C32 minus.t2 a_n1220_n4888# 0.985149f
C33 minus.n4 a_n1220_n4888# 0.380314f
C34 minus.t4 a_n1220_n4888# 0.973585f
C35 minus.n5 a_n1220_n4888# 0.361664f
C36 minus.t1 a_n1220_n4888# 0.985149f
C37 minus.n6 a_n1220_n4888# 0.380223f
C38 minus.n7 a_n1220_n4888# 0.458499f
C39 minus.n8 a_n1220_n4888# 2.83441f
C40 drain_left.t4 a_n1220_n4888# 5.15673f
C41 drain_left.t1 a_n1220_n4888# 0.440853f
C42 drain_left.t5 a_n1220_n4888# 0.440853f
C43 drain_left.n0 a_n1220_n4888# 4.03079f
C44 drain_left.n1 a_n1220_n4888# 2.39543f
C45 drain_left.t3 a_n1220_n4888# 5.158f
C46 drain_left.t2 a_n1220_n4888# 0.440853f
C47 drain_left.t0 a_n1220_n4888# 0.440853f
C48 drain_left.n2 a_n1220_n4888# 4.03037f
C49 drain_left.n3 a_n1220_n4888# 0.93534f
C50 source.t10 a_n1220_n4888# 5.04151f
C51 source.n0 a_n1220_n4888# 2.14432f
C52 source.t11 a_n1220_n4888# 0.441139f
C53 source.t6 a_n1220_n4888# 0.441139f
C54 source.n1 a_n1220_n4888# 3.94397f
C55 source.n2 a_n1220_n4888# 0.402143f
C56 source.t2 a_n1220_n4888# 5.04152f
C57 source.n3 a_n1220_n4888# 0.507706f
C58 source.t4 a_n1220_n4888# 0.441139f
C59 source.t0 a_n1220_n4888# 0.441139f
C60 source.n4 a_n1220_n4888# 3.94397f
C61 source.n5 a_n1220_n4888# 2.58224f
C62 source.t8 a_n1220_n4888# 0.441139f
C63 source.t7 a_n1220_n4888# 0.441139f
C64 source.n6 a_n1220_n4888# 3.94398f
C65 source.n7 a_n1220_n4888# 2.58223f
C66 source.t9 a_n1220_n4888# 5.04149f
C67 source.n8 a_n1220_n4888# 0.507734f
C68 source.t3 a_n1220_n4888# 0.441139f
C69 source.t1 a_n1220_n4888# 0.441139f
C70 source.n9 a_n1220_n4888# 3.94398f
C71 source.n10 a_n1220_n4888# 0.402136f
C72 source.t5 a_n1220_n4888# 5.04149f
C73 source.n11 a_n1220_n4888# 0.640874f
C74 source.n12 a_n1220_n4888# 2.51261f
C75 plus.t2 a_n1220_n4888# 1.00777f
C76 plus.n0 a_n1220_n4888# 0.389047f
C77 plus.t3 a_n1220_n4888# 0.995942f
C78 plus.n1 a_n1220_n4888# 0.369968f
C79 plus.t5 a_n1220_n4888# 1.00777f
C80 plus.n2 a_n1220_n4888# 0.388954f
C81 plus.n3 a_n1220_n4888# 0.978514f
C82 plus.t0 a_n1220_n4888# 1.00777f
C83 plus.n4 a_n1220_n4888# 0.389047f
C84 plus.t1 a_n1220_n4888# 1.00777f
C85 plus.t4 a_n1220_n4888# 0.995942f
C86 plus.n5 a_n1220_n4888# 0.369968f
C87 plus.n6 a_n1220_n4888# 0.388954f
C88 plus.n7 a_n1220_n4888# 1.97277f
.ends

