* NGSPICE file created from diffpair201.ext - technology: sky130A

.subckt diffpair201 minus drain_right drain_left source plus
X0 source minus drain_right a_n1214_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X1 source plus drain_left a_n1214_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X2 source minus drain_right a_n1214_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X3 drain_left plus source a_n1214_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X4 drain_right minus source a_n1214_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X5 a_n1214_n1488# a_n1214_n1488# a_n1214_n1488# a_n1214_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.5
X6 source plus drain_left a_n1214_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X7 a_n1214_n1488# a_n1214_n1488# a_n1214_n1488# a_n1214_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X8 a_n1214_n1488# a_n1214_n1488# a_n1214_n1488# a_n1214_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X9 drain_right minus source a_n1214_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X10 drain_left plus source a_n1214_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X11 a_n1214_n1488# a_n1214_n1488# a_n1214_n1488# a_n1214_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
.ends

