* NGSPICE file created from diffpair626.ext - technology: sky130A

.subckt diffpair626 minus drain_right drain_left source plus
X0 drain_left.t13 plus.t0 source.t23 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X1 a_n2364_n4888# a_n2364_n4888# a_n2364_n4888# a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.7
X2 drain_right.t13 minus.t0 source.t8 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X3 source.t13 plus.t1 drain_left.t12 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X4 drain_left.t11 plus.t2 source.t25 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X5 source.t0 minus.t1 drain_right.t12 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X6 drain_left.t10 plus.t3 source.t19 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X7 source.t1 minus.t2 drain_right.t11 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X8 drain_right.t10 minus.t3 source.t2 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X9 drain_left.t9 plus.t4 source.t26 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X10 drain_left.t8 plus.t5 source.t17 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X11 source.t20 plus.t6 drain_left.t7 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X12 drain_left.t6 plus.t7 source.t16 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X13 source.t7 minus.t4 drain_right.t9 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X14 drain_right.t8 minus.t5 source.t10 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X15 a_n2364_n4888# a_n2364_n4888# a_n2364_n4888# a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X16 drain_right.t7 minus.t6 source.t27 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X17 drain_right.t6 minus.t7 source.t6 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X18 drain_right.t5 minus.t8 source.t5 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X19 source.t22 plus.t8 drain_left.t5 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X20 source.t14 plus.t9 drain_left.t4 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X21 source.t24 plus.t10 drain_left.t3 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X22 drain_left.t2 plus.t11 source.t15 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X23 drain_right.t4 minus.t9 source.t12 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X24 a_n2364_n4888# a_n2364_n4888# a_n2364_n4888# a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X25 source.t18 plus.t12 drain_left.t1 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X26 a_n2364_n4888# a_n2364_n4888# a_n2364_n4888# a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X27 drain_left.t0 plus.t13 source.t21 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X28 source.t3 minus.t10 drain_right.t3 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X29 source.t9 minus.t11 drain_right.t2 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X30 source.t11 minus.t12 drain_right.t1 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X31 drain_right.t0 minus.t13 source.t4 a_n2364_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
R0 plus.n5 plus.t5 768.537
R1 plus.n27 plus.t0 768.537
R2 plus.n20 plus.t2 744.691
R3 plus.n18 plus.t9 744.691
R4 plus.n2 plus.t4 744.691
R5 plus.n12 plus.t8 744.691
R6 plus.n4 plus.t3 744.691
R7 plus.n6 plus.t12 744.691
R8 plus.n42 plus.t7 744.691
R9 plus.n40 plus.t6 744.691
R10 plus.n24 plus.t11 744.691
R11 plus.n34 plus.t10 744.691
R12 plus.n26 plus.t13 744.691
R13 plus.n28 plus.t1 744.691
R14 plus.n8 plus.n7 161.3
R15 plus.n9 plus.n4 161.3
R16 plus.n11 plus.n10 161.3
R17 plus.n12 plus.n3 161.3
R18 plus.n14 plus.n13 161.3
R19 plus.n15 plus.n2 161.3
R20 plus.n17 plus.n16 161.3
R21 plus.n18 plus.n1 161.3
R22 plus.n19 plus.n0 161.3
R23 plus.n21 plus.n20 161.3
R24 plus.n30 plus.n29 161.3
R25 plus.n31 plus.n26 161.3
R26 plus.n33 plus.n32 161.3
R27 plus.n34 plus.n25 161.3
R28 plus.n36 plus.n35 161.3
R29 plus.n37 plus.n24 161.3
R30 plus.n39 plus.n38 161.3
R31 plus.n40 plus.n23 161.3
R32 plus.n41 plus.n22 161.3
R33 plus.n43 plus.n42 161.3
R34 plus.n30 plus.n27 44.9119
R35 plus.n8 plus.n5 44.9119
R36 plus plus.n43 35.1373
R37 plus.n20 plus.n19 35.055
R38 plus.n42 plus.n41 35.055
R39 plus.n18 plus.n17 30.6732
R40 plus.n7 plus.n6 30.6732
R41 plus.n40 plus.n39 30.6732
R42 plus.n29 plus.n28 30.6732
R43 plus.n13 plus.n2 26.2914
R44 plus.n11 plus.n4 26.2914
R45 plus.n35 plus.n24 26.2914
R46 plus.n33 plus.n26 26.2914
R47 plus.n13 plus.n12 21.9096
R48 plus.n12 plus.n11 21.9096
R49 plus.n35 plus.n34 21.9096
R50 plus.n34 plus.n33 21.9096
R51 plus.n28 plus.n27 17.739
R52 plus.n6 plus.n5 17.739
R53 plus.n17 plus.n2 17.5278
R54 plus.n7 plus.n4 17.5278
R55 plus.n39 plus.n24 17.5278
R56 plus.n29 plus.n26 17.5278
R57 plus plus.n21 15.3244
R58 plus.n19 plus.n18 13.146
R59 plus.n41 plus.n40 13.146
R60 plus.n9 plus.n8 0.189894
R61 plus.n10 plus.n9 0.189894
R62 plus.n10 plus.n3 0.189894
R63 plus.n14 plus.n3 0.189894
R64 plus.n15 plus.n14 0.189894
R65 plus.n16 plus.n15 0.189894
R66 plus.n16 plus.n1 0.189894
R67 plus.n1 plus.n0 0.189894
R68 plus.n21 plus.n0 0.189894
R69 plus.n43 plus.n22 0.189894
R70 plus.n23 plus.n22 0.189894
R71 plus.n38 plus.n23 0.189894
R72 plus.n38 plus.n37 0.189894
R73 plus.n37 plus.n36 0.189894
R74 plus.n36 plus.n25 0.189894
R75 plus.n32 plus.n25 0.189894
R76 plus.n32 plus.n31 0.189894
R77 plus.n31 plus.n30 0.189894
R78 source.n0 source.t25 44.1297
R79 source.n7 source.t12 44.1296
R80 source.n27 source.t4 44.1295
R81 source.n20 source.t23 44.1295
R82 source.n2 source.n1 43.1397
R83 source.n4 source.n3 43.1397
R84 source.n6 source.n5 43.1397
R85 source.n9 source.n8 43.1397
R86 source.n11 source.n10 43.1397
R87 source.n13 source.n12 43.1397
R88 source.n26 source.n25 43.1396
R89 source.n24 source.n23 43.1396
R90 source.n22 source.n21 43.1396
R91 source.n19 source.n18 43.1396
R92 source.n17 source.n16 43.1396
R93 source.n15 source.n14 43.1396
R94 source.n15 source.n13 29.1242
R95 source.n28 source.n0 22.5294
R96 source.n28 source.n27 5.7074
R97 source.n25 source.t2 0.9905
R98 source.n25 source.t3 0.9905
R99 source.n23 source.t8 0.9905
R100 source.n23 source.t0 0.9905
R101 source.n21 source.t10 0.9905
R102 source.n21 source.t7 0.9905
R103 source.n18 source.t21 0.9905
R104 source.n18 source.t13 0.9905
R105 source.n16 source.t15 0.9905
R106 source.n16 source.t24 0.9905
R107 source.n14 source.t16 0.9905
R108 source.n14 source.t20 0.9905
R109 source.n1 source.t26 0.9905
R110 source.n1 source.t14 0.9905
R111 source.n3 source.t19 0.9905
R112 source.n3 source.t22 0.9905
R113 source.n5 source.t17 0.9905
R114 source.n5 source.t18 0.9905
R115 source.n8 source.t5 0.9905
R116 source.n8 source.t1 0.9905
R117 source.n10 source.t6 0.9905
R118 source.n10 source.t9 0.9905
R119 source.n12 source.t27 0.9905
R120 source.n12 source.t11 0.9905
R121 source.n7 source.n6 0.914293
R122 source.n22 source.n20 0.914293
R123 source.n13 source.n11 0.888431
R124 source.n11 source.n9 0.888431
R125 source.n9 source.n7 0.888431
R126 source.n6 source.n4 0.888431
R127 source.n4 source.n2 0.888431
R128 source.n2 source.n0 0.888431
R129 source.n17 source.n15 0.888431
R130 source.n19 source.n17 0.888431
R131 source.n20 source.n19 0.888431
R132 source.n24 source.n22 0.888431
R133 source.n26 source.n24 0.888431
R134 source.n27 source.n26 0.888431
R135 source source.n28 0.188
R136 drain_left.n7 drain_left.t8 61.6963
R137 drain_left.n1 drain_left.t6 61.6962
R138 drain_left.n4 drain_left.n2 60.7063
R139 drain_left.n11 drain_left.n10 59.8185
R140 drain_left.n9 drain_left.n8 59.8185
R141 drain_left.n7 drain_left.n6 59.8185
R142 drain_left.n4 drain_left.n3 59.8184
R143 drain_left.n1 drain_left.n0 59.8184
R144 drain_left drain_left.n5 38.5333
R145 drain_left drain_left.n11 6.54115
R146 drain_left.n2 drain_left.t12 0.9905
R147 drain_left.n2 drain_left.t13 0.9905
R148 drain_left.n3 drain_left.t3 0.9905
R149 drain_left.n3 drain_left.t0 0.9905
R150 drain_left.n0 drain_left.t7 0.9905
R151 drain_left.n0 drain_left.t2 0.9905
R152 drain_left.n10 drain_left.t4 0.9905
R153 drain_left.n10 drain_left.t11 0.9905
R154 drain_left.n8 drain_left.t5 0.9905
R155 drain_left.n8 drain_left.t9 0.9905
R156 drain_left.n6 drain_left.t1 0.9905
R157 drain_left.n6 drain_left.t10 0.9905
R158 drain_left.n9 drain_left.n7 0.888431
R159 drain_left.n11 drain_left.n9 0.888431
R160 drain_left.n5 drain_left.n1 0.611102
R161 drain_left.n5 drain_left.n4 0.167137
R162 minus.n5 minus.t9 768.537
R163 minus.n27 minus.t5 768.537
R164 minus.n6 minus.t2 744.691
R165 minus.n8 minus.t8 744.691
R166 minus.n12 minus.t11 744.691
R167 minus.n14 minus.t7 744.691
R168 minus.n18 minus.t12 744.691
R169 minus.n20 minus.t6 744.691
R170 minus.n28 minus.t4 744.691
R171 minus.n30 minus.t0 744.691
R172 minus.n34 minus.t1 744.691
R173 minus.n36 minus.t3 744.691
R174 minus.n40 minus.t10 744.691
R175 minus.n42 minus.t13 744.691
R176 minus.n21 minus.n20 161.3
R177 minus.n19 minus.n0 161.3
R178 minus.n18 minus.n17 161.3
R179 minus.n16 minus.n1 161.3
R180 minus.n15 minus.n14 161.3
R181 minus.n13 minus.n2 161.3
R182 minus.n12 minus.n11 161.3
R183 minus.n10 minus.n3 161.3
R184 minus.n9 minus.n8 161.3
R185 minus.n7 minus.n4 161.3
R186 minus.n43 minus.n42 161.3
R187 minus.n41 minus.n22 161.3
R188 minus.n40 minus.n39 161.3
R189 minus.n38 minus.n23 161.3
R190 minus.n37 minus.n36 161.3
R191 minus.n35 minus.n24 161.3
R192 minus.n34 minus.n33 161.3
R193 minus.n32 minus.n25 161.3
R194 minus.n31 minus.n30 161.3
R195 minus.n29 minus.n26 161.3
R196 minus.n5 minus.n4 44.9119
R197 minus.n27 minus.n26 44.9119
R198 minus.n44 minus.n21 44.2865
R199 minus.n20 minus.n19 35.055
R200 minus.n42 minus.n41 35.055
R201 minus.n7 minus.n6 30.6732
R202 minus.n18 minus.n1 30.6732
R203 minus.n29 minus.n28 30.6732
R204 minus.n40 minus.n23 30.6732
R205 minus.n8 minus.n3 26.2914
R206 minus.n14 minus.n13 26.2914
R207 minus.n30 minus.n25 26.2914
R208 minus.n36 minus.n35 26.2914
R209 minus.n12 minus.n3 21.9096
R210 minus.n13 minus.n12 21.9096
R211 minus.n34 minus.n25 21.9096
R212 minus.n35 minus.n34 21.9096
R213 minus.n6 minus.n5 17.739
R214 minus.n28 minus.n27 17.739
R215 minus.n8 minus.n7 17.5278
R216 minus.n14 minus.n1 17.5278
R217 minus.n30 minus.n29 17.5278
R218 minus.n36 minus.n23 17.5278
R219 minus.n19 minus.n18 13.146
R220 minus.n41 minus.n40 13.146
R221 minus.n44 minus.n43 6.65012
R222 minus.n21 minus.n0 0.189894
R223 minus.n17 minus.n0 0.189894
R224 minus.n17 minus.n16 0.189894
R225 minus.n16 minus.n15 0.189894
R226 minus.n15 minus.n2 0.189894
R227 minus.n11 minus.n2 0.189894
R228 minus.n11 minus.n10 0.189894
R229 minus.n10 minus.n9 0.189894
R230 minus.n9 minus.n4 0.189894
R231 minus.n31 minus.n26 0.189894
R232 minus.n32 minus.n31 0.189894
R233 minus.n33 minus.n32 0.189894
R234 minus.n33 minus.n24 0.189894
R235 minus.n37 minus.n24 0.189894
R236 minus.n38 minus.n37 0.189894
R237 minus.n39 minus.n38 0.189894
R238 minus.n39 minus.n22 0.189894
R239 minus.n43 minus.n22 0.189894
R240 minus minus.n44 0.188
R241 drain_right.n1 drain_right.t8 61.6962
R242 drain_right.n11 drain_right.t7 60.8084
R243 drain_right.n8 drain_right.n6 60.7064
R244 drain_right.n4 drain_right.n2 60.7063
R245 drain_right.n8 drain_right.n7 59.8185
R246 drain_right.n10 drain_right.n9 59.8185
R247 drain_right.n4 drain_right.n3 59.8184
R248 drain_right.n1 drain_right.n0 59.8184
R249 drain_right drain_right.n5 37.9801
R250 drain_right drain_right.n11 6.09718
R251 drain_right.n2 drain_right.t3 0.9905
R252 drain_right.n2 drain_right.t0 0.9905
R253 drain_right.n3 drain_right.t12 0.9905
R254 drain_right.n3 drain_right.t10 0.9905
R255 drain_right.n0 drain_right.t9 0.9905
R256 drain_right.n0 drain_right.t13 0.9905
R257 drain_right.n6 drain_right.t11 0.9905
R258 drain_right.n6 drain_right.t4 0.9905
R259 drain_right.n7 drain_right.t2 0.9905
R260 drain_right.n7 drain_right.t5 0.9905
R261 drain_right.n9 drain_right.t1 0.9905
R262 drain_right.n9 drain_right.t6 0.9905
R263 drain_right.n11 drain_right.n10 0.888431
R264 drain_right.n10 drain_right.n8 0.888431
R265 drain_right.n5 drain_right.n1 0.611102
R266 drain_right.n5 drain_right.n4 0.167137
C0 minus source 14.398499f
C1 drain_left drain_right 1.23643f
C2 plus source 14.413401f
C3 plus minus 7.57396f
C4 drain_right source 28.9182f
C5 drain_right minus 14.750099f
C6 drain_left source 28.9296f
C7 drain_left minus 0.172675f
C8 plus drain_right 0.392237f
C9 plus drain_left 14.9794f
C10 drain_right a_n2364_n4888# 9.75187f
C11 drain_left a_n2364_n4888# 10.0999f
C12 source a_n2364_n4888# 9.577408f
C13 minus a_n2364_n4888# 9.92189f
C14 plus a_n2364_n4888# 12.05124f
C15 drain_right.t8 a_n2364_n4888# 4.6131f
C16 drain_right.t9 a_n2364_n4888# 0.39409f
C17 drain_right.t13 a_n2364_n4888# 0.39409f
C18 drain_right.n0 a_n2364_n4888# 3.60286f
C19 drain_right.n1 a_n2364_n4888# 0.68812f
C20 drain_right.t3 a_n2364_n4888# 0.39409f
C21 drain_right.t0 a_n2364_n4888# 0.39409f
C22 drain_right.n2 a_n2364_n4888# 3.60817f
C23 drain_right.t12 a_n2364_n4888# 0.39409f
C24 drain_right.t10 a_n2364_n4888# 0.39409f
C25 drain_right.n3 a_n2364_n4888# 3.60286f
C26 drain_right.n4 a_n2364_n4888# 0.65645f
C27 drain_right.n5 a_n2364_n4888# 1.81553f
C28 drain_right.t11 a_n2364_n4888# 0.39409f
C29 drain_right.t4 a_n2364_n4888# 0.39409f
C30 drain_right.n6 a_n2364_n4888# 3.60817f
C31 drain_right.t2 a_n2364_n4888# 0.39409f
C32 drain_right.t5 a_n2364_n4888# 0.39409f
C33 drain_right.n7 a_n2364_n4888# 3.60285f
C34 drain_right.n8 a_n2364_n4888# 0.710945f
C35 drain_right.t1 a_n2364_n4888# 0.39409f
C36 drain_right.t6 a_n2364_n4888# 0.39409f
C37 drain_right.n9 a_n2364_n4888# 3.60285f
C38 drain_right.n10 a_n2364_n4888# 0.353106f
C39 drain_right.t7 a_n2364_n4888# 4.60791f
C40 drain_right.n11 a_n2364_n4888# 0.590708f
C41 minus.n0 a_n2364_n4888# 0.040827f
C42 minus.n1 a_n2364_n4888# 0.009264f
C43 minus.t12 a_n2364_n4888# 1.61864f
C44 minus.n2 a_n2364_n4888# 0.040827f
C45 minus.n3 a_n2364_n4888# 0.009264f
C46 minus.t11 a_n2364_n4888# 1.61864f
C47 minus.n4 a_n2364_n4888# 0.172021f
C48 minus.t9 a_n2364_n4888# 1.63737f
C49 minus.n5 a_n2364_n4888# 0.588404f
C50 minus.t2 a_n2364_n4888# 1.61864f
C51 minus.n6 a_n2364_n4888# 0.608642f
C52 minus.n7 a_n2364_n4888# 0.009264f
C53 minus.t8 a_n2364_n4888# 1.61864f
C54 minus.n8 a_n2364_n4888# 0.603585f
C55 minus.n9 a_n2364_n4888# 0.040827f
C56 minus.n10 a_n2364_n4888# 0.040827f
C57 minus.n11 a_n2364_n4888# 0.040827f
C58 minus.n12 a_n2364_n4888# 0.603585f
C59 minus.n13 a_n2364_n4888# 0.009264f
C60 minus.t7 a_n2364_n4888# 1.61864f
C61 minus.n14 a_n2364_n4888# 0.603585f
C62 minus.n15 a_n2364_n4888# 0.040827f
C63 minus.n16 a_n2364_n4888# 0.040827f
C64 minus.n17 a_n2364_n4888# 0.040827f
C65 minus.n18 a_n2364_n4888# 0.603585f
C66 minus.n19 a_n2364_n4888# 0.009264f
C67 minus.t6 a_n2364_n4888# 1.61864f
C68 minus.n20 a_n2364_n4888# 0.602075f
C69 minus.n21 a_n2364_n4888# 1.95724f
C70 minus.n22 a_n2364_n4888# 0.040827f
C71 minus.n23 a_n2364_n4888# 0.009264f
C72 minus.n24 a_n2364_n4888# 0.040827f
C73 minus.n25 a_n2364_n4888# 0.009264f
C74 minus.n26 a_n2364_n4888# 0.172021f
C75 minus.t5 a_n2364_n4888# 1.63737f
C76 minus.n27 a_n2364_n4888# 0.588404f
C77 minus.t4 a_n2364_n4888# 1.61864f
C78 minus.n28 a_n2364_n4888# 0.608642f
C79 minus.n29 a_n2364_n4888# 0.009264f
C80 minus.t0 a_n2364_n4888# 1.61864f
C81 minus.n30 a_n2364_n4888# 0.603585f
C82 minus.n31 a_n2364_n4888# 0.040827f
C83 minus.n32 a_n2364_n4888# 0.040827f
C84 minus.n33 a_n2364_n4888# 0.040827f
C85 minus.t1 a_n2364_n4888# 1.61864f
C86 minus.n34 a_n2364_n4888# 0.603585f
C87 minus.n35 a_n2364_n4888# 0.009264f
C88 minus.t3 a_n2364_n4888# 1.61864f
C89 minus.n36 a_n2364_n4888# 0.603585f
C90 minus.n37 a_n2364_n4888# 0.040827f
C91 minus.n38 a_n2364_n4888# 0.040827f
C92 minus.n39 a_n2364_n4888# 0.040827f
C93 minus.t10 a_n2364_n4888# 1.61864f
C94 minus.n40 a_n2364_n4888# 0.603585f
C95 minus.n41 a_n2364_n4888# 0.009264f
C96 minus.t13 a_n2364_n4888# 1.61864f
C97 minus.n42 a_n2364_n4888# 0.602075f
C98 minus.n43 a_n2364_n4888# 0.281253f
C99 minus.n44 a_n2364_n4888# 2.31946f
C100 drain_left.t6 a_n2364_n4888# 4.62389f
C101 drain_left.t7 a_n2364_n4888# 0.395012f
C102 drain_left.t2 a_n2364_n4888# 0.395012f
C103 drain_left.n0 a_n2364_n4888# 3.61129f
C104 drain_left.n1 a_n2364_n4888# 0.68973f
C105 drain_left.t12 a_n2364_n4888# 0.395012f
C106 drain_left.t13 a_n2364_n4888# 0.395012f
C107 drain_left.n2 a_n2364_n4888# 3.61661f
C108 drain_left.t3 a_n2364_n4888# 0.395012f
C109 drain_left.t0 a_n2364_n4888# 0.395012f
C110 drain_left.n3 a_n2364_n4888# 3.61129f
C111 drain_left.n4 a_n2364_n4888# 0.657986f
C112 drain_left.n5 a_n2364_n4888# 1.87142f
C113 drain_left.t8 a_n2364_n4888# 4.62391f
C114 drain_left.t1 a_n2364_n4888# 0.395012f
C115 drain_left.t10 a_n2364_n4888# 0.395012f
C116 drain_left.n6 a_n2364_n4888# 3.61128f
C117 drain_left.n7 a_n2364_n4888# 0.711103f
C118 drain_left.t5 a_n2364_n4888# 0.395012f
C119 drain_left.t9 a_n2364_n4888# 0.395012f
C120 drain_left.n8 a_n2364_n4888# 3.61128f
C121 drain_left.n9 a_n2364_n4888# 0.353933f
C122 drain_left.t4 a_n2364_n4888# 0.395012f
C123 drain_left.t11 a_n2364_n4888# 0.395012f
C124 drain_left.n10 a_n2364_n4888# 3.61128f
C125 drain_left.n11 a_n2364_n4888# 0.575001f
C126 source.t25 a_n2364_n4888# 4.62117f
C127 source.n0 a_n2364_n4888# 2.01034f
C128 source.t26 a_n2364_n4888# 0.40436f
C129 source.t14 a_n2364_n4888# 0.40436f
C130 source.n1 a_n2364_n4888# 3.61515f
C131 source.n2 a_n2364_n4888# 0.409125f
C132 source.t19 a_n2364_n4888# 0.40436f
C133 source.t22 a_n2364_n4888# 0.40436f
C134 source.n3 a_n2364_n4888# 3.61515f
C135 source.n4 a_n2364_n4888# 0.409125f
C136 source.t17 a_n2364_n4888# 0.40436f
C137 source.t18 a_n2364_n4888# 0.40436f
C138 source.n5 a_n2364_n4888# 3.61515f
C139 source.n6 a_n2364_n4888# 0.411257f
C140 source.t12 a_n2364_n4888# 4.62119f
C141 source.n7 a_n2364_n4888# 0.508018f
C142 source.t5 a_n2364_n4888# 0.40436f
C143 source.t1 a_n2364_n4888# 0.40436f
C144 source.n8 a_n2364_n4888# 3.61515f
C145 source.n9 a_n2364_n4888# 0.409125f
C146 source.t6 a_n2364_n4888# 0.40436f
C147 source.t9 a_n2364_n4888# 0.40436f
C148 source.n10 a_n2364_n4888# 3.61515f
C149 source.n11 a_n2364_n4888# 0.409125f
C150 source.t27 a_n2364_n4888# 0.40436f
C151 source.t11 a_n2364_n4888# 0.40436f
C152 source.n12 a_n2364_n4888# 3.61515f
C153 source.n13 a_n2364_n4888# 2.45223f
C154 source.t16 a_n2364_n4888# 0.40436f
C155 source.t20 a_n2364_n4888# 0.40436f
C156 source.n14 a_n2364_n4888# 3.61515f
C157 source.n15 a_n2364_n4888# 2.45222f
C158 source.t15 a_n2364_n4888# 0.40436f
C159 source.t24 a_n2364_n4888# 0.40436f
C160 source.n16 a_n2364_n4888# 3.61515f
C161 source.n17 a_n2364_n4888# 0.409117f
C162 source.t21 a_n2364_n4888# 0.40436f
C163 source.t13 a_n2364_n4888# 0.40436f
C164 source.n18 a_n2364_n4888# 3.61515f
C165 source.n19 a_n2364_n4888# 0.409117f
C166 source.t23 a_n2364_n4888# 4.62116f
C167 source.n20 a_n2364_n4888# 0.508044f
C168 source.t10 a_n2364_n4888# 0.40436f
C169 source.t7 a_n2364_n4888# 0.40436f
C170 source.n21 a_n2364_n4888# 3.61515f
C171 source.n22 a_n2364_n4888# 0.411249f
C172 source.t8 a_n2364_n4888# 0.40436f
C173 source.t0 a_n2364_n4888# 0.40436f
C174 source.n23 a_n2364_n4888# 3.61515f
C175 source.n24 a_n2364_n4888# 0.409117f
C176 source.t2 a_n2364_n4888# 0.40436f
C177 source.t3 a_n2364_n4888# 0.40436f
C178 source.n25 a_n2364_n4888# 3.61515f
C179 source.n26 a_n2364_n4888# 0.409117f
C180 source.t4 a_n2364_n4888# 4.62116f
C181 source.n27 a_n2364_n4888# 0.638335f
C182 source.n28 a_n2364_n4888# 2.32114f
C183 plus.n0 a_n2364_n4888# 0.041141f
C184 plus.t2 a_n2364_n4888# 1.63109f
C185 plus.t9 a_n2364_n4888# 1.63109f
C186 plus.n1 a_n2364_n4888# 0.041141f
C187 plus.t4 a_n2364_n4888# 1.63109f
C188 plus.n2 a_n2364_n4888# 0.60823f
C189 plus.n3 a_n2364_n4888# 0.041141f
C190 plus.t8 a_n2364_n4888# 1.63109f
C191 plus.t3 a_n2364_n4888# 1.63109f
C192 plus.n4 a_n2364_n4888# 0.60823f
C193 plus.t5 a_n2364_n4888# 1.64997f
C194 plus.n5 a_n2364_n4888# 0.592932f
C195 plus.t12 a_n2364_n4888# 1.63109f
C196 plus.n6 a_n2364_n4888# 0.613326f
C197 plus.n7 a_n2364_n4888# 0.009336f
C198 plus.n8 a_n2364_n4888# 0.173345f
C199 plus.n9 a_n2364_n4888# 0.041141f
C200 plus.n10 a_n2364_n4888# 0.041141f
C201 plus.n11 a_n2364_n4888# 0.009336f
C202 plus.n12 a_n2364_n4888# 0.60823f
C203 plus.n13 a_n2364_n4888# 0.009336f
C204 plus.n14 a_n2364_n4888# 0.041141f
C205 plus.n15 a_n2364_n4888# 0.041141f
C206 plus.n16 a_n2364_n4888# 0.041141f
C207 plus.n17 a_n2364_n4888# 0.009336f
C208 plus.n18 a_n2364_n4888# 0.60823f
C209 plus.n19 a_n2364_n4888# 0.009336f
C210 plus.n20 a_n2364_n4888# 0.606708f
C211 plus.n21 a_n2364_n4888# 0.638863f
C212 plus.n22 a_n2364_n4888# 0.041141f
C213 plus.t7 a_n2364_n4888# 1.63109f
C214 plus.n23 a_n2364_n4888# 0.041141f
C215 plus.t6 a_n2364_n4888# 1.63109f
C216 plus.t11 a_n2364_n4888# 1.63109f
C217 plus.n24 a_n2364_n4888# 0.60823f
C218 plus.n25 a_n2364_n4888# 0.041141f
C219 plus.t10 a_n2364_n4888# 1.63109f
C220 plus.t13 a_n2364_n4888# 1.63109f
C221 plus.n26 a_n2364_n4888# 0.60823f
C222 plus.t0 a_n2364_n4888# 1.64997f
C223 plus.n27 a_n2364_n4888# 0.592932f
C224 plus.t1 a_n2364_n4888# 1.63109f
C225 plus.n28 a_n2364_n4888# 0.613326f
C226 plus.n29 a_n2364_n4888# 0.009336f
C227 plus.n30 a_n2364_n4888# 0.173345f
C228 plus.n31 a_n2364_n4888# 0.041141f
C229 plus.n32 a_n2364_n4888# 0.041141f
C230 plus.n33 a_n2364_n4888# 0.009336f
C231 plus.n34 a_n2364_n4888# 0.60823f
C232 plus.n35 a_n2364_n4888# 0.009336f
C233 plus.n36 a_n2364_n4888# 0.041141f
C234 plus.n37 a_n2364_n4888# 0.041141f
C235 plus.n38 a_n2364_n4888# 0.041141f
C236 plus.n39 a_n2364_n4888# 0.009336f
C237 plus.n40 a_n2364_n4888# 0.60823f
C238 plus.n41 a_n2364_n4888# 0.009336f
C239 plus.n42 a_n2364_n4888# 0.606708f
C240 plus.n43 a_n2364_n4888# 1.5747f
.ends

