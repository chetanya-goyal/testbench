* NGSPICE file created from diffpair202.ext - technology: sky130A

.subckt diffpair202 minus drain_right drain_left source plus
X0 drain_right.t5 minus.t0 source.t10 a_n1380_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X1 source.t9 minus.t1 drain_right.t4 a_n1380_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X2 drain_left.t5 plus.t0 source.t5 a_n1380_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X3 drain_left.t4 plus.t1 source.t1 a_n1380_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X4 drain_right.t3 minus.t2 source.t11 a_n1380_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X5 drain_left.t3 plus.t2 source.t3 a_n1380_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X6 drain_right.t2 minus.t3 source.t8 a_n1380_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X7 a_n1380_n1488# a_n1380_n1488# a_n1380_n1488# a_n1380_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.5
X8 source.t7 minus.t4 drain_right.t1 a_n1380_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X9 source.t4 plus.t3 drain_left.t2 a_n1380_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X10 drain_right.t0 minus.t5 source.t6 a_n1380_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X11 source.t0 plus.t4 drain_left.t1 a_n1380_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X12 a_n1380_n1488# a_n1380_n1488# a_n1380_n1488# a_n1380_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X13 a_n1380_n1488# a_n1380_n1488# a_n1380_n1488# a_n1380_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X14 drain_left.t0 plus.t5 source.t2 a_n1380_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X15 a_n1380_n1488# a_n1380_n1488# a_n1380_n1488# a_n1380_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
R0 minus.n0 minus.t5 249.988
R1 minus.n4 minus.t2 249.988
R2 minus.n1 minus.t1 223.167
R3 minus.n2 minus.t3 223.167
R4 minus.n5 minus.t4 223.167
R5 minus.n6 minus.t0 223.167
R6 minus.n3 minus.n2 161.3
R7 minus.n7 minus.n6 161.3
R8 minus.n2 minus.n1 48.2005
R9 minus.n6 minus.n5 48.2005
R10 minus.n3 minus.n0 45.1367
R11 minus.n7 minus.n4 45.1367
R12 minus.n8 minus.n3 27.563
R13 minus.n1 minus.n0 13.3799
R14 minus.n5 minus.n4 13.3799
R15 minus.n8 minus.n7 6.5327
R16 minus minus.n8 0.188
R17 source.n0 source.t2 69.6943
R18 source.n3 source.t6 69.6943
R19 source.n11 source.t10 69.6942
R20 source.n8 source.t3 69.6942
R21 source.n2 source.n1 63.0943
R22 source.n5 source.n4 63.0943
R23 source.n10 source.n9 63.0942
R24 source.n7 source.n6 63.0942
R25 source.n7 source.n5 15.9006
R26 source.n12 source.n0 9.56437
R27 source.n9 source.t11 6.6005
R28 source.n9 source.t7 6.6005
R29 source.n6 source.t5 6.6005
R30 source.n6 source.t4 6.6005
R31 source.n1 source.t1 6.6005
R32 source.n1 source.t0 6.6005
R33 source.n4 source.t8 6.6005
R34 source.n4 source.t9 6.6005
R35 source.n12 source.n11 5.62119
R36 source.n3 source.n2 0.828086
R37 source.n10 source.n8 0.828086
R38 source.n5 source.n3 0.716017
R39 source.n2 source.n0 0.716017
R40 source.n8 source.n7 0.716017
R41 source.n11 source.n10 0.716017
R42 source source.n12 0.188
R43 drain_right.n1 drain_right.t3 86.8543
R44 drain_right.n3 drain_right.t2 86.3731
R45 drain_right.n3 drain_right.n2 80.4886
R46 drain_right.n1 drain_right.n0 79.8965
R47 drain_right drain_right.n1 21.9633
R48 drain_right.n0 drain_right.t1 6.6005
R49 drain_right.n0 drain_right.t5 6.6005
R50 drain_right.n2 drain_right.t4 6.6005
R51 drain_right.n2 drain_right.t0 6.6005
R52 drain_right drain_right.n3 6.01097
R53 plus.n0 plus.t1 249.988
R54 plus.n4 plus.t2 249.988
R55 plus.n2 plus.t5 223.167
R56 plus.n1 plus.t4 223.167
R57 plus.n6 plus.t0 223.167
R58 plus.n5 plus.t3 223.167
R59 plus.n3 plus.n2 161.3
R60 plus.n7 plus.n6 161.3
R61 plus.n2 plus.n1 48.2005
R62 plus.n6 plus.n5 48.2005
R63 plus.n3 plus.n0 45.1367
R64 plus.n7 plus.n4 45.1367
R65 plus plus.n7 24.8532
R66 plus.n1 plus.n0 13.3799
R67 plus.n5 plus.n4 13.3799
R68 plus plus.n3 8.76755
R69 drain_left.n3 drain_left.t4 87.0886
R70 drain_left.n1 drain_left.t5 86.8543
R71 drain_left.n1 drain_left.n0 79.8965
R72 drain_left.n3 drain_left.n2 79.7731
R73 drain_left drain_left.n1 22.5166
R74 drain_left.n0 drain_left.t2 6.6005
R75 drain_left.n0 drain_left.t3 6.6005
R76 drain_left.n2 drain_left.t1 6.6005
R77 drain_left.n2 drain_left.t0 6.6005
R78 drain_left drain_left.n3 6.36873
C0 drain_left plus 1.28677f
C1 drain_left drain_right 0.636022f
C2 drain_left source 4.20351f
C3 drain_right plus 0.290883f
C4 minus drain_left 0.176275f
C5 source plus 1.23607f
C6 minus plus 3.20885f
C7 source drain_right 4.20066f
C8 minus drain_right 1.15673f
C9 minus source 1.22193f
C10 drain_right a_n1380_n1488# 3.38577f
C11 drain_left a_n1380_n1488# 3.55733f
C12 source a_n1380_n1488# 2.798104f
C13 minus a_n1380_n1488# 4.567214f
C14 plus a_n1380_n1488# 5.208106f
C15 drain_left.t5 a_n1380_n1488# 0.409856f
C16 drain_left.t2 a_n1380_n1488# 0.04415f
C17 drain_left.t3 a_n1380_n1488# 0.04415f
C18 drain_left.n0 a_n1380_n1488# 0.31873f
C19 drain_left.n1 a_n1380_n1488# 0.91041f
C20 drain_left.t4 a_n1380_n1488# 0.410545f
C21 drain_left.t1 a_n1380_n1488# 0.04415f
C22 drain_left.t0 a_n1380_n1488# 0.04415f
C23 drain_left.n2 a_n1380_n1488# 0.318407f
C24 drain_left.n3 a_n1380_n1488# 0.622732f
C25 plus.t1 a_n1380_n1488# 0.145524f
C26 plus.n0 a_n1380_n1488# 0.0738f
C27 plus.t5 a_n1380_n1488# 0.136718f
C28 plus.t4 a_n1380_n1488# 0.136718f
C29 plus.n1 a_n1380_n1488# 0.088898f
C30 plus.n2 a_n1380_n1488# 0.082f
C31 plus.n3 a_n1380_n1488# 0.323092f
C32 plus.t2 a_n1380_n1488# 0.145524f
C33 plus.n4 a_n1380_n1488# 0.0738f
C34 plus.t0 a_n1380_n1488# 0.136718f
C35 plus.t3 a_n1380_n1488# 0.136718f
C36 plus.n5 a_n1380_n1488# 0.088898f
C37 plus.n6 a_n1380_n1488# 0.082f
C38 plus.n7 a_n1380_n1488# 0.738773f
C39 drain_right.t3 a_n1380_n1488# 0.417091f
C40 drain_right.t1 a_n1380_n1488# 0.044929f
C41 drain_right.t5 a_n1380_n1488# 0.044929f
C42 drain_right.n0 a_n1380_n1488# 0.324357f
C43 drain_right.n1 a_n1380_n1488# 0.888698f
C44 drain_right.t4 a_n1380_n1488# 0.044929f
C45 drain_right.t0 a_n1380_n1488# 0.044929f
C46 drain_right.n2 a_n1380_n1488# 0.32622f
C47 drain_right.t2 a_n1380_n1488# 0.415871f
C48 drain_right.n3 a_n1380_n1488# 0.644443f
C49 source.t2 a_n1380_n1488# 0.443153f
C50 source.n0 a_n1380_n1488# 0.626606f
C51 source.t1 a_n1380_n1488# 0.053367f
C52 source.t0 a_n1380_n1488# 0.053367f
C53 source.n1 a_n1380_n1488# 0.33838f
C54 source.n2 a_n1380_n1488# 0.308034f
C55 source.t6 a_n1380_n1488# 0.443153f
C56 source.n3 a_n1380_n1488# 0.348808f
C57 source.t8 a_n1380_n1488# 0.053367f
C58 source.t9 a_n1380_n1488# 0.053367f
C59 source.n4 a_n1380_n1488# 0.33838f
C60 source.n5 a_n1380_n1488# 0.875399f
C61 source.t5 a_n1380_n1488# 0.053367f
C62 source.t4 a_n1380_n1488# 0.053367f
C63 source.n6 a_n1380_n1488# 0.338377f
C64 source.n7 a_n1380_n1488# 0.875401f
C65 source.t3 a_n1380_n1488# 0.443151f
C66 source.n8 a_n1380_n1488# 0.34881f
C67 source.t11 a_n1380_n1488# 0.053367f
C68 source.t7 a_n1380_n1488# 0.053367f
C69 source.n9 a_n1380_n1488# 0.338377f
C70 source.n10 a_n1380_n1488# 0.308036f
C71 source.t10 a_n1380_n1488# 0.443151f
C72 source.n11 a_n1380_n1488# 0.459874f
C73 source.n12 a_n1380_n1488# 0.658078f
C74 minus.t5 a_n1380_n1488# 0.142782f
C75 minus.n0 a_n1380_n1488# 0.072409f
C76 minus.t1 a_n1380_n1488# 0.134142f
C77 minus.n1 a_n1380_n1488# 0.087222f
C78 minus.t3 a_n1380_n1488# 0.134142f
C79 minus.n2 a_n1380_n1488# 0.080455f
C80 minus.n3 a_n1380_n1488# 0.76195f
C81 minus.t2 a_n1380_n1488# 0.142782f
C82 minus.n4 a_n1380_n1488# 0.072409f
C83 minus.t4 a_n1380_n1488# 0.134142f
C84 minus.n5 a_n1380_n1488# 0.087222f
C85 minus.t0 a_n1380_n1488# 0.134142f
C86 minus.n6 a_n1380_n1488# 0.080455f
C87 minus.n7 a_n1380_n1488# 0.289083f
C88 minus.n8 a_n1380_n1488# 0.82708f
.ends

