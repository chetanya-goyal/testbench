* NGSPICE file created from diffpair331.ext - technology: sky130A

.subckt diffpair331 minus drain_right drain_left source plus
X0 drain_right minus source a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X1 a_n1034_n2692# a_n1034_n2692# a_n1034_n2692# a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.2
X2 a_n1034_n2692# a_n1034_n2692# a_n1034_n2692# a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X3 drain_left plus source a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X4 a_n1034_n2692# a_n1034_n2692# a_n1034_n2692# a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X5 source plus drain_left a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X6 source minus drain_right a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X7 drain_right minus source a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X8 drain_left plus source a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X9 a_n1034_n2692# a_n1034_n2692# a_n1034_n2692# a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X10 source minus drain_right a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X11 source plus drain_left a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
.ends

