* NGSPICE file created from diffpair324.ext - technology: sky130A

.subckt diffpair324 minus drain_right drain_left source plus
X0 drain_left.t9 plus.t0 source.t18 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X1 source.t9 plus.t1 drain_left.t8 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X2 drain_right.t9 minus.t0 source.t6 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X3 a_n1496_n2688# a_n1496_n2688# a_n1496_n2688# a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=34.2 ps=151.6 w=9 l=0.15
X4 drain_left.t7 plus.t2 source.t14 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X5 a_n1496_n2688# a_n1496_n2688# a_n1496_n2688# a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X6 a_n1496_n2688# a_n1496_n2688# a_n1496_n2688# a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X7 source.t0 minus.t1 drain_right.t8 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X8 drain_left.t6 plus.t3 source.t12 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X9 source.t1 minus.t2 drain_right.t7 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X10 source.t15 plus.t4 drain_left.t5 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X11 drain_right.t6 minus.t3 source.t2 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
X12 drain_right.t5 minus.t4 source.t5 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X13 drain_right.t4 minus.t5 source.t7 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X14 source.t19 minus.t6 drain_right.t3 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X15 a_n1496_n2688# a_n1496_n2688# a_n1496_n2688# a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=0 ps=0 w=9 l=0.15
X16 drain_left.t4 plus.t5 source.t16 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X17 drain_right.t2 minus.t7 source.t4 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X18 source.t10 plus.t6 drain_left.t3 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X19 source.t3 minus.t8 drain_right.t1 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X20 drain_left.t2 plus.t7 source.t11 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X21 source.t13 plus.t8 drain_left.t1 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=2.25 ps=9.5 w=9 l=0.15
X22 drain_right.t0 minus.t9 source.t8 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=4.275 pd=18.95 as=2.25 ps=9.5 w=9 l=0.15
X23 drain_left.t0 plus.t9 source.t17 a_n1496_n2688# sky130_fd_pr__nfet_01v8 ad=2.25 pd=9.5 as=4.275 ps=18.95 w=9 l=0.15
R0 plus.n3 plus.t5 1698.68
R1 plus.n9 plus.t9 1698.68
R2 plus.n14 plus.t2 1698.68
R3 plus.n20 plus.t3 1698.68
R4 plus.n6 plus.t7 1654.87
R5 plus.n2 plus.t8 1654.87
R6 plus.n8 plus.t6 1654.87
R7 plus.n17 plus.t0 1654.87
R8 plus.n13 plus.t4 1654.87
R9 plus.n19 plus.t1 1654.87
R10 plus.n4 plus.n3 161.489
R11 plus.n15 plus.n14 161.489
R12 plus.n4 plus.n1 161.3
R13 plus.n6 plus.n5 161.3
R14 plus.n7 plus.n0 161.3
R15 plus.n10 plus.n9 161.3
R16 plus.n15 plus.n12 161.3
R17 plus.n17 plus.n16 161.3
R18 plus.n18 plus.n11 161.3
R19 plus.n21 plus.n20 161.3
R20 plus.n6 plus.n1 73.0308
R21 plus.n7 plus.n6 73.0308
R22 plus.n18 plus.n17 73.0308
R23 plus.n17 plus.n12 73.0308
R24 plus.n3 plus.n2 51.1217
R25 plus.n9 plus.n8 51.1217
R26 plus.n20 plus.n19 51.1217
R27 plus.n14 plus.n13 51.1217
R28 plus plus.n21 27.5464
R29 plus.n2 plus.n1 21.9096
R30 plus.n8 plus.n7 21.9096
R31 plus.n19 plus.n18 21.9096
R32 plus.n13 plus.n12 21.9096
R33 plus plus.n10 11.0213
R34 plus.n5 plus.n4 0.189894
R35 plus.n5 plus.n0 0.189894
R36 plus.n10 plus.n0 0.189894
R37 plus.n21 plus.n11 0.189894
R38 plus.n16 plus.n11 0.189894
R39 plus.n16 plus.n15 0.189894
R40 source.n5 source.t2 52.1921
R41 source.n19 source.t6 52.1919
R42 source.n14 source.t14 52.1919
R43 source.n0 source.t17 52.1919
R44 source.n2 source.n1 48.8588
R45 source.n4 source.n3 48.8588
R46 source.n7 source.n6 48.8588
R47 source.n9 source.n8 48.8588
R48 source.n18 source.n17 48.8586
R49 source.n16 source.n15 48.8586
R50 source.n13 source.n12 48.8586
R51 source.n11 source.n10 48.8586
R52 source.n11 source.n9 20.1357
R53 source.n20 source.n0 14.0322
R54 source.n20 source.n19 5.5436
R55 source.n17 source.t7 3.33383
R56 source.n17 source.t3 3.33383
R57 source.n15 source.t8 3.33383
R58 source.n15 source.t0 3.33383
R59 source.n12 source.t18 3.33383
R60 source.n12 source.t15 3.33383
R61 source.n10 source.t12 3.33383
R62 source.n10 source.t9 3.33383
R63 source.n1 source.t11 3.33383
R64 source.n1 source.t10 3.33383
R65 source.n3 source.t16 3.33383
R66 source.n3 source.t13 3.33383
R67 source.n6 source.t4 3.33383
R68 source.n6 source.t1 3.33383
R69 source.n8 source.t5 3.33383
R70 source.n8 source.t19 3.33383
R71 source.n5 source.n4 0.7505
R72 source.n16 source.n14 0.7505
R73 source.n9 source.n7 0.560845
R74 source.n7 source.n5 0.560845
R75 source.n4 source.n2 0.560845
R76 source.n2 source.n0 0.560845
R77 source.n13 source.n11 0.560845
R78 source.n14 source.n13 0.560845
R79 source.n18 source.n16 0.560845
R80 source.n19 source.n18 0.560845
R81 source source.n20 0.188
R82 drain_left.n5 drain_left.t4 69.4313
R83 drain_left.n1 drain_left.t6 69.431
R84 drain_left.n3 drain_left.n2 65.9022
R85 drain_left.n5 drain_left.n4 65.5376
R86 drain_left.n7 drain_left.n6 65.5374
R87 drain_left.n1 drain_left.n0 65.5373
R88 drain_left drain_left.n3 27.4758
R89 drain_left drain_left.n7 6.21356
R90 drain_left.n2 drain_left.t5 3.33383
R91 drain_left.n2 drain_left.t7 3.33383
R92 drain_left.n0 drain_left.t8 3.33383
R93 drain_left.n0 drain_left.t9 3.33383
R94 drain_left.n6 drain_left.t3 3.33383
R95 drain_left.n6 drain_left.t0 3.33383
R96 drain_left.n4 drain_left.t1 3.33383
R97 drain_left.n4 drain_left.t2 3.33383
R98 drain_left.n7 drain_left.n5 0.560845
R99 drain_left.n3 drain_left.n1 0.0852402
R100 minus.n9 minus.t4 1698.68
R101 minus.n3 minus.t3 1698.68
R102 minus.n20 minus.t0 1698.68
R103 minus.n14 minus.t9 1698.68
R104 minus.n6 minus.t7 1654.87
R105 minus.n8 minus.t6 1654.87
R106 minus.n2 minus.t2 1654.87
R107 minus.n17 minus.t5 1654.87
R108 minus.n19 minus.t8 1654.87
R109 minus.n13 minus.t1 1654.87
R110 minus.n4 minus.n3 161.489
R111 minus.n15 minus.n14 161.489
R112 minus.n10 minus.n9 161.3
R113 minus.n7 minus.n0 161.3
R114 minus.n6 minus.n5 161.3
R115 minus.n4 minus.n1 161.3
R116 minus.n21 minus.n20 161.3
R117 minus.n18 minus.n11 161.3
R118 minus.n17 minus.n16 161.3
R119 minus.n15 minus.n12 161.3
R120 minus.n7 minus.n6 73.0308
R121 minus.n6 minus.n1 73.0308
R122 minus.n17 minus.n12 73.0308
R123 minus.n18 minus.n17 73.0308
R124 minus.n9 minus.n8 51.1217
R125 minus.n3 minus.n2 51.1217
R126 minus.n14 minus.n13 51.1217
R127 minus.n20 minus.n19 51.1217
R128 minus.n22 minus.n10 32.5289
R129 minus.n8 minus.n7 21.9096
R130 minus.n2 minus.n1 21.9096
R131 minus.n13 minus.n12 21.9096
R132 minus.n19 minus.n18 21.9096
R133 minus.n22 minus.n21 6.51376
R134 minus.n10 minus.n0 0.189894
R135 minus.n5 minus.n0 0.189894
R136 minus.n5 minus.n4 0.189894
R137 minus.n16 minus.n15 0.189894
R138 minus.n16 minus.n11 0.189894
R139 minus.n21 minus.n11 0.189894
R140 minus minus.n22 0.188
R141 drain_right.n1 drain_right.t0 69.431
R142 drain_right.n7 drain_right.t5 68.8709
R143 drain_right.n6 drain_right.n4 66.0978
R144 drain_right.n3 drain_right.n2 65.9022
R145 drain_right.n6 drain_right.n5 65.5376
R146 drain_right.n1 drain_right.n0 65.5373
R147 drain_right drain_right.n3 26.9226
R148 drain_right drain_right.n7 5.93339
R149 drain_right.n2 drain_right.t1 3.33383
R150 drain_right.n2 drain_right.t9 3.33383
R151 drain_right.n0 drain_right.t8 3.33383
R152 drain_right.n0 drain_right.t4 3.33383
R153 drain_right.n4 drain_right.t7 3.33383
R154 drain_right.n4 drain_right.t6 3.33383
R155 drain_right.n5 drain_right.t3 3.33383
R156 drain_right.n5 drain_right.t2 3.33383
R157 drain_right.n7 drain_right.n6 0.560845
R158 drain_right.n3 drain_right.n1 0.0852402
C0 plus minus 4.44792f
C1 drain_right plus 0.298099f
C2 source drain_left 16.6504f
C3 minus drain_left 0.170828f
C4 drain_right drain_left 0.735254f
C5 source minus 1.59805f
C6 drain_right source 16.642f
C7 plus drain_left 2.12472f
C8 drain_right minus 1.98386f
C9 source plus 1.61258f
C10 drain_right a_n1496_n2688# 5.47698f
C11 drain_left a_n1496_n2688# 5.94163f
C12 source a_n1496_n2688# 5.104126f
C13 minus a_n1496_n2688# 5.280847f
C14 plus a_n1496_n2688# 6.78543f
C15 drain_right.t0 a_n1496_n2688# 1.92989f
C16 drain_right.t8 a_n1496_n2688# 0.243912f
C17 drain_right.t4 a_n1496_n2688# 0.243912f
C18 drain_right.n0 a_n1496_n2688# 1.57391f
C19 drain_right.n1 a_n1496_n2688# 0.548909f
C20 drain_right.t1 a_n1496_n2688# 0.243912f
C21 drain_right.t9 a_n1496_n2688# 0.243912f
C22 drain_right.n2 a_n1496_n2688# 1.57535f
C23 drain_right.n3 a_n1496_n2688# 1.0831f
C24 drain_right.t7 a_n1496_n2688# 0.243912f
C25 drain_right.t6 a_n1496_n2688# 0.243912f
C26 drain_right.n4 a_n1496_n2688# 1.57622f
C27 drain_right.t3 a_n1496_n2688# 0.243912f
C28 drain_right.t2 a_n1496_n2688# 0.243912f
C29 drain_right.n5 a_n1496_n2688# 1.57391f
C30 drain_right.n6 a_n1496_n2688# 0.532902f
C31 drain_right.t5 a_n1496_n2688# 1.92733f
C32 drain_right.n7 a_n1496_n2688# 0.506714f
C33 minus.n0 a_n1496_n2688# 0.031076f
C34 minus.t4 a_n1496_n2688# 0.120255f
C35 minus.t6 a_n1496_n2688# 0.118875f
C36 minus.t7 a_n1496_n2688# 0.118875f
C37 minus.n1 a_n1496_n2688# 0.013183f
C38 minus.t2 a_n1496_n2688# 0.118875f
C39 minus.n2 a_n1496_n2688# 0.05443f
C40 minus.t3 a_n1496_n2688# 0.120255f
C41 minus.n3 a_n1496_n2688# 0.065318f
C42 minus.n4 a_n1496_n2688# 0.066899f
C43 minus.n5 a_n1496_n2688# 0.031076f
C44 minus.n6 a_n1496_n2688# 0.064739f
C45 minus.n7 a_n1496_n2688# 0.013183f
C46 minus.n8 a_n1496_n2688# 0.05443f
C47 minus.n9 a_n1496_n2688# 0.065276f
C48 minus.n10 a_n1496_n2688# 0.926035f
C49 minus.n11 a_n1496_n2688# 0.031076f
C50 minus.t8 a_n1496_n2688# 0.118875f
C51 minus.t5 a_n1496_n2688# 0.118875f
C52 minus.n12 a_n1496_n2688# 0.013183f
C53 minus.t9 a_n1496_n2688# 0.120255f
C54 minus.t1 a_n1496_n2688# 0.118875f
C55 minus.n13 a_n1496_n2688# 0.05443f
C56 minus.n14 a_n1496_n2688# 0.065318f
C57 minus.n15 a_n1496_n2688# 0.066899f
C58 minus.n16 a_n1496_n2688# 0.031076f
C59 minus.n17 a_n1496_n2688# 0.064739f
C60 minus.n18 a_n1496_n2688# 0.013183f
C61 minus.n19 a_n1496_n2688# 0.05443f
C62 minus.t0 a_n1496_n2688# 0.120255f
C63 minus.n20 a_n1496_n2688# 0.065276f
C64 minus.n21 a_n1496_n2688# 0.204171f
C65 minus.n22 a_n1496_n2688# 1.1359f
C66 drain_left.t6 a_n1496_n2688# 2.17406f
C67 drain_left.t8 a_n1496_n2688# 0.274772f
C68 drain_left.t9 a_n1496_n2688# 0.274772f
C69 drain_left.n0 a_n1496_n2688# 1.77304f
C70 drain_left.n1 a_n1496_n2688# 0.618358f
C71 drain_left.t5 a_n1496_n2688# 0.274772f
C72 drain_left.t7 a_n1496_n2688# 0.274772f
C73 drain_left.n2 a_n1496_n2688# 1.77466f
C74 drain_left.n3 a_n1496_n2688# 1.27296f
C75 drain_left.t4 a_n1496_n2688# 2.17406f
C76 drain_left.t1 a_n1496_n2688# 0.274772f
C77 drain_left.t2 a_n1496_n2688# 0.274772f
C78 drain_left.n4 a_n1496_n2688# 1.77305f
C79 drain_left.n5 a_n1496_n2688# 0.650452f
C80 drain_left.t3 a_n1496_n2688# 0.274772f
C81 drain_left.t0 a_n1496_n2688# 0.274772f
C82 drain_left.n6 a_n1496_n2688# 1.77304f
C83 drain_left.n7 a_n1496_n2688# 0.509272f
C84 source.t17 a_n1496_n2688# 1.95823f
C85 source.n0 a_n1496_n2688# 1.09234f
C86 source.t11 a_n1496_n2688# 0.259105f
C87 source.t10 a_n1496_n2688# 0.259105f
C88 source.n1 a_n1496_n2688# 1.60777f
C89 source.n2 a_n1496_n2688# 0.310932f
C90 source.t16 a_n1496_n2688# 0.259105f
C91 source.t13 a_n1496_n2688# 0.259105f
C92 source.n3 a_n1496_n2688# 1.60777f
C93 source.n4 a_n1496_n2688# 0.325626f
C94 source.t2 a_n1496_n2688# 1.95824f
C95 source.n5 a_n1496_n2688# 0.441548f
C96 source.t4 a_n1496_n2688# 0.259105f
C97 source.t1 a_n1496_n2688# 0.259105f
C98 source.n6 a_n1496_n2688# 1.60777f
C99 source.n7 a_n1496_n2688# 0.310932f
C100 source.t5 a_n1496_n2688# 0.259105f
C101 source.t19 a_n1496_n2688# 0.259105f
C102 source.n8 a_n1496_n2688# 1.60777f
C103 source.n9 a_n1496_n2688# 1.36964f
C104 source.t12 a_n1496_n2688# 0.259105f
C105 source.t9 a_n1496_n2688# 0.259105f
C106 source.n10 a_n1496_n2688# 1.60777f
C107 source.n11 a_n1496_n2688# 1.36964f
C108 source.t18 a_n1496_n2688# 0.259105f
C109 source.t15 a_n1496_n2688# 0.259105f
C110 source.n12 a_n1496_n2688# 1.60777f
C111 source.n13 a_n1496_n2688# 0.310936f
C112 source.t14 a_n1496_n2688# 1.95823f
C113 source.n14 a_n1496_n2688# 0.441553f
C114 source.t8 a_n1496_n2688# 0.259105f
C115 source.t0 a_n1496_n2688# 0.259105f
C116 source.n15 a_n1496_n2688# 1.60777f
C117 source.n16 a_n1496_n2688# 0.32563f
C118 source.t7 a_n1496_n2688# 0.259105f
C119 source.t3 a_n1496_n2688# 0.259105f
C120 source.n17 a_n1496_n2688# 1.60777f
C121 source.n18 a_n1496_n2688# 0.310936f
C122 source.t6 a_n1496_n2688# 1.95823f
C123 source.n19 a_n1496_n2688# 0.556646f
C124 source.n20 a_n1496_n2688# 1.25241f
C125 plus.n0 a_n1496_n2688# 0.046572f
C126 plus.t6 a_n1496_n2688# 0.178156f
C127 plus.t7 a_n1496_n2688# 0.178156f
C128 plus.n1 a_n1496_n2688# 0.019757f
C129 plus.t5 a_n1496_n2688# 0.180223f
C130 plus.t8 a_n1496_n2688# 0.178156f
C131 plus.n2 a_n1496_n2688# 0.081573f
C132 plus.n3 a_n1496_n2688# 0.09789f
C133 plus.n4 a_n1496_n2688# 0.10026f
C134 plus.n5 a_n1496_n2688# 0.046572f
C135 plus.n6 a_n1496_n2688# 0.097023f
C136 plus.n7 a_n1496_n2688# 0.019757f
C137 plus.n8 a_n1496_n2688# 0.081573f
C138 plus.t9 a_n1496_n2688# 0.180223f
C139 plus.n9 a_n1496_n2688# 0.097827f
C140 plus.n10 a_n1496_n2688# 0.459032f
C141 plus.n11 a_n1496_n2688# 0.046572f
C142 plus.t3 a_n1496_n2688# 0.180223f
C143 plus.t1 a_n1496_n2688# 0.178156f
C144 plus.t0 a_n1496_n2688# 0.178156f
C145 plus.n12 a_n1496_n2688# 0.019757f
C146 plus.t4 a_n1496_n2688# 0.178156f
C147 plus.n13 a_n1496_n2688# 0.081573f
C148 plus.t2 a_n1496_n2688# 0.180223f
C149 plus.n14 a_n1496_n2688# 0.09789f
C150 plus.n15 a_n1496_n2688# 0.10026f
C151 plus.n16 a_n1496_n2688# 0.046572f
C152 plus.n17 a_n1496_n2688# 0.097023f
C153 plus.n18 a_n1496_n2688# 0.019757f
C154 plus.n19 a_n1496_n2688# 0.081573f
C155 plus.n20 a_n1496_n2688# 0.097827f
C156 plus.n21 a_n1496_n2688# 1.20904f
.ends

