* NGSPICE file created from diffpair679.ext - technology: sky130A

.subckt diffpair679 minus drain_right drain_left source plus
X0 source.t47 plus.t0 drain_left.t2 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X1 drain_left.t1 plus.t1 source.t46 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X2 source.t6 minus.t0 drain_right.t23 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X3 drain_right.t22 minus.t1 source.t0 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X4 drain_right.t21 minus.t2 source.t20 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X5 source.t10 minus.t3 drain_right.t20 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X6 source.t14 minus.t4 drain_right.t19 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X7 source.t8 minus.t5 drain_right.t18 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X8 drain_right.t17 minus.t6 source.t19 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X9 source.t45 plus.t2 drain_left.t0 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X10 drain_right.t16 minus.t7 source.t23 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X11 source.t44 plus.t3 drain_left.t5 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X12 drain_left.t4 plus.t4 source.t43 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X13 drain_left.t3 plus.t5 source.t42 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X14 a_n2354_n5888# a_n2354_n5888# a_n2354_n5888# a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.3
X15 drain_right.t15 minus.t8 source.t13 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X16 drain_left.t20 plus.t6 source.t41 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X17 source.t15 minus.t9 drain_right.t14 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X18 drain_left.t19 plus.t7 source.t40 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X19 source.t39 plus.t8 drain_left.t18 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X20 drain_left.t11 plus.t9 source.t38 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X21 source.t7 minus.t10 drain_right.t13 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X22 source.t12 minus.t11 drain_right.t12 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X23 a_n2354_n5888# a_n2354_n5888# a_n2354_n5888# a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X24 source.t16 minus.t12 drain_right.t11 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X25 source.t21 minus.t13 drain_right.t10 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X26 source.t37 plus.t10 drain_left.t10 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X27 source.t36 plus.t11 drain_left.t9 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X28 drain_left.t8 plus.t12 source.t35 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X29 drain_right.t9 minus.t14 source.t2 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X30 drain_left.t7 plus.t13 source.t34 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X31 source.t33 plus.t14 drain_left.t6 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X32 source.t32 plus.t15 drain_left.t14 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X33 source.t31 plus.t16 drain_left.t13 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X34 drain_right.t8 minus.t15 source.t9 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X35 drain_right.t7 minus.t16 source.t11 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X36 drain_left.t12 plus.t17 source.t30 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X37 source.t3 minus.t17 drain_right.t6 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X38 drain_right.t5 minus.t18 source.t1 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X39 drain_right.t4 minus.t19 source.t5 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X40 a_n2354_n5888# a_n2354_n5888# a_n2354_n5888# a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X41 a_n2354_n5888# a_n2354_n5888# a_n2354_n5888# a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X42 drain_right.t3 minus.t20 source.t18 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X43 source.t29 plus.t18 drain_left.t23 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X44 source.t17 minus.t21 drain_right.t2 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X45 source.t22 minus.t22 drain_right.t1 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X46 drain_right.t0 minus.t23 source.t4 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X47 source.t28 plus.t19 drain_left.t22 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X48 source.t27 plus.t20 drain_left.t21 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X49 drain_left.t17 plus.t21 source.t26 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X50 drain_left.t16 plus.t22 source.t25 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X51 drain_left.t15 plus.t23 source.t24 a_n2354_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
R0 plus.n9 plus.t2 2144.17
R1 plus.n35 plus.t5 2144.17
R2 plus.n46 plus.t22 2144.17
R3 plus.n72 plus.t3 2144.17
R4 plus.n8 plus.t9 2112.77
R5 plus.n13 plus.t15 2112.77
R6 plus.n15 plus.t21 2112.77
R7 plus.n5 plus.t8 2112.77
R8 plus.n20 plus.t13 2112.77
R9 plus.n3 plus.t20 2112.77
R10 plus.n26 plus.t1 2112.77
R11 plus.n28 plus.t10 2112.77
R12 plus.n1 plus.t17 2112.77
R13 plus.n34 plus.t0 2112.77
R14 plus.n45 plus.t11 2112.77
R15 plus.n50 plus.t23 2112.77
R16 plus.n52 plus.t14 2112.77
R17 plus.n42 plus.t6 2112.77
R18 plus.n57 plus.t16 2112.77
R19 plus.n40 plus.t7 2112.77
R20 plus.n63 plus.t18 2112.77
R21 plus.n65 plus.t4 2112.77
R22 plus.n38 plus.t19 2112.77
R23 plus.n71 plus.t12 2112.77
R24 plus.n10 plus.n9 161.489
R25 plus.n47 plus.n46 161.489
R26 plus.n10 plus.n7 161.3
R27 plus.n12 plus.n11 161.3
R28 plus.n14 plus.n6 161.3
R29 plus.n17 plus.n16 161.3
R30 plus.n19 plus.n18 161.3
R31 plus.n21 plus.n4 161.3
R32 plus.n23 plus.n22 161.3
R33 plus.n25 plus.n24 161.3
R34 plus.n27 plus.n2 161.3
R35 plus.n30 plus.n29 161.3
R36 plus.n32 plus.n31 161.3
R37 plus.n33 plus.n0 161.3
R38 plus.n36 plus.n35 161.3
R39 plus.n47 plus.n44 161.3
R40 plus.n49 plus.n48 161.3
R41 plus.n51 plus.n43 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n56 plus.n55 161.3
R44 plus.n58 plus.n41 161.3
R45 plus.n60 plus.n59 161.3
R46 plus.n62 plus.n61 161.3
R47 plus.n64 plus.n39 161.3
R48 plus.n67 plus.n66 161.3
R49 plus.n69 plus.n68 161.3
R50 plus.n70 plus.n37 161.3
R51 plus.n73 plus.n72 161.3
R52 plus.n12 plus.n7 73.0308
R53 plus.n22 plus.n21 73.0308
R54 plus.n33 plus.n32 73.0308
R55 plus.n70 plus.n69 73.0308
R56 plus.n59 plus.n58 73.0308
R57 plus.n49 plus.n44 73.0308
R58 plus.n14 plus.n13 66.4581
R59 plus.n29 plus.n1 66.4581
R60 plus.n66 plus.n38 66.4581
R61 plus.n51 plus.n50 66.4581
R62 plus.n20 plus.n19 63.5369
R63 plus.n25 plus.n3 63.5369
R64 plus.n62 plus.n40 63.5369
R65 plus.n57 plus.n56 63.5369
R66 plus.n9 plus.n8 60.6157
R67 plus.n35 plus.n34 60.6157
R68 plus.n72 plus.n71 60.6157
R69 plus.n46 plus.n45 60.6157
R70 plus.n16 plus.n15 47.4702
R71 plus.n28 plus.n27 47.4702
R72 plus.n65 plus.n64 47.4702
R73 plus.n53 plus.n52 47.4702
R74 plus.n16 plus.n5 44.549
R75 plus.n27 plus.n26 44.549
R76 plus.n64 plus.n63 44.549
R77 plus.n53 plus.n42 44.549
R78 plus plus.n73 36.8134
R79 plus.n19 plus.n5 28.4823
R80 plus.n26 plus.n25 28.4823
R81 plus.n63 plus.n62 28.4823
R82 plus.n56 plus.n42 28.4823
R83 plus.n15 plus.n14 25.5611
R84 plus.n29 plus.n28 25.5611
R85 plus.n66 plus.n65 25.5611
R86 plus.n52 plus.n51 25.5611
R87 plus plus.n36 17.0384
R88 plus.n8 plus.n7 12.4157
R89 plus.n34 plus.n33 12.4157
R90 plus.n71 plus.n70 12.4157
R91 plus.n45 plus.n44 12.4157
R92 plus.n21 plus.n20 9.49444
R93 plus.n22 plus.n3 9.49444
R94 plus.n59 plus.n40 9.49444
R95 plus.n58 plus.n57 9.49444
R96 plus.n13 plus.n12 6.57323
R97 plus.n32 plus.n1 6.57323
R98 plus.n69 plus.n38 6.57323
R99 plus.n50 plus.n49 6.57323
R100 plus.n11 plus.n10 0.189894
R101 plus.n11 plus.n6 0.189894
R102 plus.n17 plus.n6 0.189894
R103 plus.n18 plus.n17 0.189894
R104 plus.n18 plus.n4 0.189894
R105 plus.n23 plus.n4 0.189894
R106 plus.n24 plus.n23 0.189894
R107 plus.n24 plus.n2 0.189894
R108 plus.n30 plus.n2 0.189894
R109 plus.n31 plus.n30 0.189894
R110 plus.n31 plus.n0 0.189894
R111 plus.n36 plus.n0 0.189894
R112 plus.n73 plus.n37 0.189894
R113 plus.n68 plus.n37 0.189894
R114 plus.n68 plus.n67 0.189894
R115 plus.n67 plus.n39 0.189894
R116 plus.n61 plus.n39 0.189894
R117 plus.n61 plus.n60 0.189894
R118 plus.n60 plus.n41 0.189894
R119 plus.n55 plus.n41 0.189894
R120 plus.n55 plus.n54 0.189894
R121 plus.n54 plus.n43 0.189894
R122 plus.n48 plus.n43 0.189894
R123 plus.n48 plus.n47 0.189894
R124 drain_left.n7 drain_left.n5 59.2585
R125 drain_left.n2 drain_left.n0 59.2585
R126 drain_left.n13 drain_left.n11 59.2585
R127 drain_left.n7 drain_left.n6 58.7154
R128 drain_left.n9 drain_left.n8 58.7154
R129 drain_left.n4 drain_left.n3 58.7154
R130 drain_left.n2 drain_left.n1 58.7154
R131 drain_left.n19 drain_left.n18 58.7154
R132 drain_left.n17 drain_left.n16 58.7154
R133 drain_left.n15 drain_left.n14 58.7154
R134 drain_left.n13 drain_left.n12 58.7154
R135 drain_left.n21 drain_left.n20 58.7153
R136 drain_left drain_left.n10 42.375
R137 drain_left drain_left.n21 6.19632
R138 drain_left.n5 drain_left.t9 0.7925
R139 drain_left.n5 drain_left.t16 0.7925
R140 drain_left.n6 drain_left.t6 0.7925
R141 drain_left.n6 drain_left.t15 0.7925
R142 drain_left.n8 drain_left.t13 0.7925
R143 drain_left.n8 drain_left.t20 0.7925
R144 drain_left.n3 drain_left.t23 0.7925
R145 drain_left.n3 drain_left.t19 0.7925
R146 drain_left.n1 drain_left.t22 0.7925
R147 drain_left.n1 drain_left.t4 0.7925
R148 drain_left.n0 drain_left.t5 0.7925
R149 drain_left.n0 drain_left.t8 0.7925
R150 drain_left.n20 drain_left.t2 0.7925
R151 drain_left.n20 drain_left.t3 0.7925
R152 drain_left.n18 drain_left.t10 0.7925
R153 drain_left.n18 drain_left.t12 0.7925
R154 drain_left.n16 drain_left.t21 0.7925
R155 drain_left.n16 drain_left.t1 0.7925
R156 drain_left.n14 drain_left.t18 0.7925
R157 drain_left.n14 drain_left.t7 0.7925
R158 drain_left.n12 drain_left.t14 0.7925
R159 drain_left.n12 drain_left.t17 0.7925
R160 drain_left.n11 drain_left.t0 0.7925
R161 drain_left.n11 drain_left.t11 0.7925
R162 drain_left.n9 drain_left.n7 0.543603
R163 drain_left.n4 drain_left.n2 0.543603
R164 drain_left.n15 drain_left.n13 0.543603
R165 drain_left.n17 drain_left.n15 0.543603
R166 drain_left.n19 drain_left.n17 0.543603
R167 drain_left.n21 drain_left.n19 0.543603
R168 drain_left.n10 drain_left.n9 0.216706
R169 drain_left.n10 drain_left.n4 0.216706
R170 source.n1154 source.n1020 289.615
R171 source.n1004 source.n870 289.615
R172 source.n864 source.n730 289.615
R173 source.n714 source.n580 289.615
R174 source.n134 source.n0 289.615
R175 source.n284 source.n150 289.615
R176 source.n424 source.n290 289.615
R177 source.n574 source.n440 289.615
R178 source.n1064 source.n1063 185
R179 source.n1069 source.n1068 185
R180 source.n1071 source.n1070 185
R181 source.n1060 source.n1059 185
R182 source.n1077 source.n1076 185
R183 source.n1079 source.n1078 185
R184 source.n1056 source.n1055 185
R185 source.n1086 source.n1085 185
R186 source.n1087 source.n1054 185
R187 source.n1089 source.n1088 185
R188 source.n1052 source.n1051 185
R189 source.n1095 source.n1094 185
R190 source.n1097 source.n1096 185
R191 source.n1048 source.n1047 185
R192 source.n1103 source.n1102 185
R193 source.n1105 source.n1104 185
R194 source.n1044 source.n1043 185
R195 source.n1111 source.n1110 185
R196 source.n1113 source.n1112 185
R197 source.n1040 source.n1039 185
R198 source.n1119 source.n1118 185
R199 source.n1121 source.n1120 185
R200 source.n1036 source.n1035 185
R201 source.n1127 source.n1126 185
R202 source.n1130 source.n1129 185
R203 source.n1128 source.n1032 185
R204 source.n1135 source.n1031 185
R205 source.n1137 source.n1136 185
R206 source.n1139 source.n1138 185
R207 source.n1028 source.n1027 185
R208 source.n1145 source.n1144 185
R209 source.n1147 source.n1146 185
R210 source.n1024 source.n1023 185
R211 source.n1153 source.n1152 185
R212 source.n1155 source.n1154 185
R213 source.n914 source.n913 185
R214 source.n919 source.n918 185
R215 source.n921 source.n920 185
R216 source.n910 source.n909 185
R217 source.n927 source.n926 185
R218 source.n929 source.n928 185
R219 source.n906 source.n905 185
R220 source.n936 source.n935 185
R221 source.n937 source.n904 185
R222 source.n939 source.n938 185
R223 source.n902 source.n901 185
R224 source.n945 source.n944 185
R225 source.n947 source.n946 185
R226 source.n898 source.n897 185
R227 source.n953 source.n952 185
R228 source.n955 source.n954 185
R229 source.n894 source.n893 185
R230 source.n961 source.n960 185
R231 source.n963 source.n962 185
R232 source.n890 source.n889 185
R233 source.n969 source.n968 185
R234 source.n971 source.n970 185
R235 source.n886 source.n885 185
R236 source.n977 source.n976 185
R237 source.n980 source.n979 185
R238 source.n978 source.n882 185
R239 source.n985 source.n881 185
R240 source.n987 source.n986 185
R241 source.n989 source.n988 185
R242 source.n878 source.n877 185
R243 source.n995 source.n994 185
R244 source.n997 source.n996 185
R245 source.n874 source.n873 185
R246 source.n1003 source.n1002 185
R247 source.n1005 source.n1004 185
R248 source.n774 source.n773 185
R249 source.n779 source.n778 185
R250 source.n781 source.n780 185
R251 source.n770 source.n769 185
R252 source.n787 source.n786 185
R253 source.n789 source.n788 185
R254 source.n766 source.n765 185
R255 source.n796 source.n795 185
R256 source.n797 source.n764 185
R257 source.n799 source.n798 185
R258 source.n762 source.n761 185
R259 source.n805 source.n804 185
R260 source.n807 source.n806 185
R261 source.n758 source.n757 185
R262 source.n813 source.n812 185
R263 source.n815 source.n814 185
R264 source.n754 source.n753 185
R265 source.n821 source.n820 185
R266 source.n823 source.n822 185
R267 source.n750 source.n749 185
R268 source.n829 source.n828 185
R269 source.n831 source.n830 185
R270 source.n746 source.n745 185
R271 source.n837 source.n836 185
R272 source.n840 source.n839 185
R273 source.n838 source.n742 185
R274 source.n845 source.n741 185
R275 source.n847 source.n846 185
R276 source.n849 source.n848 185
R277 source.n738 source.n737 185
R278 source.n855 source.n854 185
R279 source.n857 source.n856 185
R280 source.n734 source.n733 185
R281 source.n863 source.n862 185
R282 source.n865 source.n864 185
R283 source.n624 source.n623 185
R284 source.n629 source.n628 185
R285 source.n631 source.n630 185
R286 source.n620 source.n619 185
R287 source.n637 source.n636 185
R288 source.n639 source.n638 185
R289 source.n616 source.n615 185
R290 source.n646 source.n645 185
R291 source.n647 source.n614 185
R292 source.n649 source.n648 185
R293 source.n612 source.n611 185
R294 source.n655 source.n654 185
R295 source.n657 source.n656 185
R296 source.n608 source.n607 185
R297 source.n663 source.n662 185
R298 source.n665 source.n664 185
R299 source.n604 source.n603 185
R300 source.n671 source.n670 185
R301 source.n673 source.n672 185
R302 source.n600 source.n599 185
R303 source.n679 source.n678 185
R304 source.n681 source.n680 185
R305 source.n596 source.n595 185
R306 source.n687 source.n686 185
R307 source.n690 source.n689 185
R308 source.n688 source.n592 185
R309 source.n695 source.n591 185
R310 source.n697 source.n696 185
R311 source.n699 source.n698 185
R312 source.n588 source.n587 185
R313 source.n705 source.n704 185
R314 source.n707 source.n706 185
R315 source.n584 source.n583 185
R316 source.n713 source.n712 185
R317 source.n715 source.n714 185
R318 source.n135 source.n134 185
R319 source.n133 source.n132 185
R320 source.n4 source.n3 185
R321 source.n127 source.n126 185
R322 source.n125 source.n124 185
R323 source.n8 source.n7 185
R324 source.n119 source.n118 185
R325 source.n117 source.n116 185
R326 source.n115 source.n11 185
R327 source.n15 source.n12 185
R328 source.n110 source.n109 185
R329 source.n108 source.n107 185
R330 source.n17 source.n16 185
R331 source.n102 source.n101 185
R332 source.n100 source.n99 185
R333 source.n21 source.n20 185
R334 source.n94 source.n93 185
R335 source.n92 source.n91 185
R336 source.n25 source.n24 185
R337 source.n86 source.n85 185
R338 source.n84 source.n83 185
R339 source.n29 source.n28 185
R340 source.n78 source.n77 185
R341 source.n76 source.n75 185
R342 source.n33 source.n32 185
R343 source.n70 source.n69 185
R344 source.n68 source.n35 185
R345 source.n67 source.n66 185
R346 source.n38 source.n36 185
R347 source.n61 source.n60 185
R348 source.n59 source.n58 185
R349 source.n42 source.n41 185
R350 source.n53 source.n52 185
R351 source.n51 source.n50 185
R352 source.n46 source.n45 185
R353 source.n285 source.n284 185
R354 source.n283 source.n282 185
R355 source.n154 source.n153 185
R356 source.n277 source.n276 185
R357 source.n275 source.n274 185
R358 source.n158 source.n157 185
R359 source.n269 source.n268 185
R360 source.n267 source.n266 185
R361 source.n265 source.n161 185
R362 source.n165 source.n162 185
R363 source.n260 source.n259 185
R364 source.n258 source.n257 185
R365 source.n167 source.n166 185
R366 source.n252 source.n251 185
R367 source.n250 source.n249 185
R368 source.n171 source.n170 185
R369 source.n244 source.n243 185
R370 source.n242 source.n241 185
R371 source.n175 source.n174 185
R372 source.n236 source.n235 185
R373 source.n234 source.n233 185
R374 source.n179 source.n178 185
R375 source.n228 source.n227 185
R376 source.n226 source.n225 185
R377 source.n183 source.n182 185
R378 source.n220 source.n219 185
R379 source.n218 source.n185 185
R380 source.n217 source.n216 185
R381 source.n188 source.n186 185
R382 source.n211 source.n210 185
R383 source.n209 source.n208 185
R384 source.n192 source.n191 185
R385 source.n203 source.n202 185
R386 source.n201 source.n200 185
R387 source.n196 source.n195 185
R388 source.n425 source.n424 185
R389 source.n423 source.n422 185
R390 source.n294 source.n293 185
R391 source.n417 source.n416 185
R392 source.n415 source.n414 185
R393 source.n298 source.n297 185
R394 source.n409 source.n408 185
R395 source.n407 source.n406 185
R396 source.n405 source.n301 185
R397 source.n305 source.n302 185
R398 source.n400 source.n399 185
R399 source.n398 source.n397 185
R400 source.n307 source.n306 185
R401 source.n392 source.n391 185
R402 source.n390 source.n389 185
R403 source.n311 source.n310 185
R404 source.n384 source.n383 185
R405 source.n382 source.n381 185
R406 source.n315 source.n314 185
R407 source.n376 source.n375 185
R408 source.n374 source.n373 185
R409 source.n319 source.n318 185
R410 source.n368 source.n367 185
R411 source.n366 source.n365 185
R412 source.n323 source.n322 185
R413 source.n360 source.n359 185
R414 source.n358 source.n325 185
R415 source.n357 source.n356 185
R416 source.n328 source.n326 185
R417 source.n351 source.n350 185
R418 source.n349 source.n348 185
R419 source.n332 source.n331 185
R420 source.n343 source.n342 185
R421 source.n341 source.n340 185
R422 source.n336 source.n335 185
R423 source.n575 source.n574 185
R424 source.n573 source.n572 185
R425 source.n444 source.n443 185
R426 source.n567 source.n566 185
R427 source.n565 source.n564 185
R428 source.n448 source.n447 185
R429 source.n559 source.n558 185
R430 source.n557 source.n556 185
R431 source.n555 source.n451 185
R432 source.n455 source.n452 185
R433 source.n550 source.n549 185
R434 source.n548 source.n547 185
R435 source.n457 source.n456 185
R436 source.n542 source.n541 185
R437 source.n540 source.n539 185
R438 source.n461 source.n460 185
R439 source.n534 source.n533 185
R440 source.n532 source.n531 185
R441 source.n465 source.n464 185
R442 source.n526 source.n525 185
R443 source.n524 source.n523 185
R444 source.n469 source.n468 185
R445 source.n518 source.n517 185
R446 source.n516 source.n515 185
R447 source.n473 source.n472 185
R448 source.n510 source.n509 185
R449 source.n508 source.n475 185
R450 source.n507 source.n506 185
R451 source.n478 source.n476 185
R452 source.n501 source.n500 185
R453 source.n499 source.n498 185
R454 source.n482 source.n481 185
R455 source.n493 source.n492 185
R456 source.n491 source.n490 185
R457 source.n486 source.n485 185
R458 source.n1065 source.t23 149.524
R459 source.n915 source.t8 149.524
R460 source.n775 source.t25 149.524
R461 source.n625 source.t44 149.524
R462 source.n47 source.t42 149.524
R463 source.n197 source.t45 149.524
R464 source.n337 source.t2 149.524
R465 source.n487 source.t10 149.524
R466 source.n1069 source.n1063 104.615
R467 source.n1070 source.n1069 104.615
R468 source.n1070 source.n1059 104.615
R469 source.n1077 source.n1059 104.615
R470 source.n1078 source.n1077 104.615
R471 source.n1078 source.n1055 104.615
R472 source.n1086 source.n1055 104.615
R473 source.n1087 source.n1086 104.615
R474 source.n1088 source.n1087 104.615
R475 source.n1088 source.n1051 104.615
R476 source.n1095 source.n1051 104.615
R477 source.n1096 source.n1095 104.615
R478 source.n1096 source.n1047 104.615
R479 source.n1103 source.n1047 104.615
R480 source.n1104 source.n1103 104.615
R481 source.n1104 source.n1043 104.615
R482 source.n1111 source.n1043 104.615
R483 source.n1112 source.n1111 104.615
R484 source.n1112 source.n1039 104.615
R485 source.n1119 source.n1039 104.615
R486 source.n1120 source.n1119 104.615
R487 source.n1120 source.n1035 104.615
R488 source.n1127 source.n1035 104.615
R489 source.n1129 source.n1127 104.615
R490 source.n1129 source.n1128 104.615
R491 source.n1128 source.n1031 104.615
R492 source.n1137 source.n1031 104.615
R493 source.n1138 source.n1137 104.615
R494 source.n1138 source.n1027 104.615
R495 source.n1145 source.n1027 104.615
R496 source.n1146 source.n1145 104.615
R497 source.n1146 source.n1023 104.615
R498 source.n1153 source.n1023 104.615
R499 source.n1154 source.n1153 104.615
R500 source.n919 source.n913 104.615
R501 source.n920 source.n919 104.615
R502 source.n920 source.n909 104.615
R503 source.n927 source.n909 104.615
R504 source.n928 source.n927 104.615
R505 source.n928 source.n905 104.615
R506 source.n936 source.n905 104.615
R507 source.n937 source.n936 104.615
R508 source.n938 source.n937 104.615
R509 source.n938 source.n901 104.615
R510 source.n945 source.n901 104.615
R511 source.n946 source.n945 104.615
R512 source.n946 source.n897 104.615
R513 source.n953 source.n897 104.615
R514 source.n954 source.n953 104.615
R515 source.n954 source.n893 104.615
R516 source.n961 source.n893 104.615
R517 source.n962 source.n961 104.615
R518 source.n962 source.n889 104.615
R519 source.n969 source.n889 104.615
R520 source.n970 source.n969 104.615
R521 source.n970 source.n885 104.615
R522 source.n977 source.n885 104.615
R523 source.n979 source.n977 104.615
R524 source.n979 source.n978 104.615
R525 source.n978 source.n881 104.615
R526 source.n987 source.n881 104.615
R527 source.n988 source.n987 104.615
R528 source.n988 source.n877 104.615
R529 source.n995 source.n877 104.615
R530 source.n996 source.n995 104.615
R531 source.n996 source.n873 104.615
R532 source.n1003 source.n873 104.615
R533 source.n1004 source.n1003 104.615
R534 source.n779 source.n773 104.615
R535 source.n780 source.n779 104.615
R536 source.n780 source.n769 104.615
R537 source.n787 source.n769 104.615
R538 source.n788 source.n787 104.615
R539 source.n788 source.n765 104.615
R540 source.n796 source.n765 104.615
R541 source.n797 source.n796 104.615
R542 source.n798 source.n797 104.615
R543 source.n798 source.n761 104.615
R544 source.n805 source.n761 104.615
R545 source.n806 source.n805 104.615
R546 source.n806 source.n757 104.615
R547 source.n813 source.n757 104.615
R548 source.n814 source.n813 104.615
R549 source.n814 source.n753 104.615
R550 source.n821 source.n753 104.615
R551 source.n822 source.n821 104.615
R552 source.n822 source.n749 104.615
R553 source.n829 source.n749 104.615
R554 source.n830 source.n829 104.615
R555 source.n830 source.n745 104.615
R556 source.n837 source.n745 104.615
R557 source.n839 source.n837 104.615
R558 source.n839 source.n838 104.615
R559 source.n838 source.n741 104.615
R560 source.n847 source.n741 104.615
R561 source.n848 source.n847 104.615
R562 source.n848 source.n737 104.615
R563 source.n855 source.n737 104.615
R564 source.n856 source.n855 104.615
R565 source.n856 source.n733 104.615
R566 source.n863 source.n733 104.615
R567 source.n864 source.n863 104.615
R568 source.n629 source.n623 104.615
R569 source.n630 source.n629 104.615
R570 source.n630 source.n619 104.615
R571 source.n637 source.n619 104.615
R572 source.n638 source.n637 104.615
R573 source.n638 source.n615 104.615
R574 source.n646 source.n615 104.615
R575 source.n647 source.n646 104.615
R576 source.n648 source.n647 104.615
R577 source.n648 source.n611 104.615
R578 source.n655 source.n611 104.615
R579 source.n656 source.n655 104.615
R580 source.n656 source.n607 104.615
R581 source.n663 source.n607 104.615
R582 source.n664 source.n663 104.615
R583 source.n664 source.n603 104.615
R584 source.n671 source.n603 104.615
R585 source.n672 source.n671 104.615
R586 source.n672 source.n599 104.615
R587 source.n679 source.n599 104.615
R588 source.n680 source.n679 104.615
R589 source.n680 source.n595 104.615
R590 source.n687 source.n595 104.615
R591 source.n689 source.n687 104.615
R592 source.n689 source.n688 104.615
R593 source.n688 source.n591 104.615
R594 source.n697 source.n591 104.615
R595 source.n698 source.n697 104.615
R596 source.n698 source.n587 104.615
R597 source.n705 source.n587 104.615
R598 source.n706 source.n705 104.615
R599 source.n706 source.n583 104.615
R600 source.n713 source.n583 104.615
R601 source.n714 source.n713 104.615
R602 source.n134 source.n133 104.615
R603 source.n133 source.n3 104.615
R604 source.n126 source.n3 104.615
R605 source.n126 source.n125 104.615
R606 source.n125 source.n7 104.615
R607 source.n118 source.n7 104.615
R608 source.n118 source.n117 104.615
R609 source.n117 source.n11 104.615
R610 source.n15 source.n11 104.615
R611 source.n109 source.n15 104.615
R612 source.n109 source.n108 104.615
R613 source.n108 source.n16 104.615
R614 source.n101 source.n16 104.615
R615 source.n101 source.n100 104.615
R616 source.n100 source.n20 104.615
R617 source.n93 source.n20 104.615
R618 source.n93 source.n92 104.615
R619 source.n92 source.n24 104.615
R620 source.n85 source.n24 104.615
R621 source.n85 source.n84 104.615
R622 source.n84 source.n28 104.615
R623 source.n77 source.n28 104.615
R624 source.n77 source.n76 104.615
R625 source.n76 source.n32 104.615
R626 source.n69 source.n32 104.615
R627 source.n69 source.n68 104.615
R628 source.n68 source.n67 104.615
R629 source.n67 source.n36 104.615
R630 source.n60 source.n36 104.615
R631 source.n60 source.n59 104.615
R632 source.n59 source.n41 104.615
R633 source.n52 source.n41 104.615
R634 source.n52 source.n51 104.615
R635 source.n51 source.n45 104.615
R636 source.n284 source.n283 104.615
R637 source.n283 source.n153 104.615
R638 source.n276 source.n153 104.615
R639 source.n276 source.n275 104.615
R640 source.n275 source.n157 104.615
R641 source.n268 source.n157 104.615
R642 source.n268 source.n267 104.615
R643 source.n267 source.n161 104.615
R644 source.n165 source.n161 104.615
R645 source.n259 source.n165 104.615
R646 source.n259 source.n258 104.615
R647 source.n258 source.n166 104.615
R648 source.n251 source.n166 104.615
R649 source.n251 source.n250 104.615
R650 source.n250 source.n170 104.615
R651 source.n243 source.n170 104.615
R652 source.n243 source.n242 104.615
R653 source.n242 source.n174 104.615
R654 source.n235 source.n174 104.615
R655 source.n235 source.n234 104.615
R656 source.n234 source.n178 104.615
R657 source.n227 source.n178 104.615
R658 source.n227 source.n226 104.615
R659 source.n226 source.n182 104.615
R660 source.n219 source.n182 104.615
R661 source.n219 source.n218 104.615
R662 source.n218 source.n217 104.615
R663 source.n217 source.n186 104.615
R664 source.n210 source.n186 104.615
R665 source.n210 source.n209 104.615
R666 source.n209 source.n191 104.615
R667 source.n202 source.n191 104.615
R668 source.n202 source.n201 104.615
R669 source.n201 source.n195 104.615
R670 source.n424 source.n423 104.615
R671 source.n423 source.n293 104.615
R672 source.n416 source.n293 104.615
R673 source.n416 source.n415 104.615
R674 source.n415 source.n297 104.615
R675 source.n408 source.n297 104.615
R676 source.n408 source.n407 104.615
R677 source.n407 source.n301 104.615
R678 source.n305 source.n301 104.615
R679 source.n399 source.n305 104.615
R680 source.n399 source.n398 104.615
R681 source.n398 source.n306 104.615
R682 source.n391 source.n306 104.615
R683 source.n391 source.n390 104.615
R684 source.n390 source.n310 104.615
R685 source.n383 source.n310 104.615
R686 source.n383 source.n382 104.615
R687 source.n382 source.n314 104.615
R688 source.n375 source.n314 104.615
R689 source.n375 source.n374 104.615
R690 source.n374 source.n318 104.615
R691 source.n367 source.n318 104.615
R692 source.n367 source.n366 104.615
R693 source.n366 source.n322 104.615
R694 source.n359 source.n322 104.615
R695 source.n359 source.n358 104.615
R696 source.n358 source.n357 104.615
R697 source.n357 source.n326 104.615
R698 source.n350 source.n326 104.615
R699 source.n350 source.n349 104.615
R700 source.n349 source.n331 104.615
R701 source.n342 source.n331 104.615
R702 source.n342 source.n341 104.615
R703 source.n341 source.n335 104.615
R704 source.n574 source.n573 104.615
R705 source.n573 source.n443 104.615
R706 source.n566 source.n443 104.615
R707 source.n566 source.n565 104.615
R708 source.n565 source.n447 104.615
R709 source.n558 source.n447 104.615
R710 source.n558 source.n557 104.615
R711 source.n557 source.n451 104.615
R712 source.n455 source.n451 104.615
R713 source.n549 source.n455 104.615
R714 source.n549 source.n548 104.615
R715 source.n548 source.n456 104.615
R716 source.n541 source.n456 104.615
R717 source.n541 source.n540 104.615
R718 source.n540 source.n460 104.615
R719 source.n533 source.n460 104.615
R720 source.n533 source.n532 104.615
R721 source.n532 source.n464 104.615
R722 source.n525 source.n464 104.615
R723 source.n525 source.n524 104.615
R724 source.n524 source.n468 104.615
R725 source.n517 source.n468 104.615
R726 source.n517 source.n516 104.615
R727 source.n516 source.n472 104.615
R728 source.n509 source.n472 104.615
R729 source.n509 source.n508 104.615
R730 source.n508 source.n507 104.615
R731 source.n507 source.n476 104.615
R732 source.n500 source.n476 104.615
R733 source.n500 source.n499 104.615
R734 source.n499 source.n481 104.615
R735 source.n492 source.n481 104.615
R736 source.n492 source.n491 104.615
R737 source.n491 source.n485 104.615
R738 source.t23 source.n1063 52.3082
R739 source.t8 source.n913 52.3082
R740 source.t25 source.n773 52.3082
R741 source.t44 source.n623 52.3082
R742 source.t42 source.n45 52.3082
R743 source.t45 source.n195 52.3082
R744 source.t2 source.n335 52.3082
R745 source.t10 source.n485 52.3082
R746 source.n1019 source.n1018 42.0366
R747 source.n1017 source.n1016 42.0366
R748 source.n1015 source.n1014 42.0366
R749 source.n1013 source.n1012 42.0366
R750 source.n1011 source.n1010 42.0366
R751 source.n729 source.n728 42.0366
R752 source.n727 source.n726 42.0366
R753 source.n725 source.n724 42.0366
R754 source.n723 source.n722 42.0366
R755 source.n721 source.n720 42.0366
R756 source.n141 source.n140 42.0366
R757 source.n143 source.n142 42.0366
R758 source.n145 source.n144 42.0366
R759 source.n147 source.n146 42.0366
R760 source.n149 source.n148 42.0366
R761 source.n431 source.n430 42.0366
R762 source.n433 source.n432 42.0366
R763 source.n435 source.n434 42.0366
R764 source.n437 source.n436 42.0366
R765 source.n439 source.n438 42.0366
R766 source.n719 source.n579 31.6793
R767 source.n1159 source.n1158 30.6338
R768 source.n1009 source.n1008 30.6338
R769 source.n869 source.n868 30.6338
R770 source.n719 source.n718 30.6338
R771 source.n139 source.n138 30.6338
R772 source.n289 source.n288 30.6338
R773 source.n429 source.n428 30.6338
R774 source.n579 source.n578 30.6338
R775 source.n1160 source.n139 26.1448
R776 source.n1089 source.n1054 13.1884
R777 source.n1136 source.n1135 13.1884
R778 source.n939 source.n904 13.1884
R779 source.n986 source.n985 13.1884
R780 source.n799 source.n764 13.1884
R781 source.n846 source.n845 13.1884
R782 source.n649 source.n614 13.1884
R783 source.n696 source.n695 13.1884
R784 source.n116 source.n115 13.1884
R785 source.n70 source.n35 13.1884
R786 source.n266 source.n265 13.1884
R787 source.n220 source.n185 13.1884
R788 source.n406 source.n405 13.1884
R789 source.n360 source.n325 13.1884
R790 source.n556 source.n555 13.1884
R791 source.n510 source.n475 13.1884
R792 source.n1085 source.n1084 12.8005
R793 source.n1090 source.n1052 12.8005
R794 source.n1134 source.n1032 12.8005
R795 source.n1139 source.n1030 12.8005
R796 source.n935 source.n934 12.8005
R797 source.n940 source.n902 12.8005
R798 source.n984 source.n882 12.8005
R799 source.n989 source.n880 12.8005
R800 source.n795 source.n794 12.8005
R801 source.n800 source.n762 12.8005
R802 source.n844 source.n742 12.8005
R803 source.n849 source.n740 12.8005
R804 source.n645 source.n644 12.8005
R805 source.n650 source.n612 12.8005
R806 source.n694 source.n592 12.8005
R807 source.n699 source.n590 12.8005
R808 source.n119 source.n10 12.8005
R809 source.n114 source.n12 12.8005
R810 source.n71 source.n33 12.8005
R811 source.n66 source.n37 12.8005
R812 source.n269 source.n160 12.8005
R813 source.n264 source.n162 12.8005
R814 source.n221 source.n183 12.8005
R815 source.n216 source.n187 12.8005
R816 source.n409 source.n300 12.8005
R817 source.n404 source.n302 12.8005
R818 source.n361 source.n323 12.8005
R819 source.n356 source.n327 12.8005
R820 source.n559 source.n450 12.8005
R821 source.n554 source.n452 12.8005
R822 source.n511 source.n473 12.8005
R823 source.n506 source.n477 12.8005
R824 source.n1083 source.n1056 12.0247
R825 source.n1094 source.n1093 12.0247
R826 source.n1131 source.n1130 12.0247
R827 source.n1140 source.n1028 12.0247
R828 source.n933 source.n906 12.0247
R829 source.n944 source.n943 12.0247
R830 source.n981 source.n980 12.0247
R831 source.n990 source.n878 12.0247
R832 source.n793 source.n766 12.0247
R833 source.n804 source.n803 12.0247
R834 source.n841 source.n840 12.0247
R835 source.n850 source.n738 12.0247
R836 source.n643 source.n616 12.0247
R837 source.n654 source.n653 12.0247
R838 source.n691 source.n690 12.0247
R839 source.n700 source.n588 12.0247
R840 source.n120 source.n8 12.0247
R841 source.n111 source.n110 12.0247
R842 source.n75 source.n74 12.0247
R843 source.n65 source.n38 12.0247
R844 source.n270 source.n158 12.0247
R845 source.n261 source.n260 12.0247
R846 source.n225 source.n224 12.0247
R847 source.n215 source.n188 12.0247
R848 source.n410 source.n298 12.0247
R849 source.n401 source.n400 12.0247
R850 source.n365 source.n364 12.0247
R851 source.n355 source.n328 12.0247
R852 source.n560 source.n448 12.0247
R853 source.n551 source.n550 12.0247
R854 source.n515 source.n514 12.0247
R855 source.n505 source.n478 12.0247
R856 source.n1080 source.n1079 11.249
R857 source.n1097 source.n1050 11.249
R858 source.n1126 source.n1034 11.249
R859 source.n1144 source.n1143 11.249
R860 source.n930 source.n929 11.249
R861 source.n947 source.n900 11.249
R862 source.n976 source.n884 11.249
R863 source.n994 source.n993 11.249
R864 source.n790 source.n789 11.249
R865 source.n807 source.n760 11.249
R866 source.n836 source.n744 11.249
R867 source.n854 source.n853 11.249
R868 source.n640 source.n639 11.249
R869 source.n657 source.n610 11.249
R870 source.n686 source.n594 11.249
R871 source.n704 source.n703 11.249
R872 source.n124 source.n123 11.249
R873 source.n107 source.n14 11.249
R874 source.n78 source.n31 11.249
R875 source.n62 source.n61 11.249
R876 source.n274 source.n273 11.249
R877 source.n257 source.n164 11.249
R878 source.n228 source.n181 11.249
R879 source.n212 source.n211 11.249
R880 source.n414 source.n413 11.249
R881 source.n397 source.n304 11.249
R882 source.n368 source.n321 11.249
R883 source.n352 source.n351 11.249
R884 source.n564 source.n563 11.249
R885 source.n547 source.n454 11.249
R886 source.n518 source.n471 11.249
R887 source.n502 source.n501 11.249
R888 source.n1076 source.n1058 10.4732
R889 source.n1098 source.n1048 10.4732
R890 source.n1125 source.n1036 10.4732
R891 source.n1147 source.n1026 10.4732
R892 source.n926 source.n908 10.4732
R893 source.n948 source.n898 10.4732
R894 source.n975 source.n886 10.4732
R895 source.n997 source.n876 10.4732
R896 source.n786 source.n768 10.4732
R897 source.n808 source.n758 10.4732
R898 source.n835 source.n746 10.4732
R899 source.n857 source.n736 10.4732
R900 source.n636 source.n618 10.4732
R901 source.n658 source.n608 10.4732
R902 source.n685 source.n596 10.4732
R903 source.n707 source.n586 10.4732
R904 source.n127 source.n6 10.4732
R905 source.n106 source.n17 10.4732
R906 source.n79 source.n29 10.4732
R907 source.n58 source.n40 10.4732
R908 source.n277 source.n156 10.4732
R909 source.n256 source.n167 10.4732
R910 source.n229 source.n179 10.4732
R911 source.n208 source.n190 10.4732
R912 source.n417 source.n296 10.4732
R913 source.n396 source.n307 10.4732
R914 source.n369 source.n319 10.4732
R915 source.n348 source.n330 10.4732
R916 source.n567 source.n446 10.4732
R917 source.n546 source.n457 10.4732
R918 source.n519 source.n469 10.4732
R919 source.n498 source.n480 10.4732
R920 source.n1065 source.n1064 10.2747
R921 source.n915 source.n914 10.2747
R922 source.n775 source.n774 10.2747
R923 source.n625 source.n624 10.2747
R924 source.n47 source.n46 10.2747
R925 source.n197 source.n196 10.2747
R926 source.n337 source.n336 10.2747
R927 source.n487 source.n486 10.2747
R928 source.n1075 source.n1060 9.69747
R929 source.n1102 source.n1101 9.69747
R930 source.n1122 source.n1121 9.69747
R931 source.n1148 source.n1024 9.69747
R932 source.n925 source.n910 9.69747
R933 source.n952 source.n951 9.69747
R934 source.n972 source.n971 9.69747
R935 source.n998 source.n874 9.69747
R936 source.n785 source.n770 9.69747
R937 source.n812 source.n811 9.69747
R938 source.n832 source.n831 9.69747
R939 source.n858 source.n734 9.69747
R940 source.n635 source.n620 9.69747
R941 source.n662 source.n661 9.69747
R942 source.n682 source.n681 9.69747
R943 source.n708 source.n584 9.69747
R944 source.n128 source.n4 9.69747
R945 source.n103 source.n102 9.69747
R946 source.n83 source.n82 9.69747
R947 source.n57 source.n42 9.69747
R948 source.n278 source.n154 9.69747
R949 source.n253 source.n252 9.69747
R950 source.n233 source.n232 9.69747
R951 source.n207 source.n192 9.69747
R952 source.n418 source.n294 9.69747
R953 source.n393 source.n392 9.69747
R954 source.n373 source.n372 9.69747
R955 source.n347 source.n332 9.69747
R956 source.n568 source.n444 9.69747
R957 source.n543 source.n542 9.69747
R958 source.n523 source.n522 9.69747
R959 source.n497 source.n482 9.69747
R960 source.n1158 source.n1157 9.45567
R961 source.n1008 source.n1007 9.45567
R962 source.n868 source.n867 9.45567
R963 source.n718 source.n717 9.45567
R964 source.n138 source.n137 9.45567
R965 source.n288 source.n287 9.45567
R966 source.n428 source.n427 9.45567
R967 source.n578 source.n577 9.45567
R968 source.n1022 source.n1021 9.3005
R969 source.n1151 source.n1150 9.3005
R970 source.n1149 source.n1148 9.3005
R971 source.n1026 source.n1025 9.3005
R972 source.n1143 source.n1142 9.3005
R973 source.n1141 source.n1140 9.3005
R974 source.n1030 source.n1029 9.3005
R975 source.n1109 source.n1108 9.3005
R976 source.n1107 source.n1106 9.3005
R977 source.n1046 source.n1045 9.3005
R978 source.n1101 source.n1100 9.3005
R979 source.n1099 source.n1098 9.3005
R980 source.n1050 source.n1049 9.3005
R981 source.n1093 source.n1092 9.3005
R982 source.n1091 source.n1090 9.3005
R983 source.n1067 source.n1066 9.3005
R984 source.n1062 source.n1061 9.3005
R985 source.n1073 source.n1072 9.3005
R986 source.n1075 source.n1074 9.3005
R987 source.n1058 source.n1057 9.3005
R988 source.n1081 source.n1080 9.3005
R989 source.n1083 source.n1082 9.3005
R990 source.n1084 source.n1053 9.3005
R991 source.n1042 source.n1041 9.3005
R992 source.n1115 source.n1114 9.3005
R993 source.n1117 source.n1116 9.3005
R994 source.n1038 source.n1037 9.3005
R995 source.n1123 source.n1122 9.3005
R996 source.n1125 source.n1124 9.3005
R997 source.n1034 source.n1033 9.3005
R998 source.n1132 source.n1131 9.3005
R999 source.n1134 source.n1133 9.3005
R1000 source.n1157 source.n1156 9.3005
R1001 source.n872 source.n871 9.3005
R1002 source.n1001 source.n1000 9.3005
R1003 source.n999 source.n998 9.3005
R1004 source.n876 source.n875 9.3005
R1005 source.n993 source.n992 9.3005
R1006 source.n991 source.n990 9.3005
R1007 source.n880 source.n879 9.3005
R1008 source.n959 source.n958 9.3005
R1009 source.n957 source.n956 9.3005
R1010 source.n896 source.n895 9.3005
R1011 source.n951 source.n950 9.3005
R1012 source.n949 source.n948 9.3005
R1013 source.n900 source.n899 9.3005
R1014 source.n943 source.n942 9.3005
R1015 source.n941 source.n940 9.3005
R1016 source.n917 source.n916 9.3005
R1017 source.n912 source.n911 9.3005
R1018 source.n923 source.n922 9.3005
R1019 source.n925 source.n924 9.3005
R1020 source.n908 source.n907 9.3005
R1021 source.n931 source.n930 9.3005
R1022 source.n933 source.n932 9.3005
R1023 source.n934 source.n903 9.3005
R1024 source.n892 source.n891 9.3005
R1025 source.n965 source.n964 9.3005
R1026 source.n967 source.n966 9.3005
R1027 source.n888 source.n887 9.3005
R1028 source.n973 source.n972 9.3005
R1029 source.n975 source.n974 9.3005
R1030 source.n884 source.n883 9.3005
R1031 source.n982 source.n981 9.3005
R1032 source.n984 source.n983 9.3005
R1033 source.n1007 source.n1006 9.3005
R1034 source.n732 source.n731 9.3005
R1035 source.n861 source.n860 9.3005
R1036 source.n859 source.n858 9.3005
R1037 source.n736 source.n735 9.3005
R1038 source.n853 source.n852 9.3005
R1039 source.n851 source.n850 9.3005
R1040 source.n740 source.n739 9.3005
R1041 source.n819 source.n818 9.3005
R1042 source.n817 source.n816 9.3005
R1043 source.n756 source.n755 9.3005
R1044 source.n811 source.n810 9.3005
R1045 source.n809 source.n808 9.3005
R1046 source.n760 source.n759 9.3005
R1047 source.n803 source.n802 9.3005
R1048 source.n801 source.n800 9.3005
R1049 source.n777 source.n776 9.3005
R1050 source.n772 source.n771 9.3005
R1051 source.n783 source.n782 9.3005
R1052 source.n785 source.n784 9.3005
R1053 source.n768 source.n767 9.3005
R1054 source.n791 source.n790 9.3005
R1055 source.n793 source.n792 9.3005
R1056 source.n794 source.n763 9.3005
R1057 source.n752 source.n751 9.3005
R1058 source.n825 source.n824 9.3005
R1059 source.n827 source.n826 9.3005
R1060 source.n748 source.n747 9.3005
R1061 source.n833 source.n832 9.3005
R1062 source.n835 source.n834 9.3005
R1063 source.n744 source.n743 9.3005
R1064 source.n842 source.n841 9.3005
R1065 source.n844 source.n843 9.3005
R1066 source.n867 source.n866 9.3005
R1067 source.n582 source.n581 9.3005
R1068 source.n711 source.n710 9.3005
R1069 source.n709 source.n708 9.3005
R1070 source.n586 source.n585 9.3005
R1071 source.n703 source.n702 9.3005
R1072 source.n701 source.n700 9.3005
R1073 source.n590 source.n589 9.3005
R1074 source.n669 source.n668 9.3005
R1075 source.n667 source.n666 9.3005
R1076 source.n606 source.n605 9.3005
R1077 source.n661 source.n660 9.3005
R1078 source.n659 source.n658 9.3005
R1079 source.n610 source.n609 9.3005
R1080 source.n653 source.n652 9.3005
R1081 source.n651 source.n650 9.3005
R1082 source.n627 source.n626 9.3005
R1083 source.n622 source.n621 9.3005
R1084 source.n633 source.n632 9.3005
R1085 source.n635 source.n634 9.3005
R1086 source.n618 source.n617 9.3005
R1087 source.n641 source.n640 9.3005
R1088 source.n643 source.n642 9.3005
R1089 source.n644 source.n613 9.3005
R1090 source.n602 source.n601 9.3005
R1091 source.n675 source.n674 9.3005
R1092 source.n677 source.n676 9.3005
R1093 source.n598 source.n597 9.3005
R1094 source.n683 source.n682 9.3005
R1095 source.n685 source.n684 9.3005
R1096 source.n594 source.n593 9.3005
R1097 source.n692 source.n691 9.3005
R1098 source.n694 source.n693 9.3005
R1099 source.n717 source.n716 9.3005
R1100 source.n49 source.n48 9.3005
R1101 source.n44 source.n43 9.3005
R1102 source.n55 source.n54 9.3005
R1103 source.n57 source.n56 9.3005
R1104 source.n40 source.n39 9.3005
R1105 source.n63 source.n62 9.3005
R1106 source.n65 source.n64 9.3005
R1107 source.n37 source.n34 9.3005
R1108 source.n96 source.n95 9.3005
R1109 source.n98 source.n97 9.3005
R1110 source.n19 source.n18 9.3005
R1111 source.n104 source.n103 9.3005
R1112 source.n106 source.n105 9.3005
R1113 source.n14 source.n13 9.3005
R1114 source.n112 source.n111 9.3005
R1115 source.n114 source.n113 9.3005
R1116 source.n137 source.n136 9.3005
R1117 source.n2 source.n1 9.3005
R1118 source.n131 source.n130 9.3005
R1119 source.n129 source.n128 9.3005
R1120 source.n6 source.n5 9.3005
R1121 source.n123 source.n122 9.3005
R1122 source.n121 source.n120 9.3005
R1123 source.n10 source.n9 9.3005
R1124 source.n23 source.n22 9.3005
R1125 source.n90 source.n89 9.3005
R1126 source.n88 source.n87 9.3005
R1127 source.n27 source.n26 9.3005
R1128 source.n82 source.n81 9.3005
R1129 source.n80 source.n79 9.3005
R1130 source.n31 source.n30 9.3005
R1131 source.n74 source.n73 9.3005
R1132 source.n72 source.n71 9.3005
R1133 source.n199 source.n198 9.3005
R1134 source.n194 source.n193 9.3005
R1135 source.n205 source.n204 9.3005
R1136 source.n207 source.n206 9.3005
R1137 source.n190 source.n189 9.3005
R1138 source.n213 source.n212 9.3005
R1139 source.n215 source.n214 9.3005
R1140 source.n187 source.n184 9.3005
R1141 source.n246 source.n245 9.3005
R1142 source.n248 source.n247 9.3005
R1143 source.n169 source.n168 9.3005
R1144 source.n254 source.n253 9.3005
R1145 source.n256 source.n255 9.3005
R1146 source.n164 source.n163 9.3005
R1147 source.n262 source.n261 9.3005
R1148 source.n264 source.n263 9.3005
R1149 source.n287 source.n286 9.3005
R1150 source.n152 source.n151 9.3005
R1151 source.n281 source.n280 9.3005
R1152 source.n279 source.n278 9.3005
R1153 source.n156 source.n155 9.3005
R1154 source.n273 source.n272 9.3005
R1155 source.n271 source.n270 9.3005
R1156 source.n160 source.n159 9.3005
R1157 source.n173 source.n172 9.3005
R1158 source.n240 source.n239 9.3005
R1159 source.n238 source.n237 9.3005
R1160 source.n177 source.n176 9.3005
R1161 source.n232 source.n231 9.3005
R1162 source.n230 source.n229 9.3005
R1163 source.n181 source.n180 9.3005
R1164 source.n224 source.n223 9.3005
R1165 source.n222 source.n221 9.3005
R1166 source.n339 source.n338 9.3005
R1167 source.n334 source.n333 9.3005
R1168 source.n345 source.n344 9.3005
R1169 source.n347 source.n346 9.3005
R1170 source.n330 source.n329 9.3005
R1171 source.n353 source.n352 9.3005
R1172 source.n355 source.n354 9.3005
R1173 source.n327 source.n324 9.3005
R1174 source.n386 source.n385 9.3005
R1175 source.n388 source.n387 9.3005
R1176 source.n309 source.n308 9.3005
R1177 source.n394 source.n393 9.3005
R1178 source.n396 source.n395 9.3005
R1179 source.n304 source.n303 9.3005
R1180 source.n402 source.n401 9.3005
R1181 source.n404 source.n403 9.3005
R1182 source.n427 source.n426 9.3005
R1183 source.n292 source.n291 9.3005
R1184 source.n421 source.n420 9.3005
R1185 source.n419 source.n418 9.3005
R1186 source.n296 source.n295 9.3005
R1187 source.n413 source.n412 9.3005
R1188 source.n411 source.n410 9.3005
R1189 source.n300 source.n299 9.3005
R1190 source.n313 source.n312 9.3005
R1191 source.n380 source.n379 9.3005
R1192 source.n378 source.n377 9.3005
R1193 source.n317 source.n316 9.3005
R1194 source.n372 source.n371 9.3005
R1195 source.n370 source.n369 9.3005
R1196 source.n321 source.n320 9.3005
R1197 source.n364 source.n363 9.3005
R1198 source.n362 source.n361 9.3005
R1199 source.n489 source.n488 9.3005
R1200 source.n484 source.n483 9.3005
R1201 source.n495 source.n494 9.3005
R1202 source.n497 source.n496 9.3005
R1203 source.n480 source.n479 9.3005
R1204 source.n503 source.n502 9.3005
R1205 source.n505 source.n504 9.3005
R1206 source.n477 source.n474 9.3005
R1207 source.n536 source.n535 9.3005
R1208 source.n538 source.n537 9.3005
R1209 source.n459 source.n458 9.3005
R1210 source.n544 source.n543 9.3005
R1211 source.n546 source.n545 9.3005
R1212 source.n454 source.n453 9.3005
R1213 source.n552 source.n551 9.3005
R1214 source.n554 source.n553 9.3005
R1215 source.n577 source.n576 9.3005
R1216 source.n442 source.n441 9.3005
R1217 source.n571 source.n570 9.3005
R1218 source.n569 source.n568 9.3005
R1219 source.n446 source.n445 9.3005
R1220 source.n563 source.n562 9.3005
R1221 source.n561 source.n560 9.3005
R1222 source.n450 source.n449 9.3005
R1223 source.n463 source.n462 9.3005
R1224 source.n530 source.n529 9.3005
R1225 source.n528 source.n527 9.3005
R1226 source.n467 source.n466 9.3005
R1227 source.n522 source.n521 9.3005
R1228 source.n520 source.n519 9.3005
R1229 source.n471 source.n470 9.3005
R1230 source.n514 source.n513 9.3005
R1231 source.n512 source.n511 9.3005
R1232 source.n1072 source.n1071 8.92171
R1233 source.n1105 source.n1046 8.92171
R1234 source.n1118 source.n1038 8.92171
R1235 source.n1152 source.n1151 8.92171
R1236 source.n922 source.n921 8.92171
R1237 source.n955 source.n896 8.92171
R1238 source.n968 source.n888 8.92171
R1239 source.n1002 source.n1001 8.92171
R1240 source.n782 source.n781 8.92171
R1241 source.n815 source.n756 8.92171
R1242 source.n828 source.n748 8.92171
R1243 source.n862 source.n861 8.92171
R1244 source.n632 source.n631 8.92171
R1245 source.n665 source.n606 8.92171
R1246 source.n678 source.n598 8.92171
R1247 source.n712 source.n711 8.92171
R1248 source.n132 source.n131 8.92171
R1249 source.n99 source.n19 8.92171
R1250 source.n86 source.n27 8.92171
R1251 source.n54 source.n53 8.92171
R1252 source.n282 source.n281 8.92171
R1253 source.n249 source.n169 8.92171
R1254 source.n236 source.n177 8.92171
R1255 source.n204 source.n203 8.92171
R1256 source.n422 source.n421 8.92171
R1257 source.n389 source.n309 8.92171
R1258 source.n376 source.n317 8.92171
R1259 source.n344 source.n343 8.92171
R1260 source.n572 source.n571 8.92171
R1261 source.n539 source.n459 8.92171
R1262 source.n526 source.n467 8.92171
R1263 source.n494 source.n493 8.92171
R1264 source.n1068 source.n1062 8.14595
R1265 source.n1106 source.n1044 8.14595
R1266 source.n1117 source.n1040 8.14595
R1267 source.n1155 source.n1022 8.14595
R1268 source.n918 source.n912 8.14595
R1269 source.n956 source.n894 8.14595
R1270 source.n967 source.n890 8.14595
R1271 source.n1005 source.n872 8.14595
R1272 source.n778 source.n772 8.14595
R1273 source.n816 source.n754 8.14595
R1274 source.n827 source.n750 8.14595
R1275 source.n865 source.n732 8.14595
R1276 source.n628 source.n622 8.14595
R1277 source.n666 source.n604 8.14595
R1278 source.n677 source.n600 8.14595
R1279 source.n715 source.n582 8.14595
R1280 source.n135 source.n2 8.14595
R1281 source.n98 source.n21 8.14595
R1282 source.n87 source.n25 8.14595
R1283 source.n50 source.n44 8.14595
R1284 source.n285 source.n152 8.14595
R1285 source.n248 source.n171 8.14595
R1286 source.n237 source.n175 8.14595
R1287 source.n200 source.n194 8.14595
R1288 source.n425 source.n292 8.14595
R1289 source.n388 source.n311 8.14595
R1290 source.n377 source.n315 8.14595
R1291 source.n340 source.n334 8.14595
R1292 source.n575 source.n442 8.14595
R1293 source.n538 source.n461 8.14595
R1294 source.n527 source.n465 8.14595
R1295 source.n490 source.n484 8.14595
R1296 source.n1067 source.n1064 7.3702
R1297 source.n1110 source.n1109 7.3702
R1298 source.n1114 source.n1113 7.3702
R1299 source.n1156 source.n1020 7.3702
R1300 source.n917 source.n914 7.3702
R1301 source.n960 source.n959 7.3702
R1302 source.n964 source.n963 7.3702
R1303 source.n1006 source.n870 7.3702
R1304 source.n777 source.n774 7.3702
R1305 source.n820 source.n819 7.3702
R1306 source.n824 source.n823 7.3702
R1307 source.n866 source.n730 7.3702
R1308 source.n627 source.n624 7.3702
R1309 source.n670 source.n669 7.3702
R1310 source.n674 source.n673 7.3702
R1311 source.n716 source.n580 7.3702
R1312 source.n136 source.n0 7.3702
R1313 source.n95 source.n94 7.3702
R1314 source.n91 source.n90 7.3702
R1315 source.n49 source.n46 7.3702
R1316 source.n286 source.n150 7.3702
R1317 source.n245 source.n244 7.3702
R1318 source.n241 source.n240 7.3702
R1319 source.n199 source.n196 7.3702
R1320 source.n426 source.n290 7.3702
R1321 source.n385 source.n384 7.3702
R1322 source.n381 source.n380 7.3702
R1323 source.n339 source.n336 7.3702
R1324 source.n576 source.n440 7.3702
R1325 source.n535 source.n534 7.3702
R1326 source.n531 source.n530 7.3702
R1327 source.n489 source.n486 7.3702
R1328 source.n1110 source.n1042 6.59444
R1329 source.n1113 source.n1042 6.59444
R1330 source.n1158 source.n1020 6.59444
R1331 source.n960 source.n892 6.59444
R1332 source.n963 source.n892 6.59444
R1333 source.n1008 source.n870 6.59444
R1334 source.n820 source.n752 6.59444
R1335 source.n823 source.n752 6.59444
R1336 source.n868 source.n730 6.59444
R1337 source.n670 source.n602 6.59444
R1338 source.n673 source.n602 6.59444
R1339 source.n718 source.n580 6.59444
R1340 source.n138 source.n0 6.59444
R1341 source.n94 source.n23 6.59444
R1342 source.n91 source.n23 6.59444
R1343 source.n288 source.n150 6.59444
R1344 source.n244 source.n173 6.59444
R1345 source.n241 source.n173 6.59444
R1346 source.n428 source.n290 6.59444
R1347 source.n384 source.n313 6.59444
R1348 source.n381 source.n313 6.59444
R1349 source.n578 source.n440 6.59444
R1350 source.n534 source.n463 6.59444
R1351 source.n531 source.n463 6.59444
R1352 source.n1068 source.n1067 5.81868
R1353 source.n1109 source.n1044 5.81868
R1354 source.n1114 source.n1040 5.81868
R1355 source.n1156 source.n1155 5.81868
R1356 source.n918 source.n917 5.81868
R1357 source.n959 source.n894 5.81868
R1358 source.n964 source.n890 5.81868
R1359 source.n1006 source.n1005 5.81868
R1360 source.n778 source.n777 5.81868
R1361 source.n819 source.n754 5.81868
R1362 source.n824 source.n750 5.81868
R1363 source.n866 source.n865 5.81868
R1364 source.n628 source.n627 5.81868
R1365 source.n669 source.n604 5.81868
R1366 source.n674 source.n600 5.81868
R1367 source.n716 source.n715 5.81868
R1368 source.n136 source.n135 5.81868
R1369 source.n95 source.n21 5.81868
R1370 source.n90 source.n25 5.81868
R1371 source.n50 source.n49 5.81868
R1372 source.n286 source.n285 5.81868
R1373 source.n245 source.n171 5.81868
R1374 source.n240 source.n175 5.81868
R1375 source.n200 source.n199 5.81868
R1376 source.n426 source.n425 5.81868
R1377 source.n385 source.n311 5.81868
R1378 source.n380 source.n315 5.81868
R1379 source.n340 source.n339 5.81868
R1380 source.n576 source.n575 5.81868
R1381 source.n535 source.n461 5.81868
R1382 source.n530 source.n465 5.81868
R1383 source.n490 source.n489 5.81868
R1384 source.n1160 source.n1159 5.53498
R1385 source.n1071 source.n1062 5.04292
R1386 source.n1106 source.n1105 5.04292
R1387 source.n1118 source.n1117 5.04292
R1388 source.n1152 source.n1022 5.04292
R1389 source.n921 source.n912 5.04292
R1390 source.n956 source.n955 5.04292
R1391 source.n968 source.n967 5.04292
R1392 source.n1002 source.n872 5.04292
R1393 source.n781 source.n772 5.04292
R1394 source.n816 source.n815 5.04292
R1395 source.n828 source.n827 5.04292
R1396 source.n862 source.n732 5.04292
R1397 source.n631 source.n622 5.04292
R1398 source.n666 source.n665 5.04292
R1399 source.n678 source.n677 5.04292
R1400 source.n712 source.n582 5.04292
R1401 source.n132 source.n2 5.04292
R1402 source.n99 source.n98 5.04292
R1403 source.n87 source.n86 5.04292
R1404 source.n53 source.n44 5.04292
R1405 source.n282 source.n152 5.04292
R1406 source.n249 source.n248 5.04292
R1407 source.n237 source.n236 5.04292
R1408 source.n203 source.n194 5.04292
R1409 source.n422 source.n292 5.04292
R1410 source.n389 source.n388 5.04292
R1411 source.n377 source.n376 5.04292
R1412 source.n343 source.n334 5.04292
R1413 source.n572 source.n442 5.04292
R1414 source.n539 source.n538 5.04292
R1415 source.n527 source.n526 5.04292
R1416 source.n493 source.n484 5.04292
R1417 source.n1072 source.n1060 4.26717
R1418 source.n1102 source.n1046 4.26717
R1419 source.n1121 source.n1038 4.26717
R1420 source.n1151 source.n1024 4.26717
R1421 source.n922 source.n910 4.26717
R1422 source.n952 source.n896 4.26717
R1423 source.n971 source.n888 4.26717
R1424 source.n1001 source.n874 4.26717
R1425 source.n782 source.n770 4.26717
R1426 source.n812 source.n756 4.26717
R1427 source.n831 source.n748 4.26717
R1428 source.n861 source.n734 4.26717
R1429 source.n632 source.n620 4.26717
R1430 source.n662 source.n606 4.26717
R1431 source.n681 source.n598 4.26717
R1432 source.n711 source.n584 4.26717
R1433 source.n131 source.n4 4.26717
R1434 source.n102 source.n19 4.26717
R1435 source.n83 source.n27 4.26717
R1436 source.n54 source.n42 4.26717
R1437 source.n281 source.n154 4.26717
R1438 source.n252 source.n169 4.26717
R1439 source.n233 source.n177 4.26717
R1440 source.n204 source.n192 4.26717
R1441 source.n421 source.n294 4.26717
R1442 source.n392 source.n309 4.26717
R1443 source.n373 source.n317 4.26717
R1444 source.n344 source.n332 4.26717
R1445 source.n571 source.n444 4.26717
R1446 source.n542 source.n459 4.26717
R1447 source.n523 source.n467 4.26717
R1448 source.n494 source.n482 4.26717
R1449 source.n1076 source.n1075 3.49141
R1450 source.n1101 source.n1048 3.49141
R1451 source.n1122 source.n1036 3.49141
R1452 source.n1148 source.n1147 3.49141
R1453 source.n926 source.n925 3.49141
R1454 source.n951 source.n898 3.49141
R1455 source.n972 source.n886 3.49141
R1456 source.n998 source.n997 3.49141
R1457 source.n786 source.n785 3.49141
R1458 source.n811 source.n758 3.49141
R1459 source.n832 source.n746 3.49141
R1460 source.n858 source.n857 3.49141
R1461 source.n636 source.n635 3.49141
R1462 source.n661 source.n608 3.49141
R1463 source.n682 source.n596 3.49141
R1464 source.n708 source.n707 3.49141
R1465 source.n128 source.n127 3.49141
R1466 source.n103 source.n17 3.49141
R1467 source.n82 source.n29 3.49141
R1468 source.n58 source.n57 3.49141
R1469 source.n278 source.n277 3.49141
R1470 source.n253 source.n167 3.49141
R1471 source.n232 source.n179 3.49141
R1472 source.n208 source.n207 3.49141
R1473 source.n418 source.n417 3.49141
R1474 source.n393 source.n307 3.49141
R1475 source.n372 source.n319 3.49141
R1476 source.n348 source.n347 3.49141
R1477 source.n568 source.n567 3.49141
R1478 source.n543 source.n457 3.49141
R1479 source.n522 source.n469 3.49141
R1480 source.n498 source.n497 3.49141
R1481 source.n48 source.n47 2.84303
R1482 source.n198 source.n197 2.84303
R1483 source.n338 source.n337 2.84303
R1484 source.n488 source.n487 2.84303
R1485 source.n1066 source.n1065 2.84303
R1486 source.n916 source.n915 2.84303
R1487 source.n776 source.n775 2.84303
R1488 source.n626 source.n625 2.84303
R1489 source.n1079 source.n1058 2.71565
R1490 source.n1098 source.n1097 2.71565
R1491 source.n1126 source.n1125 2.71565
R1492 source.n1144 source.n1026 2.71565
R1493 source.n929 source.n908 2.71565
R1494 source.n948 source.n947 2.71565
R1495 source.n976 source.n975 2.71565
R1496 source.n994 source.n876 2.71565
R1497 source.n789 source.n768 2.71565
R1498 source.n808 source.n807 2.71565
R1499 source.n836 source.n835 2.71565
R1500 source.n854 source.n736 2.71565
R1501 source.n639 source.n618 2.71565
R1502 source.n658 source.n657 2.71565
R1503 source.n686 source.n685 2.71565
R1504 source.n704 source.n586 2.71565
R1505 source.n124 source.n6 2.71565
R1506 source.n107 source.n106 2.71565
R1507 source.n79 source.n78 2.71565
R1508 source.n61 source.n40 2.71565
R1509 source.n274 source.n156 2.71565
R1510 source.n257 source.n256 2.71565
R1511 source.n229 source.n228 2.71565
R1512 source.n211 source.n190 2.71565
R1513 source.n414 source.n296 2.71565
R1514 source.n397 source.n396 2.71565
R1515 source.n369 source.n368 2.71565
R1516 source.n351 source.n330 2.71565
R1517 source.n564 source.n446 2.71565
R1518 source.n547 source.n546 2.71565
R1519 source.n519 source.n518 2.71565
R1520 source.n501 source.n480 2.71565
R1521 source.n1080 source.n1056 1.93989
R1522 source.n1094 source.n1050 1.93989
R1523 source.n1130 source.n1034 1.93989
R1524 source.n1143 source.n1028 1.93989
R1525 source.n930 source.n906 1.93989
R1526 source.n944 source.n900 1.93989
R1527 source.n980 source.n884 1.93989
R1528 source.n993 source.n878 1.93989
R1529 source.n790 source.n766 1.93989
R1530 source.n804 source.n760 1.93989
R1531 source.n840 source.n744 1.93989
R1532 source.n853 source.n738 1.93989
R1533 source.n640 source.n616 1.93989
R1534 source.n654 source.n610 1.93989
R1535 source.n690 source.n594 1.93989
R1536 source.n703 source.n588 1.93989
R1537 source.n123 source.n8 1.93989
R1538 source.n110 source.n14 1.93989
R1539 source.n75 source.n31 1.93989
R1540 source.n62 source.n38 1.93989
R1541 source.n273 source.n158 1.93989
R1542 source.n260 source.n164 1.93989
R1543 source.n225 source.n181 1.93989
R1544 source.n212 source.n188 1.93989
R1545 source.n413 source.n298 1.93989
R1546 source.n400 source.n304 1.93989
R1547 source.n365 source.n321 1.93989
R1548 source.n352 source.n328 1.93989
R1549 source.n563 source.n448 1.93989
R1550 source.n550 source.n454 1.93989
R1551 source.n515 source.n471 1.93989
R1552 source.n502 source.n478 1.93989
R1553 source.n1085 source.n1083 1.16414
R1554 source.n1093 source.n1052 1.16414
R1555 source.n1131 source.n1032 1.16414
R1556 source.n1140 source.n1139 1.16414
R1557 source.n935 source.n933 1.16414
R1558 source.n943 source.n902 1.16414
R1559 source.n981 source.n882 1.16414
R1560 source.n990 source.n989 1.16414
R1561 source.n795 source.n793 1.16414
R1562 source.n803 source.n762 1.16414
R1563 source.n841 source.n742 1.16414
R1564 source.n850 source.n849 1.16414
R1565 source.n645 source.n643 1.16414
R1566 source.n653 source.n612 1.16414
R1567 source.n691 source.n592 1.16414
R1568 source.n700 source.n699 1.16414
R1569 source.n120 source.n119 1.16414
R1570 source.n111 source.n12 1.16414
R1571 source.n74 source.n33 1.16414
R1572 source.n66 source.n65 1.16414
R1573 source.n270 source.n269 1.16414
R1574 source.n261 source.n162 1.16414
R1575 source.n224 source.n183 1.16414
R1576 source.n216 source.n215 1.16414
R1577 source.n410 source.n409 1.16414
R1578 source.n401 source.n302 1.16414
R1579 source.n364 source.n323 1.16414
R1580 source.n356 source.n355 1.16414
R1581 source.n560 source.n559 1.16414
R1582 source.n551 source.n452 1.16414
R1583 source.n514 source.n473 1.16414
R1584 source.n506 source.n505 1.16414
R1585 source.n1018 source.t19 0.7925
R1586 source.n1018 source.t21 0.7925
R1587 source.n1016 source.t18 0.7925
R1588 source.n1016 source.t3 0.7925
R1589 source.n1014 source.t4 0.7925
R1590 source.n1014 source.t7 0.7925
R1591 source.n1012 source.t9 0.7925
R1592 source.n1012 source.t12 0.7925
R1593 source.n1010 source.t11 0.7925
R1594 source.n1010 source.t14 0.7925
R1595 source.n728 source.t24 0.7925
R1596 source.n728 source.t36 0.7925
R1597 source.n726 source.t41 0.7925
R1598 source.n726 source.t33 0.7925
R1599 source.n724 source.t40 0.7925
R1600 source.n724 source.t31 0.7925
R1601 source.n722 source.t43 0.7925
R1602 source.n722 source.t29 0.7925
R1603 source.n720 source.t35 0.7925
R1604 source.n720 source.t28 0.7925
R1605 source.n140 source.t30 0.7925
R1606 source.n140 source.t47 0.7925
R1607 source.n142 source.t46 0.7925
R1608 source.n142 source.t37 0.7925
R1609 source.n144 source.t34 0.7925
R1610 source.n144 source.t27 0.7925
R1611 source.n146 source.t26 0.7925
R1612 source.n146 source.t39 0.7925
R1613 source.n148 source.t38 0.7925
R1614 source.n148 source.t32 0.7925
R1615 source.n430 source.t0 0.7925
R1616 source.n430 source.t17 0.7925
R1617 source.n432 source.t1 0.7925
R1618 source.n432 source.t16 0.7925
R1619 source.n434 source.t13 0.7925
R1620 source.n434 source.t6 0.7925
R1621 source.n436 source.t20 0.7925
R1622 source.n436 source.t22 0.7925
R1623 source.n438 source.t5 0.7925
R1624 source.n438 source.t15 0.7925
R1625 source.n579 source.n439 0.543603
R1626 source.n439 source.n437 0.543603
R1627 source.n437 source.n435 0.543603
R1628 source.n435 source.n433 0.543603
R1629 source.n433 source.n431 0.543603
R1630 source.n431 source.n429 0.543603
R1631 source.n289 source.n149 0.543603
R1632 source.n149 source.n147 0.543603
R1633 source.n147 source.n145 0.543603
R1634 source.n145 source.n143 0.543603
R1635 source.n143 source.n141 0.543603
R1636 source.n141 source.n139 0.543603
R1637 source.n721 source.n719 0.543603
R1638 source.n723 source.n721 0.543603
R1639 source.n725 source.n723 0.543603
R1640 source.n727 source.n725 0.543603
R1641 source.n729 source.n727 0.543603
R1642 source.n869 source.n729 0.543603
R1643 source.n1011 source.n1009 0.543603
R1644 source.n1013 source.n1011 0.543603
R1645 source.n1015 source.n1013 0.543603
R1646 source.n1017 source.n1015 0.543603
R1647 source.n1019 source.n1017 0.543603
R1648 source.n1159 source.n1019 0.543603
R1649 source.n429 source.n289 0.470328
R1650 source.n1009 source.n869 0.470328
R1651 source.n1084 source.n1054 0.388379
R1652 source.n1090 source.n1089 0.388379
R1653 source.n1135 source.n1134 0.388379
R1654 source.n1136 source.n1030 0.388379
R1655 source.n934 source.n904 0.388379
R1656 source.n940 source.n939 0.388379
R1657 source.n985 source.n984 0.388379
R1658 source.n986 source.n880 0.388379
R1659 source.n794 source.n764 0.388379
R1660 source.n800 source.n799 0.388379
R1661 source.n845 source.n844 0.388379
R1662 source.n846 source.n740 0.388379
R1663 source.n644 source.n614 0.388379
R1664 source.n650 source.n649 0.388379
R1665 source.n695 source.n694 0.388379
R1666 source.n696 source.n590 0.388379
R1667 source.n116 source.n10 0.388379
R1668 source.n115 source.n114 0.388379
R1669 source.n71 source.n70 0.388379
R1670 source.n37 source.n35 0.388379
R1671 source.n266 source.n160 0.388379
R1672 source.n265 source.n264 0.388379
R1673 source.n221 source.n220 0.388379
R1674 source.n187 source.n185 0.388379
R1675 source.n406 source.n300 0.388379
R1676 source.n405 source.n404 0.388379
R1677 source.n361 source.n360 0.388379
R1678 source.n327 source.n325 0.388379
R1679 source.n556 source.n450 0.388379
R1680 source.n555 source.n554 0.388379
R1681 source.n511 source.n510 0.388379
R1682 source.n477 source.n475 0.388379
R1683 source source.n1160 0.188
R1684 source.n1066 source.n1061 0.155672
R1685 source.n1073 source.n1061 0.155672
R1686 source.n1074 source.n1073 0.155672
R1687 source.n1074 source.n1057 0.155672
R1688 source.n1081 source.n1057 0.155672
R1689 source.n1082 source.n1081 0.155672
R1690 source.n1082 source.n1053 0.155672
R1691 source.n1091 source.n1053 0.155672
R1692 source.n1092 source.n1091 0.155672
R1693 source.n1092 source.n1049 0.155672
R1694 source.n1099 source.n1049 0.155672
R1695 source.n1100 source.n1099 0.155672
R1696 source.n1100 source.n1045 0.155672
R1697 source.n1107 source.n1045 0.155672
R1698 source.n1108 source.n1107 0.155672
R1699 source.n1108 source.n1041 0.155672
R1700 source.n1115 source.n1041 0.155672
R1701 source.n1116 source.n1115 0.155672
R1702 source.n1116 source.n1037 0.155672
R1703 source.n1123 source.n1037 0.155672
R1704 source.n1124 source.n1123 0.155672
R1705 source.n1124 source.n1033 0.155672
R1706 source.n1132 source.n1033 0.155672
R1707 source.n1133 source.n1132 0.155672
R1708 source.n1133 source.n1029 0.155672
R1709 source.n1141 source.n1029 0.155672
R1710 source.n1142 source.n1141 0.155672
R1711 source.n1142 source.n1025 0.155672
R1712 source.n1149 source.n1025 0.155672
R1713 source.n1150 source.n1149 0.155672
R1714 source.n1150 source.n1021 0.155672
R1715 source.n1157 source.n1021 0.155672
R1716 source.n916 source.n911 0.155672
R1717 source.n923 source.n911 0.155672
R1718 source.n924 source.n923 0.155672
R1719 source.n924 source.n907 0.155672
R1720 source.n931 source.n907 0.155672
R1721 source.n932 source.n931 0.155672
R1722 source.n932 source.n903 0.155672
R1723 source.n941 source.n903 0.155672
R1724 source.n942 source.n941 0.155672
R1725 source.n942 source.n899 0.155672
R1726 source.n949 source.n899 0.155672
R1727 source.n950 source.n949 0.155672
R1728 source.n950 source.n895 0.155672
R1729 source.n957 source.n895 0.155672
R1730 source.n958 source.n957 0.155672
R1731 source.n958 source.n891 0.155672
R1732 source.n965 source.n891 0.155672
R1733 source.n966 source.n965 0.155672
R1734 source.n966 source.n887 0.155672
R1735 source.n973 source.n887 0.155672
R1736 source.n974 source.n973 0.155672
R1737 source.n974 source.n883 0.155672
R1738 source.n982 source.n883 0.155672
R1739 source.n983 source.n982 0.155672
R1740 source.n983 source.n879 0.155672
R1741 source.n991 source.n879 0.155672
R1742 source.n992 source.n991 0.155672
R1743 source.n992 source.n875 0.155672
R1744 source.n999 source.n875 0.155672
R1745 source.n1000 source.n999 0.155672
R1746 source.n1000 source.n871 0.155672
R1747 source.n1007 source.n871 0.155672
R1748 source.n776 source.n771 0.155672
R1749 source.n783 source.n771 0.155672
R1750 source.n784 source.n783 0.155672
R1751 source.n784 source.n767 0.155672
R1752 source.n791 source.n767 0.155672
R1753 source.n792 source.n791 0.155672
R1754 source.n792 source.n763 0.155672
R1755 source.n801 source.n763 0.155672
R1756 source.n802 source.n801 0.155672
R1757 source.n802 source.n759 0.155672
R1758 source.n809 source.n759 0.155672
R1759 source.n810 source.n809 0.155672
R1760 source.n810 source.n755 0.155672
R1761 source.n817 source.n755 0.155672
R1762 source.n818 source.n817 0.155672
R1763 source.n818 source.n751 0.155672
R1764 source.n825 source.n751 0.155672
R1765 source.n826 source.n825 0.155672
R1766 source.n826 source.n747 0.155672
R1767 source.n833 source.n747 0.155672
R1768 source.n834 source.n833 0.155672
R1769 source.n834 source.n743 0.155672
R1770 source.n842 source.n743 0.155672
R1771 source.n843 source.n842 0.155672
R1772 source.n843 source.n739 0.155672
R1773 source.n851 source.n739 0.155672
R1774 source.n852 source.n851 0.155672
R1775 source.n852 source.n735 0.155672
R1776 source.n859 source.n735 0.155672
R1777 source.n860 source.n859 0.155672
R1778 source.n860 source.n731 0.155672
R1779 source.n867 source.n731 0.155672
R1780 source.n626 source.n621 0.155672
R1781 source.n633 source.n621 0.155672
R1782 source.n634 source.n633 0.155672
R1783 source.n634 source.n617 0.155672
R1784 source.n641 source.n617 0.155672
R1785 source.n642 source.n641 0.155672
R1786 source.n642 source.n613 0.155672
R1787 source.n651 source.n613 0.155672
R1788 source.n652 source.n651 0.155672
R1789 source.n652 source.n609 0.155672
R1790 source.n659 source.n609 0.155672
R1791 source.n660 source.n659 0.155672
R1792 source.n660 source.n605 0.155672
R1793 source.n667 source.n605 0.155672
R1794 source.n668 source.n667 0.155672
R1795 source.n668 source.n601 0.155672
R1796 source.n675 source.n601 0.155672
R1797 source.n676 source.n675 0.155672
R1798 source.n676 source.n597 0.155672
R1799 source.n683 source.n597 0.155672
R1800 source.n684 source.n683 0.155672
R1801 source.n684 source.n593 0.155672
R1802 source.n692 source.n593 0.155672
R1803 source.n693 source.n692 0.155672
R1804 source.n693 source.n589 0.155672
R1805 source.n701 source.n589 0.155672
R1806 source.n702 source.n701 0.155672
R1807 source.n702 source.n585 0.155672
R1808 source.n709 source.n585 0.155672
R1809 source.n710 source.n709 0.155672
R1810 source.n710 source.n581 0.155672
R1811 source.n717 source.n581 0.155672
R1812 source.n137 source.n1 0.155672
R1813 source.n130 source.n1 0.155672
R1814 source.n130 source.n129 0.155672
R1815 source.n129 source.n5 0.155672
R1816 source.n122 source.n5 0.155672
R1817 source.n122 source.n121 0.155672
R1818 source.n121 source.n9 0.155672
R1819 source.n113 source.n9 0.155672
R1820 source.n113 source.n112 0.155672
R1821 source.n112 source.n13 0.155672
R1822 source.n105 source.n13 0.155672
R1823 source.n105 source.n104 0.155672
R1824 source.n104 source.n18 0.155672
R1825 source.n97 source.n18 0.155672
R1826 source.n97 source.n96 0.155672
R1827 source.n96 source.n22 0.155672
R1828 source.n89 source.n22 0.155672
R1829 source.n89 source.n88 0.155672
R1830 source.n88 source.n26 0.155672
R1831 source.n81 source.n26 0.155672
R1832 source.n81 source.n80 0.155672
R1833 source.n80 source.n30 0.155672
R1834 source.n73 source.n30 0.155672
R1835 source.n73 source.n72 0.155672
R1836 source.n72 source.n34 0.155672
R1837 source.n64 source.n34 0.155672
R1838 source.n64 source.n63 0.155672
R1839 source.n63 source.n39 0.155672
R1840 source.n56 source.n39 0.155672
R1841 source.n56 source.n55 0.155672
R1842 source.n55 source.n43 0.155672
R1843 source.n48 source.n43 0.155672
R1844 source.n287 source.n151 0.155672
R1845 source.n280 source.n151 0.155672
R1846 source.n280 source.n279 0.155672
R1847 source.n279 source.n155 0.155672
R1848 source.n272 source.n155 0.155672
R1849 source.n272 source.n271 0.155672
R1850 source.n271 source.n159 0.155672
R1851 source.n263 source.n159 0.155672
R1852 source.n263 source.n262 0.155672
R1853 source.n262 source.n163 0.155672
R1854 source.n255 source.n163 0.155672
R1855 source.n255 source.n254 0.155672
R1856 source.n254 source.n168 0.155672
R1857 source.n247 source.n168 0.155672
R1858 source.n247 source.n246 0.155672
R1859 source.n246 source.n172 0.155672
R1860 source.n239 source.n172 0.155672
R1861 source.n239 source.n238 0.155672
R1862 source.n238 source.n176 0.155672
R1863 source.n231 source.n176 0.155672
R1864 source.n231 source.n230 0.155672
R1865 source.n230 source.n180 0.155672
R1866 source.n223 source.n180 0.155672
R1867 source.n223 source.n222 0.155672
R1868 source.n222 source.n184 0.155672
R1869 source.n214 source.n184 0.155672
R1870 source.n214 source.n213 0.155672
R1871 source.n213 source.n189 0.155672
R1872 source.n206 source.n189 0.155672
R1873 source.n206 source.n205 0.155672
R1874 source.n205 source.n193 0.155672
R1875 source.n198 source.n193 0.155672
R1876 source.n427 source.n291 0.155672
R1877 source.n420 source.n291 0.155672
R1878 source.n420 source.n419 0.155672
R1879 source.n419 source.n295 0.155672
R1880 source.n412 source.n295 0.155672
R1881 source.n412 source.n411 0.155672
R1882 source.n411 source.n299 0.155672
R1883 source.n403 source.n299 0.155672
R1884 source.n403 source.n402 0.155672
R1885 source.n402 source.n303 0.155672
R1886 source.n395 source.n303 0.155672
R1887 source.n395 source.n394 0.155672
R1888 source.n394 source.n308 0.155672
R1889 source.n387 source.n308 0.155672
R1890 source.n387 source.n386 0.155672
R1891 source.n386 source.n312 0.155672
R1892 source.n379 source.n312 0.155672
R1893 source.n379 source.n378 0.155672
R1894 source.n378 source.n316 0.155672
R1895 source.n371 source.n316 0.155672
R1896 source.n371 source.n370 0.155672
R1897 source.n370 source.n320 0.155672
R1898 source.n363 source.n320 0.155672
R1899 source.n363 source.n362 0.155672
R1900 source.n362 source.n324 0.155672
R1901 source.n354 source.n324 0.155672
R1902 source.n354 source.n353 0.155672
R1903 source.n353 source.n329 0.155672
R1904 source.n346 source.n329 0.155672
R1905 source.n346 source.n345 0.155672
R1906 source.n345 source.n333 0.155672
R1907 source.n338 source.n333 0.155672
R1908 source.n577 source.n441 0.155672
R1909 source.n570 source.n441 0.155672
R1910 source.n570 source.n569 0.155672
R1911 source.n569 source.n445 0.155672
R1912 source.n562 source.n445 0.155672
R1913 source.n562 source.n561 0.155672
R1914 source.n561 source.n449 0.155672
R1915 source.n553 source.n449 0.155672
R1916 source.n553 source.n552 0.155672
R1917 source.n552 source.n453 0.155672
R1918 source.n545 source.n453 0.155672
R1919 source.n545 source.n544 0.155672
R1920 source.n544 source.n458 0.155672
R1921 source.n537 source.n458 0.155672
R1922 source.n537 source.n536 0.155672
R1923 source.n536 source.n462 0.155672
R1924 source.n529 source.n462 0.155672
R1925 source.n529 source.n528 0.155672
R1926 source.n528 source.n466 0.155672
R1927 source.n521 source.n466 0.155672
R1928 source.n521 source.n520 0.155672
R1929 source.n520 source.n470 0.155672
R1930 source.n513 source.n470 0.155672
R1931 source.n513 source.n512 0.155672
R1932 source.n512 source.n474 0.155672
R1933 source.n504 source.n474 0.155672
R1934 source.n504 source.n503 0.155672
R1935 source.n503 source.n479 0.155672
R1936 source.n496 source.n479 0.155672
R1937 source.n496 source.n495 0.155672
R1938 source.n495 source.n483 0.155672
R1939 source.n488 source.n483 0.155672
R1940 minus.n35 minus.t3 2144.17
R1941 minus.n9 minus.t14 2144.17
R1942 minus.n72 minus.t7 2144.17
R1943 minus.n46 minus.t5 2144.17
R1944 minus.n34 minus.t19 2112.77
R1945 minus.n1 minus.t9 2112.77
R1946 minus.n28 minus.t2 2112.77
R1947 minus.n26 minus.t22 2112.77
R1948 minus.n3 minus.t8 2112.77
R1949 minus.n20 minus.t0 2112.77
R1950 minus.n5 minus.t18 2112.77
R1951 minus.n15 minus.t12 2112.77
R1952 minus.n13 minus.t1 2112.77
R1953 minus.n8 minus.t21 2112.77
R1954 minus.n71 minus.t13 2112.77
R1955 minus.n38 minus.t6 2112.77
R1956 minus.n65 minus.t17 2112.77
R1957 minus.n63 minus.t20 2112.77
R1958 minus.n40 minus.t10 2112.77
R1959 minus.n57 minus.t23 2112.77
R1960 minus.n42 minus.t11 2112.77
R1961 minus.n52 minus.t15 2112.77
R1962 minus.n50 minus.t4 2112.77
R1963 minus.n45 minus.t16 2112.77
R1964 minus.n10 minus.n9 161.489
R1965 minus.n47 minus.n46 161.489
R1966 minus.n36 minus.n35 161.3
R1967 minus.n33 minus.n0 161.3
R1968 minus.n32 minus.n31 161.3
R1969 minus.n30 minus.n29 161.3
R1970 minus.n27 minus.n2 161.3
R1971 minus.n25 minus.n24 161.3
R1972 minus.n23 minus.n22 161.3
R1973 minus.n21 minus.n4 161.3
R1974 minus.n19 minus.n18 161.3
R1975 minus.n17 minus.n16 161.3
R1976 minus.n14 minus.n6 161.3
R1977 minus.n12 minus.n11 161.3
R1978 minus.n10 minus.n7 161.3
R1979 minus.n73 minus.n72 161.3
R1980 minus.n70 minus.n37 161.3
R1981 minus.n69 minus.n68 161.3
R1982 minus.n67 minus.n66 161.3
R1983 minus.n64 minus.n39 161.3
R1984 minus.n62 minus.n61 161.3
R1985 minus.n60 minus.n59 161.3
R1986 minus.n58 minus.n41 161.3
R1987 minus.n56 minus.n55 161.3
R1988 minus.n54 minus.n53 161.3
R1989 minus.n51 minus.n43 161.3
R1990 minus.n49 minus.n48 161.3
R1991 minus.n47 minus.n44 161.3
R1992 minus.n33 minus.n32 73.0308
R1993 minus.n22 minus.n21 73.0308
R1994 minus.n12 minus.n7 73.0308
R1995 minus.n49 minus.n44 73.0308
R1996 minus.n59 minus.n58 73.0308
R1997 minus.n70 minus.n69 73.0308
R1998 minus.n29 minus.n1 66.4581
R1999 minus.n14 minus.n13 66.4581
R2000 minus.n51 minus.n50 66.4581
R2001 minus.n66 minus.n38 66.4581
R2002 minus.n25 minus.n3 63.5369
R2003 minus.n20 minus.n19 63.5369
R2004 minus.n57 minus.n56 63.5369
R2005 minus.n62 minus.n40 63.5369
R2006 minus.n35 minus.n34 60.6157
R2007 minus.n9 minus.n8 60.6157
R2008 minus.n46 minus.n45 60.6157
R2009 minus.n72 minus.n71 60.6157
R2010 minus.n74 minus.n36 47.8566
R2011 minus.n28 minus.n27 47.4702
R2012 minus.n16 minus.n15 47.4702
R2013 minus.n53 minus.n52 47.4702
R2014 minus.n65 minus.n64 47.4702
R2015 minus.n27 minus.n26 44.549
R2016 minus.n16 minus.n5 44.549
R2017 minus.n53 minus.n42 44.549
R2018 minus.n64 minus.n63 44.549
R2019 minus.n26 minus.n25 28.4823
R2020 minus.n19 minus.n5 28.4823
R2021 minus.n56 minus.n42 28.4823
R2022 minus.n63 minus.n62 28.4823
R2023 minus.n29 minus.n28 25.5611
R2024 minus.n15 minus.n14 25.5611
R2025 minus.n52 minus.n51 25.5611
R2026 minus.n66 minus.n65 25.5611
R2027 minus.n34 minus.n33 12.4157
R2028 minus.n8 minus.n7 12.4157
R2029 minus.n45 minus.n44 12.4157
R2030 minus.n71 minus.n70 12.4157
R2031 minus.n22 minus.n3 9.49444
R2032 minus.n21 minus.n20 9.49444
R2033 minus.n58 minus.n57 9.49444
R2034 minus.n59 minus.n40 9.49444
R2035 minus.n32 minus.n1 6.57323
R2036 minus.n13 minus.n12 6.57323
R2037 minus.n50 minus.n49 6.57323
R2038 minus.n69 minus.n38 6.57323
R2039 minus.n74 minus.n73 6.4702
R2040 minus.n36 minus.n0 0.189894
R2041 minus.n31 minus.n0 0.189894
R2042 minus.n31 minus.n30 0.189894
R2043 minus.n30 minus.n2 0.189894
R2044 minus.n24 minus.n2 0.189894
R2045 minus.n24 minus.n23 0.189894
R2046 minus.n23 minus.n4 0.189894
R2047 minus.n18 minus.n4 0.189894
R2048 minus.n18 minus.n17 0.189894
R2049 minus.n17 minus.n6 0.189894
R2050 minus.n11 minus.n6 0.189894
R2051 minus.n11 minus.n10 0.189894
R2052 minus.n48 minus.n47 0.189894
R2053 minus.n48 minus.n43 0.189894
R2054 minus.n54 minus.n43 0.189894
R2055 minus.n55 minus.n54 0.189894
R2056 minus.n55 minus.n41 0.189894
R2057 minus.n60 minus.n41 0.189894
R2058 minus.n61 minus.n60 0.189894
R2059 minus.n61 minus.n39 0.189894
R2060 minus.n67 minus.n39 0.189894
R2061 minus.n68 minus.n67 0.189894
R2062 minus.n68 minus.n37 0.189894
R2063 minus.n73 minus.n37 0.189894
R2064 minus minus.n74 0.188
R2065 drain_right.n7 drain_right.n5 59.2585
R2066 drain_right.n2 drain_right.n0 59.2585
R2067 drain_right.n13 drain_right.n11 59.2584
R2068 drain_right.n7 drain_right.n6 58.7154
R2069 drain_right.n9 drain_right.n8 58.7154
R2070 drain_right.n4 drain_right.n3 58.7154
R2071 drain_right.n2 drain_right.n1 58.7154
R2072 drain_right.n13 drain_right.n12 58.7154
R2073 drain_right.n15 drain_right.n14 58.7154
R2074 drain_right.n17 drain_right.n16 58.7154
R2075 drain_right.n19 drain_right.n18 58.7154
R2076 drain_right.n21 drain_right.n20 58.7154
R2077 drain_right drain_right.n10 41.8218
R2078 drain_right drain_right.n21 6.19632
R2079 drain_right.n5 drain_right.t10 0.7925
R2080 drain_right.n5 drain_right.t16 0.7925
R2081 drain_right.n6 drain_right.t6 0.7925
R2082 drain_right.n6 drain_right.t17 0.7925
R2083 drain_right.n8 drain_right.t13 0.7925
R2084 drain_right.n8 drain_right.t3 0.7925
R2085 drain_right.n3 drain_right.t12 0.7925
R2086 drain_right.n3 drain_right.t0 0.7925
R2087 drain_right.n1 drain_right.t19 0.7925
R2088 drain_right.n1 drain_right.t8 0.7925
R2089 drain_right.n0 drain_right.t18 0.7925
R2090 drain_right.n0 drain_right.t7 0.7925
R2091 drain_right.n11 drain_right.t2 0.7925
R2092 drain_right.n11 drain_right.t9 0.7925
R2093 drain_right.n12 drain_right.t11 0.7925
R2094 drain_right.n12 drain_right.t22 0.7925
R2095 drain_right.n14 drain_right.t23 0.7925
R2096 drain_right.n14 drain_right.t5 0.7925
R2097 drain_right.n16 drain_right.t1 0.7925
R2098 drain_right.n16 drain_right.t15 0.7925
R2099 drain_right.n18 drain_right.t14 0.7925
R2100 drain_right.n18 drain_right.t21 0.7925
R2101 drain_right.n20 drain_right.t20 0.7925
R2102 drain_right.n20 drain_right.t4 0.7925
R2103 drain_right.n9 drain_right.n7 0.543603
R2104 drain_right.n4 drain_right.n2 0.543603
R2105 drain_right.n21 drain_right.n19 0.543603
R2106 drain_right.n19 drain_right.n17 0.543603
R2107 drain_right.n17 drain_right.n15 0.543603
R2108 drain_right.n15 drain_right.n13 0.543603
R2109 drain_right.n10 drain_right.n9 0.216706
R2110 drain_right.n10 drain_right.n4 0.216706
C0 source drain_right 88.428795f
C1 drain_left drain_right 1.26597f
C2 drain_right plus 0.387992f
C3 drain_right minus 16.8494f
C4 source drain_left 88.4281f
C5 source plus 16.1485f
C6 drain_left plus 17.0816f
C7 source minus 16.134401f
C8 drain_left minus 0.172624f
C9 plus minus 8.50142f
C10 drain_right a_n2354_n5888# 10.063859f
C11 drain_left a_n2354_n5888# 10.41868f
C12 source a_n2354_n5888# 15.864443f
C13 minus a_n2354_n5888# 10.15463f
C14 plus a_n2354_n5888# 13.01519f
C15 drain_right.t18 a_n2354_n5888# 0.682201f
C16 drain_right.t7 a_n2354_n5888# 0.682201f
C17 drain_right.n0 a_n2354_n5888# 6.29113f
C18 drain_right.t19 a_n2354_n5888# 0.682201f
C19 drain_right.t8 a_n2354_n5888# 0.682201f
C20 drain_right.n1 a_n2354_n5888# 6.28722f
C21 drain_right.n2 a_n2354_n5888# 0.835508f
C22 drain_right.t12 a_n2354_n5888# 0.682201f
C23 drain_right.t0 a_n2354_n5888# 0.682201f
C24 drain_right.n3 a_n2354_n5888# 6.28722f
C25 drain_right.n4 a_n2354_n5888# 0.380084f
C26 drain_right.t10 a_n2354_n5888# 0.682201f
C27 drain_right.t16 a_n2354_n5888# 0.682201f
C28 drain_right.n5 a_n2354_n5888# 6.29113f
C29 drain_right.t6 a_n2354_n5888# 0.682201f
C30 drain_right.t17 a_n2354_n5888# 0.682201f
C31 drain_right.n6 a_n2354_n5888# 6.28722f
C32 drain_right.n7 a_n2354_n5888# 0.835508f
C33 drain_right.t13 a_n2354_n5888# 0.682201f
C34 drain_right.t3 a_n2354_n5888# 0.682201f
C35 drain_right.n8 a_n2354_n5888# 6.28722f
C36 drain_right.n9 a_n2354_n5888# 0.380084f
C37 drain_right.n10 a_n2354_n5888# 2.93314f
C38 drain_right.t2 a_n2354_n5888# 0.682201f
C39 drain_right.t9 a_n2354_n5888# 0.682201f
C40 drain_right.n11 a_n2354_n5888# 6.29111f
C41 drain_right.t11 a_n2354_n5888# 0.682201f
C42 drain_right.t22 a_n2354_n5888# 0.682201f
C43 drain_right.n12 a_n2354_n5888# 6.28722f
C44 drain_right.n13 a_n2354_n5888# 0.83552f
C45 drain_right.t23 a_n2354_n5888# 0.682201f
C46 drain_right.t5 a_n2354_n5888# 0.682201f
C47 drain_right.n14 a_n2354_n5888# 6.28722f
C48 drain_right.n15 a_n2354_n5888# 0.412753f
C49 drain_right.t1 a_n2354_n5888# 0.682201f
C50 drain_right.t15 a_n2354_n5888# 0.682201f
C51 drain_right.n16 a_n2354_n5888# 6.28722f
C52 drain_right.n17 a_n2354_n5888# 0.412753f
C53 drain_right.t14 a_n2354_n5888# 0.682201f
C54 drain_right.t21 a_n2354_n5888# 0.682201f
C55 drain_right.n18 a_n2354_n5888# 6.28722f
C56 drain_right.n19 a_n2354_n5888# 0.412753f
C57 drain_right.t20 a_n2354_n5888# 0.682201f
C58 drain_right.t4 a_n2354_n5888# 0.682201f
C59 drain_right.n20 a_n2354_n5888# 6.28722f
C60 drain_right.n21 a_n2354_n5888# 0.700182f
C61 minus.n0 a_n2354_n5888# 0.048622f
C62 minus.t3 a_n2354_n5888# 1.03153f
C63 minus.t19 a_n2354_n5888# 1.02606f
C64 minus.t9 a_n2354_n5888# 1.02606f
C65 minus.n1 a_n2354_n5888# 0.37336f
C66 minus.n2 a_n2354_n5888# 0.048622f
C67 minus.t2 a_n2354_n5888# 1.02606f
C68 minus.t22 a_n2354_n5888# 1.02606f
C69 minus.t8 a_n2354_n5888# 1.02606f
C70 minus.n3 a_n2354_n5888# 0.37336f
C71 minus.n4 a_n2354_n5888# 0.048622f
C72 minus.t0 a_n2354_n5888# 1.02606f
C73 minus.t18 a_n2354_n5888# 1.02606f
C74 minus.n5 a_n2354_n5888# 0.37336f
C75 minus.n6 a_n2354_n5888# 0.048622f
C76 minus.t12 a_n2354_n5888# 1.02606f
C77 minus.t1 a_n2354_n5888# 1.02606f
C78 minus.n7 a_n2354_n5888# 0.018678f
C79 minus.t21 a_n2354_n5888# 1.02606f
C80 minus.n8 a_n2354_n5888# 0.37336f
C81 minus.t14 a_n2354_n5888# 1.03153f
C82 minus.n9 a_n2354_n5888# 0.388427f
C83 minus.n10 a_n2354_n5888# 0.104075f
C84 minus.n11 a_n2354_n5888# 0.048622f
C85 minus.n12 a_n2354_n5888# 0.017479f
C86 minus.n13 a_n2354_n5888# 0.37336f
C87 minus.n14 a_n2354_n5888# 0.020027f
C88 minus.n15 a_n2354_n5888# 0.37336f
C89 minus.n16 a_n2354_n5888# 0.020027f
C90 minus.n17 a_n2354_n5888# 0.048622f
C91 minus.n18 a_n2354_n5888# 0.048622f
C92 minus.n19 a_n2354_n5888# 0.020027f
C93 minus.n20 a_n2354_n5888# 0.37336f
C94 minus.n21 a_n2354_n5888# 0.018078f
C95 minus.n22 a_n2354_n5888# 0.018078f
C96 minus.n23 a_n2354_n5888# 0.048622f
C97 minus.n24 a_n2354_n5888# 0.048622f
C98 minus.n25 a_n2354_n5888# 0.020027f
C99 minus.n26 a_n2354_n5888# 0.37336f
C100 minus.n27 a_n2354_n5888# 0.020027f
C101 minus.n28 a_n2354_n5888# 0.37336f
C102 minus.n29 a_n2354_n5888# 0.020027f
C103 minus.n30 a_n2354_n5888# 0.048622f
C104 minus.n31 a_n2354_n5888# 0.048622f
C105 minus.n32 a_n2354_n5888# 0.017479f
C106 minus.n33 a_n2354_n5888# 0.018678f
C107 minus.n34 a_n2354_n5888# 0.37336f
C108 minus.n35 a_n2354_n5888# 0.388362f
C109 minus.n36 a_n2354_n5888# 2.59722f
C110 minus.n37 a_n2354_n5888# 0.048622f
C111 minus.t13 a_n2354_n5888# 1.02606f
C112 minus.t6 a_n2354_n5888# 1.02606f
C113 minus.n38 a_n2354_n5888# 0.37336f
C114 minus.n39 a_n2354_n5888# 0.048622f
C115 minus.t17 a_n2354_n5888# 1.02606f
C116 minus.t20 a_n2354_n5888# 1.02606f
C117 minus.t10 a_n2354_n5888# 1.02606f
C118 minus.n40 a_n2354_n5888# 0.37336f
C119 minus.n41 a_n2354_n5888# 0.048622f
C120 minus.t23 a_n2354_n5888# 1.02606f
C121 minus.t11 a_n2354_n5888# 1.02606f
C122 minus.n42 a_n2354_n5888# 0.37336f
C123 minus.n43 a_n2354_n5888# 0.048622f
C124 minus.t15 a_n2354_n5888# 1.02606f
C125 minus.t4 a_n2354_n5888# 1.02606f
C126 minus.n44 a_n2354_n5888# 0.018678f
C127 minus.t5 a_n2354_n5888# 1.03153f
C128 minus.t16 a_n2354_n5888# 1.02606f
C129 minus.n45 a_n2354_n5888# 0.37336f
C130 minus.n46 a_n2354_n5888# 0.388427f
C131 minus.n47 a_n2354_n5888# 0.104075f
C132 minus.n48 a_n2354_n5888# 0.048622f
C133 minus.n49 a_n2354_n5888# 0.017479f
C134 minus.n50 a_n2354_n5888# 0.37336f
C135 minus.n51 a_n2354_n5888# 0.020027f
C136 minus.n52 a_n2354_n5888# 0.37336f
C137 minus.n53 a_n2354_n5888# 0.020027f
C138 minus.n54 a_n2354_n5888# 0.048622f
C139 minus.n55 a_n2354_n5888# 0.048622f
C140 minus.n56 a_n2354_n5888# 0.020027f
C141 minus.n57 a_n2354_n5888# 0.37336f
C142 minus.n58 a_n2354_n5888# 0.018078f
C143 minus.n59 a_n2354_n5888# 0.018078f
C144 minus.n60 a_n2354_n5888# 0.048622f
C145 minus.n61 a_n2354_n5888# 0.048622f
C146 minus.n62 a_n2354_n5888# 0.020027f
C147 minus.n63 a_n2354_n5888# 0.37336f
C148 minus.n64 a_n2354_n5888# 0.020027f
C149 minus.n65 a_n2354_n5888# 0.37336f
C150 minus.n66 a_n2354_n5888# 0.020027f
C151 minus.n67 a_n2354_n5888# 0.048622f
C152 minus.n68 a_n2354_n5888# 0.048622f
C153 minus.n69 a_n2354_n5888# 0.017479f
C154 minus.n70 a_n2354_n5888# 0.018678f
C155 minus.n71 a_n2354_n5888# 0.37336f
C156 minus.t7 a_n2354_n5888# 1.03153f
C157 minus.n72 a_n2354_n5888# 0.388362f
C158 minus.n73 a_n2354_n5888# 0.314462f
C159 minus.n74 a_n2354_n5888# 3.05319f
C160 source.n0 a_n2354_n5888# 0.041229f
C161 source.n1 a_n2354_n5888# 0.029906f
C162 source.n2 a_n2354_n5888# 0.01607f
C163 source.n3 a_n2354_n5888# 0.037984f
C164 source.n4 a_n2354_n5888# 0.017016f
C165 source.n5 a_n2354_n5888# 0.029906f
C166 source.n6 a_n2354_n5888# 0.01607f
C167 source.n7 a_n2354_n5888# 0.037984f
C168 source.n8 a_n2354_n5888# 0.017016f
C169 source.n9 a_n2354_n5888# 0.029906f
C170 source.n10 a_n2354_n5888# 0.01607f
C171 source.n11 a_n2354_n5888# 0.037984f
C172 source.n12 a_n2354_n5888# 0.017016f
C173 source.n13 a_n2354_n5888# 0.029906f
C174 source.n14 a_n2354_n5888# 0.01607f
C175 source.n15 a_n2354_n5888# 0.037984f
C176 source.n16 a_n2354_n5888# 0.037984f
C177 source.n17 a_n2354_n5888# 0.017016f
C178 source.n18 a_n2354_n5888# 0.029906f
C179 source.n19 a_n2354_n5888# 0.01607f
C180 source.n20 a_n2354_n5888# 0.037984f
C181 source.n21 a_n2354_n5888# 0.017016f
C182 source.n22 a_n2354_n5888# 0.029906f
C183 source.n23 a_n2354_n5888# 0.01607f
C184 source.n24 a_n2354_n5888# 0.037984f
C185 source.n25 a_n2354_n5888# 0.017016f
C186 source.n26 a_n2354_n5888# 0.029906f
C187 source.n27 a_n2354_n5888# 0.01607f
C188 source.n28 a_n2354_n5888# 0.037984f
C189 source.n29 a_n2354_n5888# 0.017016f
C190 source.n30 a_n2354_n5888# 0.029906f
C191 source.n31 a_n2354_n5888# 0.01607f
C192 source.n32 a_n2354_n5888# 0.037984f
C193 source.n33 a_n2354_n5888# 0.017016f
C194 source.n34 a_n2354_n5888# 0.029906f
C195 source.n35 a_n2354_n5888# 0.016543f
C196 source.n36 a_n2354_n5888# 0.037984f
C197 source.n37 a_n2354_n5888# 0.01607f
C198 source.n38 a_n2354_n5888# 0.017016f
C199 source.n39 a_n2354_n5888# 0.029906f
C200 source.n40 a_n2354_n5888# 0.01607f
C201 source.n41 a_n2354_n5888# 0.037984f
C202 source.n42 a_n2354_n5888# 0.017016f
C203 source.n43 a_n2354_n5888# 0.029906f
C204 source.n44 a_n2354_n5888# 0.01607f
C205 source.n45 a_n2354_n5888# 0.028488f
C206 source.n46 a_n2354_n5888# 0.026852f
C207 source.t42 a_n2354_n5888# 0.066247f
C208 source.n47 a_n2354_n5888# 0.364881f
C209 source.n48 a_n2354_n5888# 3.23796f
C210 source.n49 a_n2354_n5888# 0.01607f
C211 source.n50 a_n2354_n5888# 0.017016f
C212 source.n51 a_n2354_n5888# 0.037984f
C213 source.n52 a_n2354_n5888# 0.037984f
C214 source.n53 a_n2354_n5888# 0.017016f
C215 source.n54 a_n2354_n5888# 0.01607f
C216 source.n55 a_n2354_n5888# 0.029906f
C217 source.n56 a_n2354_n5888# 0.029906f
C218 source.n57 a_n2354_n5888# 0.01607f
C219 source.n58 a_n2354_n5888# 0.017016f
C220 source.n59 a_n2354_n5888# 0.037984f
C221 source.n60 a_n2354_n5888# 0.037984f
C222 source.n61 a_n2354_n5888# 0.017016f
C223 source.n62 a_n2354_n5888# 0.01607f
C224 source.n63 a_n2354_n5888# 0.029906f
C225 source.n64 a_n2354_n5888# 0.029906f
C226 source.n65 a_n2354_n5888# 0.01607f
C227 source.n66 a_n2354_n5888# 0.017016f
C228 source.n67 a_n2354_n5888# 0.037984f
C229 source.n68 a_n2354_n5888# 0.037984f
C230 source.n69 a_n2354_n5888# 0.037984f
C231 source.n70 a_n2354_n5888# 0.016543f
C232 source.n71 a_n2354_n5888# 0.01607f
C233 source.n72 a_n2354_n5888# 0.029906f
C234 source.n73 a_n2354_n5888# 0.029906f
C235 source.n74 a_n2354_n5888# 0.01607f
C236 source.n75 a_n2354_n5888# 0.017016f
C237 source.n76 a_n2354_n5888# 0.037984f
C238 source.n77 a_n2354_n5888# 0.037984f
C239 source.n78 a_n2354_n5888# 0.017016f
C240 source.n79 a_n2354_n5888# 0.01607f
C241 source.n80 a_n2354_n5888# 0.029906f
C242 source.n81 a_n2354_n5888# 0.029906f
C243 source.n82 a_n2354_n5888# 0.01607f
C244 source.n83 a_n2354_n5888# 0.017016f
C245 source.n84 a_n2354_n5888# 0.037984f
C246 source.n85 a_n2354_n5888# 0.037984f
C247 source.n86 a_n2354_n5888# 0.017016f
C248 source.n87 a_n2354_n5888# 0.01607f
C249 source.n88 a_n2354_n5888# 0.029906f
C250 source.n89 a_n2354_n5888# 0.029906f
C251 source.n90 a_n2354_n5888# 0.01607f
C252 source.n91 a_n2354_n5888# 0.017016f
C253 source.n92 a_n2354_n5888# 0.037984f
C254 source.n93 a_n2354_n5888# 0.037984f
C255 source.n94 a_n2354_n5888# 0.017016f
C256 source.n95 a_n2354_n5888# 0.01607f
C257 source.n96 a_n2354_n5888# 0.029906f
C258 source.n97 a_n2354_n5888# 0.029906f
C259 source.n98 a_n2354_n5888# 0.01607f
C260 source.n99 a_n2354_n5888# 0.017016f
C261 source.n100 a_n2354_n5888# 0.037984f
C262 source.n101 a_n2354_n5888# 0.037984f
C263 source.n102 a_n2354_n5888# 0.017016f
C264 source.n103 a_n2354_n5888# 0.01607f
C265 source.n104 a_n2354_n5888# 0.029906f
C266 source.n105 a_n2354_n5888# 0.029906f
C267 source.n106 a_n2354_n5888# 0.01607f
C268 source.n107 a_n2354_n5888# 0.017016f
C269 source.n108 a_n2354_n5888# 0.037984f
C270 source.n109 a_n2354_n5888# 0.037984f
C271 source.n110 a_n2354_n5888# 0.017016f
C272 source.n111 a_n2354_n5888# 0.01607f
C273 source.n112 a_n2354_n5888# 0.029906f
C274 source.n113 a_n2354_n5888# 0.029906f
C275 source.n114 a_n2354_n5888# 0.01607f
C276 source.n115 a_n2354_n5888# 0.016543f
C277 source.n116 a_n2354_n5888# 0.016543f
C278 source.n117 a_n2354_n5888# 0.037984f
C279 source.n118 a_n2354_n5888# 0.037984f
C280 source.n119 a_n2354_n5888# 0.017016f
C281 source.n120 a_n2354_n5888# 0.01607f
C282 source.n121 a_n2354_n5888# 0.029906f
C283 source.n122 a_n2354_n5888# 0.029906f
C284 source.n123 a_n2354_n5888# 0.01607f
C285 source.n124 a_n2354_n5888# 0.017016f
C286 source.n125 a_n2354_n5888# 0.037984f
C287 source.n126 a_n2354_n5888# 0.037984f
C288 source.n127 a_n2354_n5888# 0.017016f
C289 source.n128 a_n2354_n5888# 0.01607f
C290 source.n129 a_n2354_n5888# 0.029906f
C291 source.n130 a_n2354_n5888# 0.029906f
C292 source.n131 a_n2354_n5888# 0.01607f
C293 source.n132 a_n2354_n5888# 0.017016f
C294 source.n133 a_n2354_n5888# 0.037984f
C295 source.n134 a_n2354_n5888# 0.080802f
C296 source.n135 a_n2354_n5888# 0.017016f
C297 source.n136 a_n2354_n5888# 0.01607f
C298 source.n137 a_n2354_n5888# 0.065858f
C299 source.n138 a_n2354_n5888# 0.044963f
C300 source.n139 a_n2354_n5888# 2.35039f
C301 source.t30 a_n2354_n5888# 0.59082f
C302 source.t47 a_n2354_n5888# 0.59082f
C303 source.n140 a_n2354_n5888# 5.347f
C304 source.n141 a_n2354_n5888# 0.414858f
C305 source.t46 a_n2354_n5888# 0.59082f
C306 source.t37 a_n2354_n5888# 0.59082f
C307 source.n142 a_n2354_n5888# 5.347f
C308 source.n143 a_n2354_n5888# 0.414858f
C309 source.t34 a_n2354_n5888# 0.59082f
C310 source.t27 a_n2354_n5888# 0.59082f
C311 source.n144 a_n2354_n5888# 5.347f
C312 source.n145 a_n2354_n5888# 0.414858f
C313 source.t26 a_n2354_n5888# 0.59082f
C314 source.t39 a_n2354_n5888# 0.59082f
C315 source.n146 a_n2354_n5888# 5.347f
C316 source.n147 a_n2354_n5888# 0.414858f
C317 source.t38 a_n2354_n5888# 0.59082f
C318 source.t32 a_n2354_n5888# 0.59082f
C319 source.n148 a_n2354_n5888# 5.347f
C320 source.n149 a_n2354_n5888# 0.414858f
C321 source.n150 a_n2354_n5888# 0.041229f
C322 source.n151 a_n2354_n5888# 0.029906f
C323 source.n152 a_n2354_n5888# 0.01607f
C324 source.n153 a_n2354_n5888# 0.037984f
C325 source.n154 a_n2354_n5888# 0.017016f
C326 source.n155 a_n2354_n5888# 0.029906f
C327 source.n156 a_n2354_n5888# 0.01607f
C328 source.n157 a_n2354_n5888# 0.037984f
C329 source.n158 a_n2354_n5888# 0.017016f
C330 source.n159 a_n2354_n5888# 0.029906f
C331 source.n160 a_n2354_n5888# 0.01607f
C332 source.n161 a_n2354_n5888# 0.037984f
C333 source.n162 a_n2354_n5888# 0.017016f
C334 source.n163 a_n2354_n5888# 0.029906f
C335 source.n164 a_n2354_n5888# 0.01607f
C336 source.n165 a_n2354_n5888# 0.037984f
C337 source.n166 a_n2354_n5888# 0.037984f
C338 source.n167 a_n2354_n5888# 0.017016f
C339 source.n168 a_n2354_n5888# 0.029906f
C340 source.n169 a_n2354_n5888# 0.01607f
C341 source.n170 a_n2354_n5888# 0.037984f
C342 source.n171 a_n2354_n5888# 0.017016f
C343 source.n172 a_n2354_n5888# 0.029906f
C344 source.n173 a_n2354_n5888# 0.01607f
C345 source.n174 a_n2354_n5888# 0.037984f
C346 source.n175 a_n2354_n5888# 0.017016f
C347 source.n176 a_n2354_n5888# 0.029906f
C348 source.n177 a_n2354_n5888# 0.01607f
C349 source.n178 a_n2354_n5888# 0.037984f
C350 source.n179 a_n2354_n5888# 0.017016f
C351 source.n180 a_n2354_n5888# 0.029906f
C352 source.n181 a_n2354_n5888# 0.01607f
C353 source.n182 a_n2354_n5888# 0.037984f
C354 source.n183 a_n2354_n5888# 0.017016f
C355 source.n184 a_n2354_n5888# 0.029906f
C356 source.n185 a_n2354_n5888# 0.016543f
C357 source.n186 a_n2354_n5888# 0.037984f
C358 source.n187 a_n2354_n5888# 0.01607f
C359 source.n188 a_n2354_n5888# 0.017016f
C360 source.n189 a_n2354_n5888# 0.029906f
C361 source.n190 a_n2354_n5888# 0.01607f
C362 source.n191 a_n2354_n5888# 0.037984f
C363 source.n192 a_n2354_n5888# 0.017016f
C364 source.n193 a_n2354_n5888# 0.029906f
C365 source.n194 a_n2354_n5888# 0.01607f
C366 source.n195 a_n2354_n5888# 0.028488f
C367 source.n196 a_n2354_n5888# 0.026852f
C368 source.t45 a_n2354_n5888# 0.066247f
C369 source.n197 a_n2354_n5888# 0.364881f
C370 source.n198 a_n2354_n5888# 3.23796f
C371 source.n199 a_n2354_n5888# 0.01607f
C372 source.n200 a_n2354_n5888# 0.017016f
C373 source.n201 a_n2354_n5888# 0.037984f
C374 source.n202 a_n2354_n5888# 0.037984f
C375 source.n203 a_n2354_n5888# 0.017016f
C376 source.n204 a_n2354_n5888# 0.01607f
C377 source.n205 a_n2354_n5888# 0.029906f
C378 source.n206 a_n2354_n5888# 0.029906f
C379 source.n207 a_n2354_n5888# 0.01607f
C380 source.n208 a_n2354_n5888# 0.017016f
C381 source.n209 a_n2354_n5888# 0.037984f
C382 source.n210 a_n2354_n5888# 0.037984f
C383 source.n211 a_n2354_n5888# 0.017016f
C384 source.n212 a_n2354_n5888# 0.01607f
C385 source.n213 a_n2354_n5888# 0.029906f
C386 source.n214 a_n2354_n5888# 0.029906f
C387 source.n215 a_n2354_n5888# 0.01607f
C388 source.n216 a_n2354_n5888# 0.017016f
C389 source.n217 a_n2354_n5888# 0.037984f
C390 source.n218 a_n2354_n5888# 0.037984f
C391 source.n219 a_n2354_n5888# 0.037984f
C392 source.n220 a_n2354_n5888# 0.016543f
C393 source.n221 a_n2354_n5888# 0.01607f
C394 source.n222 a_n2354_n5888# 0.029906f
C395 source.n223 a_n2354_n5888# 0.029906f
C396 source.n224 a_n2354_n5888# 0.01607f
C397 source.n225 a_n2354_n5888# 0.017016f
C398 source.n226 a_n2354_n5888# 0.037984f
C399 source.n227 a_n2354_n5888# 0.037984f
C400 source.n228 a_n2354_n5888# 0.017016f
C401 source.n229 a_n2354_n5888# 0.01607f
C402 source.n230 a_n2354_n5888# 0.029906f
C403 source.n231 a_n2354_n5888# 0.029906f
C404 source.n232 a_n2354_n5888# 0.01607f
C405 source.n233 a_n2354_n5888# 0.017016f
C406 source.n234 a_n2354_n5888# 0.037984f
C407 source.n235 a_n2354_n5888# 0.037984f
C408 source.n236 a_n2354_n5888# 0.017016f
C409 source.n237 a_n2354_n5888# 0.01607f
C410 source.n238 a_n2354_n5888# 0.029906f
C411 source.n239 a_n2354_n5888# 0.029906f
C412 source.n240 a_n2354_n5888# 0.01607f
C413 source.n241 a_n2354_n5888# 0.017016f
C414 source.n242 a_n2354_n5888# 0.037984f
C415 source.n243 a_n2354_n5888# 0.037984f
C416 source.n244 a_n2354_n5888# 0.017016f
C417 source.n245 a_n2354_n5888# 0.01607f
C418 source.n246 a_n2354_n5888# 0.029906f
C419 source.n247 a_n2354_n5888# 0.029906f
C420 source.n248 a_n2354_n5888# 0.01607f
C421 source.n249 a_n2354_n5888# 0.017016f
C422 source.n250 a_n2354_n5888# 0.037984f
C423 source.n251 a_n2354_n5888# 0.037984f
C424 source.n252 a_n2354_n5888# 0.017016f
C425 source.n253 a_n2354_n5888# 0.01607f
C426 source.n254 a_n2354_n5888# 0.029906f
C427 source.n255 a_n2354_n5888# 0.029906f
C428 source.n256 a_n2354_n5888# 0.01607f
C429 source.n257 a_n2354_n5888# 0.017016f
C430 source.n258 a_n2354_n5888# 0.037984f
C431 source.n259 a_n2354_n5888# 0.037984f
C432 source.n260 a_n2354_n5888# 0.017016f
C433 source.n261 a_n2354_n5888# 0.01607f
C434 source.n262 a_n2354_n5888# 0.029906f
C435 source.n263 a_n2354_n5888# 0.029906f
C436 source.n264 a_n2354_n5888# 0.01607f
C437 source.n265 a_n2354_n5888# 0.016543f
C438 source.n266 a_n2354_n5888# 0.016543f
C439 source.n267 a_n2354_n5888# 0.037984f
C440 source.n268 a_n2354_n5888# 0.037984f
C441 source.n269 a_n2354_n5888# 0.017016f
C442 source.n270 a_n2354_n5888# 0.01607f
C443 source.n271 a_n2354_n5888# 0.029906f
C444 source.n272 a_n2354_n5888# 0.029906f
C445 source.n273 a_n2354_n5888# 0.01607f
C446 source.n274 a_n2354_n5888# 0.017016f
C447 source.n275 a_n2354_n5888# 0.037984f
C448 source.n276 a_n2354_n5888# 0.037984f
C449 source.n277 a_n2354_n5888# 0.017016f
C450 source.n278 a_n2354_n5888# 0.01607f
C451 source.n279 a_n2354_n5888# 0.029906f
C452 source.n280 a_n2354_n5888# 0.029906f
C453 source.n281 a_n2354_n5888# 0.01607f
C454 source.n282 a_n2354_n5888# 0.017016f
C455 source.n283 a_n2354_n5888# 0.037984f
C456 source.n284 a_n2354_n5888# 0.080802f
C457 source.n285 a_n2354_n5888# 0.017016f
C458 source.n286 a_n2354_n5888# 0.01607f
C459 source.n287 a_n2354_n5888# 0.065858f
C460 source.n288 a_n2354_n5888# 0.044963f
C461 source.n289 a_n2354_n5888# 0.12131f
C462 source.n290 a_n2354_n5888# 0.041229f
C463 source.n291 a_n2354_n5888# 0.029906f
C464 source.n292 a_n2354_n5888# 0.01607f
C465 source.n293 a_n2354_n5888# 0.037984f
C466 source.n294 a_n2354_n5888# 0.017016f
C467 source.n295 a_n2354_n5888# 0.029906f
C468 source.n296 a_n2354_n5888# 0.01607f
C469 source.n297 a_n2354_n5888# 0.037984f
C470 source.n298 a_n2354_n5888# 0.017016f
C471 source.n299 a_n2354_n5888# 0.029906f
C472 source.n300 a_n2354_n5888# 0.01607f
C473 source.n301 a_n2354_n5888# 0.037984f
C474 source.n302 a_n2354_n5888# 0.017016f
C475 source.n303 a_n2354_n5888# 0.029906f
C476 source.n304 a_n2354_n5888# 0.01607f
C477 source.n305 a_n2354_n5888# 0.037984f
C478 source.n306 a_n2354_n5888# 0.037984f
C479 source.n307 a_n2354_n5888# 0.017016f
C480 source.n308 a_n2354_n5888# 0.029906f
C481 source.n309 a_n2354_n5888# 0.01607f
C482 source.n310 a_n2354_n5888# 0.037984f
C483 source.n311 a_n2354_n5888# 0.017016f
C484 source.n312 a_n2354_n5888# 0.029906f
C485 source.n313 a_n2354_n5888# 0.01607f
C486 source.n314 a_n2354_n5888# 0.037984f
C487 source.n315 a_n2354_n5888# 0.017016f
C488 source.n316 a_n2354_n5888# 0.029906f
C489 source.n317 a_n2354_n5888# 0.01607f
C490 source.n318 a_n2354_n5888# 0.037984f
C491 source.n319 a_n2354_n5888# 0.017016f
C492 source.n320 a_n2354_n5888# 0.029906f
C493 source.n321 a_n2354_n5888# 0.01607f
C494 source.n322 a_n2354_n5888# 0.037984f
C495 source.n323 a_n2354_n5888# 0.017016f
C496 source.n324 a_n2354_n5888# 0.029906f
C497 source.n325 a_n2354_n5888# 0.016543f
C498 source.n326 a_n2354_n5888# 0.037984f
C499 source.n327 a_n2354_n5888# 0.01607f
C500 source.n328 a_n2354_n5888# 0.017016f
C501 source.n329 a_n2354_n5888# 0.029906f
C502 source.n330 a_n2354_n5888# 0.01607f
C503 source.n331 a_n2354_n5888# 0.037984f
C504 source.n332 a_n2354_n5888# 0.017016f
C505 source.n333 a_n2354_n5888# 0.029906f
C506 source.n334 a_n2354_n5888# 0.01607f
C507 source.n335 a_n2354_n5888# 0.028488f
C508 source.n336 a_n2354_n5888# 0.026852f
C509 source.t2 a_n2354_n5888# 0.066247f
C510 source.n337 a_n2354_n5888# 0.364881f
C511 source.n338 a_n2354_n5888# 3.23796f
C512 source.n339 a_n2354_n5888# 0.01607f
C513 source.n340 a_n2354_n5888# 0.017016f
C514 source.n341 a_n2354_n5888# 0.037984f
C515 source.n342 a_n2354_n5888# 0.037984f
C516 source.n343 a_n2354_n5888# 0.017016f
C517 source.n344 a_n2354_n5888# 0.01607f
C518 source.n345 a_n2354_n5888# 0.029906f
C519 source.n346 a_n2354_n5888# 0.029906f
C520 source.n347 a_n2354_n5888# 0.01607f
C521 source.n348 a_n2354_n5888# 0.017016f
C522 source.n349 a_n2354_n5888# 0.037984f
C523 source.n350 a_n2354_n5888# 0.037984f
C524 source.n351 a_n2354_n5888# 0.017016f
C525 source.n352 a_n2354_n5888# 0.01607f
C526 source.n353 a_n2354_n5888# 0.029906f
C527 source.n354 a_n2354_n5888# 0.029906f
C528 source.n355 a_n2354_n5888# 0.01607f
C529 source.n356 a_n2354_n5888# 0.017016f
C530 source.n357 a_n2354_n5888# 0.037984f
C531 source.n358 a_n2354_n5888# 0.037984f
C532 source.n359 a_n2354_n5888# 0.037984f
C533 source.n360 a_n2354_n5888# 0.016543f
C534 source.n361 a_n2354_n5888# 0.01607f
C535 source.n362 a_n2354_n5888# 0.029906f
C536 source.n363 a_n2354_n5888# 0.029906f
C537 source.n364 a_n2354_n5888# 0.01607f
C538 source.n365 a_n2354_n5888# 0.017016f
C539 source.n366 a_n2354_n5888# 0.037984f
C540 source.n367 a_n2354_n5888# 0.037984f
C541 source.n368 a_n2354_n5888# 0.017016f
C542 source.n369 a_n2354_n5888# 0.01607f
C543 source.n370 a_n2354_n5888# 0.029906f
C544 source.n371 a_n2354_n5888# 0.029906f
C545 source.n372 a_n2354_n5888# 0.01607f
C546 source.n373 a_n2354_n5888# 0.017016f
C547 source.n374 a_n2354_n5888# 0.037984f
C548 source.n375 a_n2354_n5888# 0.037984f
C549 source.n376 a_n2354_n5888# 0.017016f
C550 source.n377 a_n2354_n5888# 0.01607f
C551 source.n378 a_n2354_n5888# 0.029906f
C552 source.n379 a_n2354_n5888# 0.029906f
C553 source.n380 a_n2354_n5888# 0.01607f
C554 source.n381 a_n2354_n5888# 0.017016f
C555 source.n382 a_n2354_n5888# 0.037984f
C556 source.n383 a_n2354_n5888# 0.037984f
C557 source.n384 a_n2354_n5888# 0.017016f
C558 source.n385 a_n2354_n5888# 0.01607f
C559 source.n386 a_n2354_n5888# 0.029906f
C560 source.n387 a_n2354_n5888# 0.029906f
C561 source.n388 a_n2354_n5888# 0.01607f
C562 source.n389 a_n2354_n5888# 0.017016f
C563 source.n390 a_n2354_n5888# 0.037984f
C564 source.n391 a_n2354_n5888# 0.037984f
C565 source.n392 a_n2354_n5888# 0.017016f
C566 source.n393 a_n2354_n5888# 0.01607f
C567 source.n394 a_n2354_n5888# 0.029906f
C568 source.n395 a_n2354_n5888# 0.029906f
C569 source.n396 a_n2354_n5888# 0.01607f
C570 source.n397 a_n2354_n5888# 0.017016f
C571 source.n398 a_n2354_n5888# 0.037984f
C572 source.n399 a_n2354_n5888# 0.037984f
C573 source.n400 a_n2354_n5888# 0.017016f
C574 source.n401 a_n2354_n5888# 0.01607f
C575 source.n402 a_n2354_n5888# 0.029906f
C576 source.n403 a_n2354_n5888# 0.029906f
C577 source.n404 a_n2354_n5888# 0.01607f
C578 source.n405 a_n2354_n5888# 0.016543f
C579 source.n406 a_n2354_n5888# 0.016543f
C580 source.n407 a_n2354_n5888# 0.037984f
C581 source.n408 a_n2354_n5888# 0.037984f
C582 source.n409 a_n2354_n5888# 0.017016f
C583 source.n410 a_n2354_n5888# 0.01607f
C584 source.n411 a_n2354_n5888# 0.029906f
C585 source.n412 a_n2354_n5888# 0.029906f
C586 source.n413 a_n2354_n5888# 0.01607f
C587 source.n414 a_n2354_n5888# 0.017016f
C588 source.n415 a_n2354_n5888# 0.037984f
C589 source.n416 a_n2354_n5888# 0.037984f
C590 source.n417 a_n2354_n5888# 0.017016f
C591 source.n418 a_n2354_n5888# 0.01607f
C592 source.n419 a_n2354_n5888# 0.029906f
C593 source.n420 a_n2354_n5888# 0.029906f
C594 source.n421 a_n2354_n5888# 0.01607f
C595 source.n422 a_n2354_n5888# 0.017016f
C596 source.n423 a_n2354_n5888# 0.037984f
C597 source.n424 a_n2354_n5888# 0.080802f
C598 source.n425 a_n2354_n5888# 0.017016f
C599 source.n426 a_n2354_n5888# 0.01607f
C600 source.n427 a_n2354_n5888# 0.065858f
C601 source.n428 a_n2354_n5888# 0.044963f
C602 source.n429 a_n2354_n5888# 0.12131f
C603 source.t0 a_n2354_n5888# 0.59082f
C604 source.t17 a_n2354_n5888# 0.59082f
C605 source.n430 a_n2354_n5888# 5.347f
C606 source.n431 a_n2354_n5888# 0.414858f
C607 source.t1 a_n2354_n5888# 0.59082f
C608 source.t16 a_n2354_n5888# 0.59082f
C609 source.n432 a_n2354_n5888# 5.347f
C610 source.n433 a_n2354_n5888# 0.414858f
C611 source.t13 a_n2354_n5888# 0.59082f
C612 source.t6 a_n2354_n5888# 0.59082f
C613 source.n434 a_n2354_n5888# 5.347f
C614 source.n435 a_n2354_n5888# 0.414858f
C615 source.t20 a_n2354_n5888# 0.59082f
C616 source.t22 a_n2354_n5888# 0.59082f
C617 source.n436 a_n2354_n5888# 5.347f
C618 source.n437 a_n2354_n5888# 0.414858f
C619 source.t5 a_n2354_n5888# 0.59082f
C620 source.t15 a_n2354_n5888# 0.59082f
C621 source.n438 a_n2354_n5888# 5.347f
C622 source.n439 a_n2354_n5888# 0.414858f
C623 source.n440 a_n2354_n5888# 0.041229f
C624 source.n441 a_n2354_n5888# 0.029906f
C625 source.n442 a_n2354_n5888# 0.01607f
C626 source.n443 a_n2354_n5888# 0.037984f
C627 source.n444 a_n2354_n5888# 0.017016f
C628 source.n445 a_n2354_n5888# 0.029906f
C629 source.n446 a_n2354_n5888# 0.01607f
C630 source.n447 a_n2354_n5888# 0.037984f
C631 source.n448 a_n2354_n5888# 0.017016f
C632 source.n449 a_n2354_n5888# 0.029906f
C633 source.n450 a_n2354_n5888# 0.01607f
C634 source.n451 a_n2354_n5888# 0.037984f
C635 source.n452 a_n2354_n5888# 0.017016f
C636 source.n453 a_n2354_n5888# 0.029906f
C637 source.n454 a_n2354_n5888# 0.01607f
C638 source.n455 a_n2354_n5888# 0.037984f
C639 source.n456 a_n2354_n5888# 0.037984f
C640 source.n457 a_n2354_n5888# 0.017016f
C641 source.n458 a_n2354_n5888# 0.029906f
C642 source.n459 a_n2354_n5888# 0.01607f
C643 source.n460 a_n2354_n5888# 0.037984f
C644 source.n461 a_n2354_n5888# 0.017016f
C645 source.n462 a_n2354_n5888# 0.029906f
C646 source.n463 a_n2354_n5888# 0.01607f
C647 source.n464 a_n2354_n5888# 0.037984f
C648 source.n465 a_n2354_n5888# 0.017016f
C649 source.n466 a_n2354_n5888# 0.029906f
C650 source.n467 a_n2354_n5888# 0.01607f
C651 source.n468 a_n2354_n5888# 0.037984f
C652 source.n469 a_n2354_n5888# 0.017016f
C653 source.n470 a_n2354_n5888# 0.029906f
C654 source.n471 a_n2354_n5888# 0.01607f
C655 source.n472 a_n2354_n5888# 0.037984f
C656 source.n473 a_n2354_n5888# 0.017016f
C657 source.n474 a_n2354_n5888# 0.029906f
C658 source.n475 a_n2354_n5888# 0.016543f
C659 source.n476 a_n2354_n5888# 0.037984f
C660 source.n477 a_n2354_n5888# 0.01607f
C661 source.n478 a_n2354_n5888# 0.017016f
C662 source.n479 a_n2354_n5888# 0.029906f
C663 source.n480 a_n2354_n5888# 0.01607f
C664 source.n481 a_n2354_n5888# 0.037984f
C665 source.n482 a_n2354_n5888# 0.017016f
C666 source.n483 a_n2354_n5888# 0.029906f
C667 source.n484 a_n2354_n5888# 0.01607f
C668 source.n485 a_n2354_n5888# 0.028488f
C669 source.n486 a_n2354_n5888# 0.026852f
C670 source.t10 a_n2354_n5888# 0.066247f
C671 source.n487 a_n2354_n5888# 0.364881f
C672 source.n488 a_n2354_n5888# 3.23796f
C673 source.n489 a_n2354_n5888# 0.01607f
C674 source.n490 a_n2354_n5888# 0.017016f
C675 source.n491 a_n2354_n5888# 0.037984f
C676 source.n492 a_n2354_n5888# 0.037984f
C677 source.n493 a_n2354_n5888# 0.017016f
C678 source.n494 a_n2354_n5888# 0.01607f
C679 source.n495 a_n2354_n5888# 0.029906f
C680 source.n496 a_n2354_n5888# 0.029906f
C681 source.n497 a_n2354_n5888# 0.01607f
C682 source.n498 a_n2354_n5888# 0.017016f
C683 source.n499 a_n2354_n5888# 0.037984f
C684 source.n500 a_n2354_n5888# 0.037984f
C685 source.n501 a_n2354_n5888# 0.017016f
C686 source.n502 a_n2354_n5888# 0.01607f
C687 source.n503 a_n2354_n5888# 0.029906f
C688 source.n504 a_n2354_n5888# 0.029906f
C689 source.n505 a_n2354_n5888# 0.01607f
C690 source.n506 a_n2354_n5888# 0.017016f
C691 source.n507 a_n2354_n5888# 0.037984f
C692 source.n508 a_n2354_n5888# 0.037984f
C693 source.n509 a_n2354_n5888# 0.037984f
C694 source.n510 a_n2354_n5888# 0.016543f
C695 source.n511 a_n2354_n5888# 0.01607f
C696 source.n512 a_n2354_n5888# 0.029906f
C697 source.n513 a_n2354_n5888# 0.029906f
C698 source.n514 a_n2354_n5888# 0.01607f
C699 source.n515 a_n2354_n5888# 0.017016f
C700 source.n516 a_n2354_n5888# 0.037984f
C701 source.n517 a_n2354_n5888# 0.037984f
C702 source.n518 a_n2354_n5888# 0.017016f
C703 source.n519 a_n2354_n5888# 0.01607f
C704 source.n520 a_n2354_n5888# 0.029906f
C705 source.n521 a_n2354_n5888# 0.029906f
C706 source.n522 a_n2354_n5888# 0.01607f
C707 source.n523 a_n2354_n5888# 0.017016f
C708 source.n524 a_n2354_n5888# 0.037984f
C709 source.n525 a_n2354_n5888# 0.037984f
C710 source.n526 a_n2354_n5888# 0.017016f
C711 source.n527 a_n2354_n5888# 0.01607f
C712 source.n528 a_n2354_n5888# 0.029906f
C713 source.n529 a_n2354_n5888# 0.029906f
C714 source.n530 a_n2354_n5888# 0.01607f
C715 source.n531 a_n2354_n5888# 0.017016f
C716 source.n532 a_n2354_n5888# 0.037984f
C717 source.n533 a_n2354_n5888# 0.037984f
C718 source.n534 a_n2354_n5888# 0.017016f
C719 source.n535 a_n2354_n5888# 0.01607f
C720 source.n536 a_n2354_n5888# 0.029906f
C721 source.n537 a_n2354_n5888# 0.029906f
C722 source.n538 a_n2354_n5888# 0.01607f
C723 source.n539 a_n2354_n5888# 0.017016f
C724 source.n540 a_n2354_n5888# 0.037984f
C725 source.n541 a_n2354_n5888# 0.037984f
C726 source.n542 a_n2354_n5888# 0.017016f
C727 source.n543 a_n2354_n5888# 0.01607f
C728 source.n544 a_n2354_n5888# 0.029906f
C729 source.n545 a_n2354_n5888# 0.029906f
C730 source.n546 a_n2354_n5888# 0.01607f
C731 source.n547 a_n2354_n5888# 0.017016f
C732 source.n548 a_n2354_n5888# 0.037984f
C733 source.n549 a_n2354_n5888# 0.037984f
C734 source.n550 a_n2354_n5888# 0.017016f
C735 source.n551 a_n2354_n5888# 0.01607f
C736 source.n552 a_n2354_n5888# 0.029906f
C737 source.n553 a_n2354_n5888# 0.029906f
C738 source.n554 a_n2354_n5888# 0.01607f
C739 source.n555 a_n2354_n5888# 0.016543f
C740 source.n556 a_n2354_n5888# 0.016543f
C741 source.n557 a_n2354_n5888# 0.037984f
C742 source.n558 a_n2354_n5888# 0.037984f
C743 source.n559 a_n2354_n5888# 0.017016f
C744 source.n560 a_n2354_n5888# 0.01607f
C745 source.n561 a_n2354_n5888# 0.029906f
C746 source.n562 a_n2354_n5888# 0.029906f
C747 source.n563 a_n2354_n5888# 0.01607f
C748 source.n564 a_n2354_n5888# 0.017016f
C749 source.n565 a_n2354_n5888# 0.037984f
C750 source.n566 a_n2354_n5888# 0.037984f
C751 source.n567 a_n2354_n5888# 0.017016f
C752 source.n568 a_n2354_n5888# 0.01607f
C753 source.n569 a_n2354_n5888# 0.029906f
C754 source.n570 a_n2354_n5888# 0.029906f
C755 source.n571 a_n2354_n5888# 0.01607f
C756 source.n572 a_n2354_n5888# 0.017016f
C757 source.n573 a_n2354_n5888# 0.037984f
C758 source.n574 a_n2354_n5888# 0.080802f
C759 source.n575 a_n2354_n5888# 0.017016f
C760 source.n576 a_n2354_n5888# 0.01607f
C761 source.n577 a_n2354_n5888# 0.065858f
C762 source.n578 a_n2354_n5888# 0.044963f
C763 source.n579 a_n2354_n5888# 2.90365f
C764 source.n580 a_n2354_n5888# 0.041229f
C765 source.n581 a_n2354_n5888# 0.029906f
C766 source.n582 a_n2354_n5888# 0.01607f
C767 source.n583 a_n2354_n5888# 0.037984f
C768 source.n584 a_n2354_n5888# 0.017016f
C769 source.n585 a_n2354_n5888# 0.029906f
C770 source.n586 a_n2354_n5888# 0.01607f
C771 source.n587 a_n2354_n5888# 0.037984f
C772 source.n588 a_n2354_n5888# 0.017016f
C773 source.n589 a_n2354_n5888# 0.029906f
C774 source.n590 a_n2354_n5888# 0.01607f
C775 source.n591 a_n2354_n5888# 0.037984f
C776 source.n592 a_n2354_n5888# 0.017016f
C777 source.n593 a_n2354_n5888# 0.029906f
C778 source.n594 a_n2354_n5888# 0.01607f
C779 source.n595 a_n2354_n5888# 0.037984f
C780 source.n596 a_n2354_n5888# 0.017016f
C781 source.n597 a_n2354_n5888# 0.029906f
C782 source.n598 a_n2354_n5888# 0.01607f
C783 source.n599 a_n2354_n5888# 0.037984f
C784 source.n600 a_n2354_n5888# 0.017016f
C785 source.n601 a_n2354_n5888# 0.029906f
C786 source.n602 a_n2354_n5888# 0.01607f
C787 source.n603 a_n2354_n5888# 0.037984f
C788 source.n604 a_n2354_n5888# 0.017016f
C789 source.n605 a_n2354_n5888# 0.029906f
C790 source.n606 a_n2354_n5888# 0.01607f
C791 source.n607 a_n2354_n5888# 0.037984f
C792 source.n608 a_n2354_n5888# 0.017016f
C793 source.n609 a_n2354_n5888# 0.029906f
C794 source.n610 a_n2354_n5888# 0.01607f
C795 source.n611 a_n2354_n5888# 0.037984f
C796 source.n612 a_n2354_n5888# 0.017016f
C797 source.n613 a_n2354_n5888# 0.029906f
C798 source.n614 a_n2354_n5888# 0.016543f
C799 source.n615 a_n2354_n5888# 0.037984f
C800 source.n616 a_n2354_n5888# 0.017016f
C801 source.n617 a_n2354_n5888# 0.029906f
C802 source.n618 a_n2354_n5888# 0.01607f
C803 source.n619 a_n2354_n5888# 0.037984f
C804 source.n620 a_n2354_n5888# 0.017016f
C805 source.n621 a_n2354_n5888# 0.029906f
C806 source.n622 a_n2354_n5888# 0.01607f
C807 source.n623 a_n2354_n5888# 0.028488f
C808 source.n624 a_n2354_n5888# 0.026852f
C809 source.t44 a_n2354_n5888# 0.066247f
C810 source.n625 a_n2354_n5888# 0.364881f
C811 source.n626 a_n2354_n5888# 3.23796f
C812 source.n627 a_n2354_n5888# 0.01607f
C813 source.n628 a_n2354_n5888# 0.017016f
C814 source.n629 a_n2354_n5888# 0.037984f
C815 source.n630 a_n2354_n5888# 0.037984f
C816 source.n631 a_n2354_n5888# 0.017016f
C817 source.n632 a_n2354_n5888# 0.01607f
C818 source.n633 a_n2354_n5888# 0.029906f
C819 source.n634 a_n2354_n5888# 0.029906f
C820 source.n635 a_n2354_n5888# 0.01607f
C821 source.n636 a_n2354_n5888# 0.017016f
C822 source.n637 a_n2354_n5888# 0.037984f
C823 source.n638 a_n2354_n5888# 0.037984f
C824 source.n639 a_n2354_n5888# 0.017016f
C825 source.n640 a_n2354_n5888# 0.01607f
C826 source.n641 a_n2354_n5888# 0.029906f
C827 source.n642 a_n2354_n5888# 0.029906f
C828 source.n643 a_n2354_n5888# 0.01607f
C829 source.n644 a_n2354_n5888# 0.01607f
C830 source.n645 a_n2354_n5888# 0.017016f
C831 source.n646 a_n2354_n5888# 0.037984f
C832 source.n647 a_n2354_n5888# 0.037984f
C833 source.n648 a_n2354_n5888# 0.037984f
C834 source.n649 a_n2354_n5888# 0.016543f
C835 source.n650 a_n2354_n5888# 0.01607f
C836 source.n651 a_n2354_n5888# 0.029906f
C837 source.n652 a_n2354_n5888# 0.029906f
C838 source.n653 a_n2354_n5888# 0.01607f
C839 source.n654 a_n2354_n5888# 0.017016f
C840 source.n655 a_n2354_n5888# 0.037984f
C841 source.n656 a_n2354_n5888# 0.037984f
C842 source.n657 a_n2354_n5888# 0.017016f
C843 source.n658 a_n2354_n5888# 0.01607f
C844 source.n659 a_n2354_n5888# 0.029906f
C845 source.n660 a_n2354_n5888# 0.029906f
C846 source.n661 a_n2354_n5888# 0.01607f
C847 source.n662 a_n2354_n5888# 0.017016f
C848 source.n663 a_n2354_n5888# 0.037984f
C849 source.n664 a_n2354_n5888# 0.037984f
C850 source.n665 a_n2354_n5888# 0.017016f
C851 source.n666 a_n2354_n5888# 0.01607f
C852 source.n667 a_n2354_n5888# 0.029906f
C853 source.n668 a_n2354_n5888# 0.029906f
C854 source.n669 a_n2354_n5888# 0.01607f
C855 source.n670 a_n2354_n5888# 0.017016f
C856 source.n671 a_n2354_n5888# 0.037984f
C857 source.n672 a_n2354_n5888# 0.037984f
C858 source.n673 a_n2354_n5888# 0.017016f
C859 source.n674 a_n2354_n5888# 0.01607f
C860 source.n675 a_n2354_n5888# 0.029906f
C861 source.n676 a_n2354_n5888# 0.029906f
C862 source.n677 a_n2354_n5888# 0.01607f
C863 source.n678 a_n2354_n5888# 0.017016f
C864 source.n679 a_n2354_n5888# 0.037984f
C865 source.n680 a_n2354_n5888# 0.037984f
C866 source.n681 a_n2354_n5888# 0.017016f
C867 source.n682 a_n2354_n5888# 0.01607f
C868 source.n683 a_n2354_n5888# 0.029906f
C869 source.n684 a_n2354_n5888# 0.029906f
C870 source.n685 a_n2354_n5888# 0.01607f
C871 source.n686 a_n2354_n5888# 0.017016f
C872 source.n687 a_n2354_n5888# 0.037984f
C873 source.n688 a_n2354_n5888# 0.037984f
C874 source.n689 a_n2354_n5888# 0.037984f
C875 source.n690 a_n2354_n5888# 0.017016f
C876 source.n691 a_n2354_n5888# 0.01607f
C877 source.n692 a_n2354_n5888# 0.029906f
C878 source.n693 a_n2354_n5888# 0.029906f
C879 source.n694 a_n2354_n5888# 0.01607f
C880 source.n695 a_n2354_n5888# 0.016543f
C881 source.n696 a_n2354_n5888# 0.016543f
C882 source.n697 a_n2354_n5888# 0.037984f
C883 source.n698 a_n2354_n5888# 0.037984f
C884 source.n699 a_n2354_n5888# 0.017016f
C885 source.n700 a_n2354_n5888# 0.01607f
C886 source.n701 a_n2354_n5888# 0.029906f
C887 source.n702 a_n2354_n5888# 0.029906f
C888 source.n703 a_n2354_n5888# 0.01607f
C889 source.n704 a_n2354_n5888# 0.017016f
C890 source.n705 a_n2354_n5888# 0.037984f
C891 source.n706 a_n2354_n5888# 0.037984f
C892 source.n707 a_n2354_n5888# 0.017016f
C893 source.n708 a_n2354_n5888# 0.01607f
C894 source.n709 a_n2354_n5888# 0.029906f
C895 source.n710 a_n2354_n5888# 0.029906f
C896 source.n711 a_n2354_n5888# 0.01607f
C897 source.n712 a_n2354_n5888# 0.017016f
C898 source.n713 a_n2354_n5888# 0.037984f
C899 source.n714 a_n2354_n5888# 0.080802f
C900 source.n715 a_n2354_n5888# 0.017016f
C901 source.n716 a_n2354_n5888# 0.01607f
C902 source.n717 a_n2354_n5888# 0.065858f
C903 source.n718 a_n2354_n5888# 0.044963f
C904 source.n719 a_n2354_n5888# 2.90365f
C905 source.t35 a_n2354_n5888# 0.59082f
C906 source.t28 a_n2354_n5888# 0.59082f
C907 source.n720 a_n2354_n5888# 5.347f
C908 source.n721 a_n2354_n5888# 0.41486f
C909 source.t43 a_n2354_n5888# 0.59082f
C910 source.t29 a_n2354_n5888# 0.59082f
C911 source.n722 a_n2354_n5888# 5.347f
C912 source.n723 a_n2354_n5888# 0.41486f
C913 source.t40 a_n2354_n5888# 0.59082f
C914 source.t31 a_n2354_n5888# 0.59082f
C915 source.n724 a_n2354_n5888# 5.347f
C916 source.n725 a_n2354_n5888# 0.41486f
C917 source.t41 a_n2354_n5888# 0.59082f
C918 source.t33 a_n2354_n5888# 0.59082f
C919 source.n726 a_n2354_n5888# 5.347f
C920 source.n727 a_n2354_n5888# 0.41486f
C921 source.t24 a_n2354_n5888# 0.59082f
C922 source.t36 a_n2354_n5888# 0.59082f
C923 source.n728 a_n2354_n5888# 5.347f
C924 source.n729 a_n2354_n5888# 0.41486f
C925 source.n730 a_n2354_n5888# 0.041229f
C926 source.n731 a_n2354_n5888# 0.029906f
C927 source.n732 a_n2354_n5888# 0.01607f
C928 source.n733 a_n2354_n5888# 0.037984f
C929 source.n734 a_n2354_n5888# 0.017016f
C930 source.n735 a_n2354_n5888# 0.029906f
C931 source.n736 a_n2354_n5888# 0.01607f
C932 source.n737 a_n2354_n5888# 0.037984f
C933 source.n738 a_n2354_n5888# 0.017016f
C934 source.n739 a_n2354_n5888# 0.029906f
C935 source.n740 a_n2354_n5888# 0.01607f
C936 source.n741 a_n2354_n5888# 0.037984f
C937 source.n742 a_n2354_n5888# 0.017016f
C938 source.n743 a_n2354_n5888# 0.029906f
C939 source.n744 a_n2354_n5888# 0.01607f
C940 source.n745 a_n2354_n5888# 0.037984f
C941 source.n746 a_n2354_n5888# 0.017016f
C942 source.n747 a_n2354_n5888# 0.029906f
C943 source.n748 a_n2354_n5888# 0.01607f
C944 source.n749 a_n2354_n5888# 0.037984f
C945 source.n750 a_n2354_n5888# 0.017016f
C946 source.n751 a_n2354_n5888# 0.029906f
C947 source.n752 a_n2354_n5888# 0.01607f
C948 source.n753 a_n2354_n5888# 0.037984f
C949 source.n754 a_n2354_n5888# 0.017016f
C950 source.n755 a_n2354_n5888# 0.029906f
C951 source.n756 a_n2354_n5888# 0.01607f
C952 source.n757 a_n2354_n5888# 0.037984f
C953 source.n758 a_n2354_n5888# 0.017016f
C954 source.n759 a_n2354_n5888# 0.029906f
C955 source.n760 a_n2354_n5888# 0.01607f
C956 source.n761 a_n2354_n5888# 0.037984f
C957 source.n762 a_n2354_n5888# 0.017016f
C958 source.n763 a_n2354_n5888# 0.029906f
C959 source.n764 a_n2354_n5888# 0.016543f
C960 source.n765 a_n2354_n5888# 0.037984f
C961 source.n766 a_n2354_n5888# 0.017016f
C962 source.n767 a_n2354_n5888# 0.029906f
C963 source.n768 a_n2354_n5888# 0.01607f
C964 source.n769 a_n2354_n5888# 0.037984f
C965 source.n770 a_n2354_n5888# 0.017016f
C966 source.n771 a_n2354_n5888# 0.029906f
C967 source.n772 a_n2354_n5888# 0.01607f
C968 source.n773 a_n2354_n5888# 0.028488f
C969 source.n774 a_n2354_n5888# 0.026852f
C970 source.t25 a_n2354_n5888# 0.066247f
C971 source.n775 a_n2354_n5888# 0.364881f
C972 source.n776 a_n2354_n5888# 3.23796f
C973 source.n777 a_n2354_n5888# 0.01607f
C974 source.n778 a_n2354_n5888# 0.017016f
C975 source.n779 a_n2354_n5888# 0.037984f
C976 source.n780 a_n2354_n5888# 0.037984f
C977 source.n781 a_n2354_n5888# 0.017016f
C978 source.n782 a_n2354_n5888# 0.01607f
C979 source.n783 a_n2354_n5888# 0.029906f
C980 source.n784 a_n2354_n5888# 0.029906f
C981 source.n785 a_n2354_n5888# 0.01607f
C982 source.n786 a_n2354_n5888# 0.017016f
C983 source.n787 a_n2354_n5888# 0.037984f
C984 source.n788 a_n2354_n5888# 0.037984f
C985 source.n789 a_n2354_n5888# 0.017016f
C986 source.n790 a_n2354_n5888# 0.01607f
C987 source.n791 a_n2354_n5888# 0.029906f
C988 source.n792 a_n2354_n5888# 0.029906f
C989 source.n793 a_n2354_n5888# 0.01607f
C990 source.n794 a_n2354_n5888# 0.01607f
C991 source.n795 a_n2354_n5888# 0.017016f
C992 source.n796 a_n2354_n5888# 0.037984f
C993 source.n797 a_n2354_n5888# 0.037984f
C994 source.n798 a_n2354_n5888# 0.037984f
C995 source.n799 a_n2354_n5888# 0.016543f
C996 source.n800 a_n2354_n5888# 0.01607f
C997 source.n801 a_n2354_n5888# 0.029906f
C998 source.n802 a_n2354_n5888# 0.029906f
C999 source.n803 a_n2354_n5888# 0.01607f
C1000 source.n804 a_n2354_n5888# 0.017016f
C1001 source.n805 a_n2354_n5888# 0.037984f
C1002 source.n806 a_n2354_n5888# 0.037984f
C1003 source.n807 a_n2354_n5888# 0.017016f
C1004 source.n808 a_n2354_n5888# 0.01607f
C1005 source.n809 a_n2354_n5888# 0.029906f
C1006 source.n810 a_n2354_n5888# 0.029906f
C1007 source.n811 a_n2354_n5888# 0.01607f
C1008 source.n812 a_n2354_n5888# 0.017016f
C1009 source.n813 a_n2354_n5888# 0.037984f
C1010 source.n814 a_n2354_n5888# 0.037984f
C1011 source.n815 a_n2354_n5888# 0.017016f
C1012 source.n816 a_n2354_n5888# 0.01607f
C1013 source.n817 a_n2354_n5888# 0.029906f
C1014 source.n818 a_n2354_n5888# 0.029906f
C1015 source.n819 a_n2354_n5888# 0.01607f
C1016 source.n820 a_n2354_n5888# 0.017016f
C1017 source.n821 a_n2354_n5888# 0.037984f
C1018 source.n822 a_n2354_n5888# 0.037984f
C1019 source.n823 a_n2354_n5888# 0.017016f
C1020 source.n824 a_n2354_n5888# 0.01607f
C1021 source.n825 a_n2354_n5888# 0.029906f
C1022 source.n826 a_n2354_n5888# 0.029906f
C1023 source.n827 a_n2354_n5888# 0.01607f
C1024 source.n828 a_n2354_n5888# 0.017016f
C1025 source.n829 a_n2354_n5888# 0.037984f
C1026 source.n830 a_n2354_n5888# 0.037984f
C1027 source.n831 a_n2354_n5888# 0.017016f
C1028 source.n832 a_n2354_n5888# 0.01607f
C1029 source.n833 a_n2354_n5888# 0.029906f
C1030 source.n834 a_n2354_n5888# 0.029906f
C1031 source.n835 a_n2354_n5888# 0.01607f
C1032 source.n836 a_n2354_n5888# 0.017016f
C1033 source.n837 a_n2354_n5888# 0.037984f
C1034 source.n838 a_n2354_n5888# 0.037984f
C1035 source.n839 a_n2354_n5888# 0.037984f
C1036 source.n840 a_n2354_n5888# 0.017016f
C1037 source.n841 a_n2354_n5888# 0.01607f
C1038 source.n842 a_n2354_n5888# 0.029906f
C1039 source.n843 a_n2354_n5888# 0.029906f
C1040 source.n844 a_n2354_n5888# 0.01607f
C1041 source.n845 a_n2354_n5888# 0.016543f
C1042 source.n846 a_n2354_n5888# 0.016543f
C1043 source.n847 a_n2354_n5888# 0.037984f
C1044 source.n848 a_n2354_n5888# 0.037984f
C1045 source.n849 a_n2354_n5888# 0.017016f
C1046 source.n850 a_n2354_n5888# 0.01607f
C1047 source.n851 a_n2354_n5888# 0.029906f
C1048 source.n852 a_n2354_n5888# 0.029906f
C1049 source.n853 a_n2354_n5888# 0.01607f
C1050 source.n854 a_n2354_n5888# 0.017016f
C1051 source.n855 a_n2354_n5888# 0.037984f
C1052 source.n856 a_n2354_n5888# 0.037984f
C1053 source.n857 a_n2354_n5888# 0.017016f
C1054 source.n858 a_n2354_n5888# 0.01607f
C1055 source.n859 a_n2354_n5888# 0.029906f
C1056 source.n860 a_n2354_n5888# 0.029906f
C1057 source.n861 a_n2354_n5888# 0.01607f
C1058 source.n862 a_n2354_n5888# 0.017016f
C1059 source.n863 a_n2354_n5888# 0.037984f
C1060 source.n864 a_n2354_n5888# 0.080802f
C1061 source.n865 a_n2354_n5888# 0.017016f
C1062 source.n866 a_n2354_n5888# 0.01607f
C1063 source.n867 a_n2354_n5888# 0.065858f
C1064 source.n868 a_n2354_n5888# 0.044963f
C1065 source.n869 a_n2354_n5888# 0.12131f
C1066 source.n870 a_n2354_n5888# 0.041229f
C1067 source.n871 a_n2354_n5888# 0.029906f
C1068 source.n872 a_n2354_n5888# 0.01607f
C1069 source.n873 a_n2354_n5888# 0.037984f
C1070 source.n874 a_n2354_n5888# 0.017016f
C1071 source.n875 a_n2354_n5888# 0.029906f
C1072 source.n876 a_n2354_n5888# 0.01607f
C1073 source.n877 a_n2354_n5888# 0.037984f
C1074 source.n878 a_n2354_n5888# 0.017016f
C1075 source.n879 a_n2354_n5888# 0.029906f
C1076 source.n880 a_n2354_n5888# 0.01607f
C1077 source.n881 a_n2354_n5888# 0.037984f
C1078 source.n882 a_n2354_n5888# 0.017016f
C1079 source.n883 a_n2354_n5888# 0.029906f
C1080 source.n884 a_n2354_n5888# 0.01607f
C1081 source.n885 a_n2354_n5888# 0.037984f
C1082 source.n886 a_n2354_n5888# 0.017016f
C1083 source.n887 a_n2354_n5888# 0.029906f
C1084 source.n888 a_n2354_n5888# 0.01607f
C1085 source.n889 a_n2354_n5888# 0.037984f
C1086 source.n890 a_n2354_n5888# 0.017016f
C1087 source.n891 a_n2354_n5888# 0.029906f
C1088 source.n892 a_n2354_n5888# 0.01607f
C1089 source.n893 a_n2354_n5888# 0.037984f
C1090 source.n894 a_n2354_n5888# 0.017016f
C1091 source.n895 a_n2354_n5888# 0.029906f
C1092 source.n896 a_n2354_n5888# 0.01607f
C1093 source.n897 a_n2354_n5888# 0.037984f
C1094 source.n898 a_n2354_n5888# 0.017016f
C1095 source.n899 a_n2354_n5888# 0.029906f
C1096 source.n900 a_n2354_n5888# 0.01607f
C1097 source.n901 a_n2354_n5888# 0.037984f
C1098 source.n902 a_n2354_n5888# 0.017016f
C1099 source.n903 a_n2354_n5888# 0.029906f
C1100 source.n904 a_n2354_n5888# 0.016543f
C1101 source.n905 a_n2354_n5888# 0.037984f
C1102 source.n906 a_n2354_n5888# 0.017016f
C1103 source.n907 a_n2354_n5888# 0.029906f
C1104 source.n908 a_n2354_n5888# 0.01607f
C1105 source.n909 a_n2354_n5888# 0.037984f
C1106 source.n910 a_n2354_n5888# 0.017016f
C1107 source.n911 a_n2354_n5888# 0.029906f
C1108 source.n912 a_n2354_n5888# 0.01607f
C1109 source.n913 a_n2354_n5888# 0.028488f
C1110 source.n914 a_n2354_n5888# 0.026852f
C1111 source.t8 a_n2354_n5888# 0.066247f
C1112 source.n915 a_n2354_n5888# 0.364881f
C1113 source.n916 a_n2354_n5888# 3.23796f
C1114 source.n917 a_n2354_n5888# 0.01607f
C1115 source.n918 a_n2354_n5888# 0.017016f
C1116 source.n919 a_n2354_n5888# 0.037984f
C1117 source.n920 a_n2354_n5888# 0.037984f
C1118 source.n921 a_n2354_n5888# 0.017016f
C1119 source.n922 a_n2354_n5888# 0.01607f
C1120 source.n923 a_n2354_n5888# 0.029906f
C1121 source.n924 a_n2354_n5888# 0.029906f
C1122 source.n925 a_n2354_n5888# 0.01607f
C1123 source.n926 a_n2354_n5888# 0.017016f
C1124 source.n927 a_n2354_n5888# 0.037984f
C1125 source.n928 a_n2354_n5888# 0.037984f
C1126 source.n929 a_n2354_n5888# 0.017016f
C1127 source.n930 a_n2354_n5888# 0.01607f
C1128 source.n931 a_n2354_n5888# 0.029906f
C1129 source.n932 a_n2354_n5888# 0.029906f
C1130 source.n933 a_n2354_n5888# 0.01607f
C1131 source.n934 a_n2354_n5888# 0.01607f
C1132 source.n935 a_n2354_n5888# 0.017016f
C1133 source.n936 a_n2354_n5888# 0.037984f
C1134 source.n937 a_n2354_n5888# 0.037984f
C1135 source.n938 a_n2354_n5888# 0.037984f
C1136 source.n939 a_n2354_n5888# 0.016543f
C1137 source.n940 a_n2354_n5888# 0.01607f
C1138 source.n941 a_n2354_n5888# 0.029906f
C1139 source.n942 a_n2354_n5888# 0.029906f
C1140 source.n943 a_n2354_n5888# 0.01607f
C1141 source.n944 a_n2354_n5888# 0.017016f
C1142 source.n945 a_n2354_n5888# 0.037984f
C1143 source.n946 a_n2354_n5888# 0.037984f
C1144 source.n947 a_n2354_n5888# 0.017016f
C1145 source.n948 a_n2354_n5888# 0.01607f
C1146 source.n949 a_n2354_n5888# 0.029906f
C1147 source.n950 a_n2354_n5888# 0.029906f
C1148 source.n951 a_n2354_n5888# 0.01607f
C1149 source.n952 a_n2354_n5888# 0.017016f
C1150 source.n953 a_n2354_n5888# 0.037984f
C1151 source.n954 a_n2354_n5888# 0.037984f
C1152 source.n955 a_n2354_n5888# 0.017016f
C1153 source.n956 a_n2354_n5888# 0.01607f
C1154 source.n957 a_n2354_n5888# 0.029906f
C1155 source.n958 a_n2354_n5888# 0.029906f
C1156 source.n959 a_n2354_n5888# 0.01607f
C1157 source.n960 a_n2354_n5888# 0.017016f
C1158 source.n961 a_n2354_n5888# 0.037984f
C1159 source.n962 a_n2354_n5888# 0.037984f
C1160 source.n963 a_n2354_n5888# 0.017016f
C1161 source.n964 a_n2354_n5888# 0.01607f
C1162 source.n965 a_n2354_n5888# 0.029906f
C1163 source.n966 a_n2354_n5888# 0.029906f
C1164 source.n967 a_n2354_n5888# 0.01607f
C1165 source.n968 a_n2354_n5888# 0.017016f
C1166 source.n969 a_n2354_n5888# 0.037984f
C1167 source.n970 a_n2354_n5888# 0.037984f
C1168 source.n971 a_n2354_n5888# 0.017016f
C1169 source.n972 a_n2354_n5888# 0.01607f
C1170 source.n973 a_n2354_n5888# 0.029906f
C1171 source.n974 a_n2354_n5888# 0.029906f
C1172 source.n975 a_n2354_n5888# 0.01607f
C1173 source.n976 a_n2354_n5888# 0.017016f
C1174 source.n977 a_n2354_n5888# 0.037984f
C1175 source.n978 a_n2354_n5888# 0.037984f
C1176 source.n979 a_n2354_n5888# 0.037984f
C1177 source.n980 a_n2354_n5888# 0.017016f
C1178 source.n981 a_n2354_n5888# 0.01607f
C1179 source.n982 a_n2354_n5888# 0.029906f
C1180 source.n983 a_n2354_n5888# 0.029906f
C1181 source.n984 a_n2354_n5888# 0.01607f
C1182 source.n985 a_n2354_n5888# 0.016543f
C1183 source.n986 a_n2354_n5888# 0.016543f
C1184 source.n987 a_n2354_n5888# 0.037984f
C1185 source.n988 a_n2354_n5888# 0.037984f
C1186 source.n989 a_n2354_n5888# 0.017016f
C1187 source.n990 a_n2354_n5888# 0.01607f
C1188 source.n991 a_n2354_n5888# 0.029906f
C1189 source.n992 a_n2354_n5888# 0.029906f
C1190 source.n993 a_n2354_n5888# 0.01607f
C1191 source.n994 a_n2354_n5888# 0.017016f
C1192 source.n995 a_n2354_n5888# 0.037984f
C1193 source.n996 a_n2354_n5888# 0.037984f
C1194 source.n997 a_n2354_n5888# 0.017016f
C1195 source.n998 a_n2354_n5888# 0.01607f
C1196 source.n999 a_n2354_n5888# 0.029906f
C1197 source.n1000 a_n2354_n5888# 0.029906f
C1198 source.n1001 a_n2354_n5888# 0.01607f
C1199 source.n1002 a_n2354_n5888# 0.017016f
C1200 source.n1003 a_n2354_n5888# 0.037984f
C1201 source.n1004 a_n2354_n5888# 0.080802f
C1202 source.n1005 a_n2354_n5888# 0.017016f
C1203 source.n1006 a_n2354_n5888# 0.01607f
C1204 source.n1007 a_n2354_n5888# 0.065858f
C1205 source.n1008 a_n2354_n5888# 0.044963f
C1206 source.n1009 a_n2354_n5888# 0.12131f
C1207 source.t11 a_n2354_n5888# 0.59082f
C1208 source.t14 a_n2354_n5888# 0.59082f
C1209 source.n1010 a_n2354_n5888# 5.347f
C1210 source.n1011 a_n2354_n5888# 0.41486f
C1211 source.t9 a_n2354_n5888# 0.59082f
C1212 source.t12 a_n2354_n5888# 0.59082f
C1213 source.n1012 a_n2354_n5888# 5.347f
C1214 source.n1013 a_n2354_n5888# 0.41486f
C1215 source.t4 a_n2354_n5888# 0.59082f
C1216 source.t7 a_n2354_n5888# 0.59082f
C1217 source.n1014 a_n2354_n5888# 5.347f
C1218 source.n1015 a_n2354_n5888# 0.41486f
C1219 source.t18 a_n2354_n5888# 0.59082f
C1220 source.t3 a_n2354_n5888# 0.59082f
C1221 source.n1016 a_n2354_n5888# 5.347f
C1222 source.n1017 a_n2354_n5888# 0.41486f
C1223 source.t19 a_n2354_n5888# 0.59082f
C1224 source.t21 a_n2354_n5888# 0.59082f
C1225 source.n1018 a_n2354_n5888# 5.347f
C1226 source.n1019 a_n2354_n5888# 0.41486f
C1227 source.n1020 a_n2354_n5888# 0.041229f
C1228 source.n1021 a_n2354_n5888# 0.029906f
C1229 source.n1022 a_n2354_n5888# 0.01607f
C1230 source.n1023 a_n2354_n5888# 0.037984f
C1231 source.n1024 a_n2354_n5888# 0.017016f
C1232 source.n1025 a_n2354_n5888# 0.029906f
C1233 source.n1026 a_n2354_n5888# 0.01607f
C1234 source.n1027 a_n2354_n5888# 0.037984f
C1235 source.n1028 a_n2354_n5888# 0.017016f
C1236 source.n1029 a_n2354_n5888# 0.029906f
C1237 source.n1030 a_n2354_n5888# 0.01607f
C1238 source.n1031 a_n2354_n5888# 0.037984f
C1239 source.n1032 a_n2354_n5888# 0.017016f
C1240 source.n1033 a_n2354_n5888# 0.029906f
C1241 source.n1034 a_n2354_n5888# 0.01607f
C1242 source.n1035 a_n2354_n5888# 0.037984f
C1243 source.n1036 a_n2354_n5888# 0.017016f
C1244 source.n1037 a_n2354_n5888# 0.029906f
C1245 source.n1038 a_n2354_n5888# 0.01607f
C1246 source.n1039 a_n2354_n5888# 0.037984f
C1247 source.n1040 a_n2354_n5888# 0.017016f
C1248 source.n1041 a_n2354_n5888# 0.029906f
C1249 source.n1042 a_n2354_n5888# 0.01607f
C1250 source.n1043 a_n2354_n5888# 0.037984f
C1251 source.n1044 a_n2354_n5888# 0.017016f
C1252 source.n1045 a_n2354_n5888# 0.029906f
C1253 source.n1046 a_n2354_n5888# 0.01607f
C1254 source.n1047 a_n2354_n5888# 0.037984f
C1255 source.n1048 a_n2354_n5888# 0.017016f
C1256 source.n1049 a_n2354_n5888# 0.029906f
C1257 source.n1050 a_n2354_n5888# 0.01607f
C1258 source.n1051 a_n2354_n5888# 0.037984f
C1259 source.n1052 a_n2354_n5888# 0.017016f
C1260 source.n1053 a_n2354_n5888# 0.029906f
C1261 source.n1054 a_n2354_n5888# 0.016543f
C1262 source.n1055 a_n2354_n5888# 0.037984f
C1263 source.n1056 a_n2354_n5888# 0.017016f
C1264 source.n1057 a_n2354_n5888# 0.029906f
C1265 source.n1058 a_n2354_n5888# 0.01607f
C1266 source.n1059 a_n2354_n5888# 0.037984f
C1267 source.n1060 a_n2354_n5888# 0.017016f
C1268 source.n1061 a_n2354_n5888# 0.029906f
C1269 source.n1062 a_n2354_n5888# 0.01607f
C1270 source.n1063 a_n2354_n5888# 0.028488f
C1271 source.n1064 a_n2354_n5888# 0.026852f
C1272 source.t23 a_n2354_n5888# 0.066247f
C1273 source.n1065 a_n2354_n5888# 0.364881f
C1274 source.n1066 a_n2354_n5888# 3.23796f
C1275 source.n1067 a_n2354_n5888# 0.01607f
C1276 source.n1068 a_n2354_n5888# 0.017016f
C1277 source.n1069 a_n2354_n5888# 0.037984f
C1278 source.n1070 a_n2354_n5888# 0.037984f
C1279 source.n1071 a_n2354_n5888# 0.017016f
C1280 source.n1072 a_n2354_n5888# 0.01607f
C1281 source.n1073 a_n2354_n5888# 0.029906f
C1282 source.n1074 a_n2354_n5888# 0.029906f
C1283 source.n1075 a_n2354_n5888# 0.01607f
C1284 source.n1076 a_n2354_n5888# 0.017016f
C1285 source.n1077 a_n2354_n5888# 0.037984f
C1286 source.n1078 a_n2354_n5888# 0.037984f
C1287 source.n1079 a_n2354_n5888# 0.017016f
C1288 source.n1080 a_n2354_n5888# 0.01607f
C1289 source.n1081 a_n2354_n5888# 0.029906f
C1290 source.n1082 a_n2354_n5888# 0.029906f
C1291 source.n1083 a_n2354_n5888# 0.01607f
C1292 source.n1084 a_n2354_n5888# 0.01607f
C1293 source.n1085 a_n2354_n5888# 0.017016f
C1294 source.n1086 a_n2354_n5888# 0.037984f
C1295 source.n1087 a_n2354_n5888# 0.037984f
C1296 source.n1088 a_n2354_n5888# 0.037984f
C1297 source.n1089 a_n2354_n5888# 0.016543f
C1298 source.n1090 a_n2354_n5888# 0.01607f
C1299 source.n1091 a_n2354_n5888# 0.029906f
C1300 source.n1092 a_n2354_n5888# 0.029906f
C1301 source.n1093 a_n2354_n5888# 0.01607f
C1302 source.n1094 a_n2354_n5888# 0.017016f
C1303 source.n1095 a_n2354_n5888# 0.037984f
C1304 source.n1096 a_n2354_n5888# 0.037984f
C1305 source.n1097 a_n2354_n5888# 0.017016f
C1306 source.n1098 a_n2354_n5888# 0.01607f
C1307 source.n1099 a_n2354_n5888# 0.029906f
C1308 source.n1100 a_n2354_n5888# 0.029906f
C1309 source.n1101 a_n2354_n5888# 0.01607f
C1310 source.n1102 a_n2354_n5888# 0.017016f
C1311 source.n1103 a_n2354_n5888# 0.037984f
C1312 source.n1104 a_n2354_n5888# 0.037984f
C1313 source.n1105 a_n2354_n5888# 0.017016f
C1314 source.n1106 a_n2354_n5888# 0.01607f
C1315 source.n1107 a_n2354_n5888# 0.029906f
C1316 source.n1108 a_n2354_n5888# 0.029906f
C1317 source.n1109 a_n2354_n5888# 0.01607f
C1318 source.n1110 a_n2354_n5888# 0.017016f
C1319 source.n1111 a_n2354_n5888# 0.037984f
C1320 source.n1112 a_n2354_n5888# 0.037984f
C1321 source.n1113 a_n2354_n5888# 0.017016f
C1322 source.n1114 a_n2354_n5888# 0.01607f
C1323 source.n1115 a_n2354_n5888# 0.029906f
C1324 source.n1116 a_n2354_n5888# 0.029906f
C1325 source.n1117 a_n2354_n5888# 0.01607f
C1326 source.n1118 a_n2354_n5888# 0.017016f
C1327 source.n1119 a_n2354_n5888# 0.037984f
C1328 source.n1120 a_n2354_n5888# 0.037984f
C1329 source.n1121 a_n2354_n5888# 0.017016f
C1330 source.n1122 a_n2354_n5888# 0.01607f
C1331 source.n1123 a_n2354_n5888# 0.029906f
C1332 source.n1124 a_n2354_n5888# 0.029906f
C1333 source.n1125 a_n2354_n5888# 0.01607f
C1334 source.n1126 a_n2354_n5888# 0.017016f
C1335 source.n1127 a_n2354_n5888# 0.037984f
C1336 source.n1128 a_n2354_n5888# 0.037984f
C1337 source.n1129 a_n2354_n5888# 0.037984f
C1338 source.n1130 a_n2354_n5888# 0.017016f
C1339 source.n1131 a_n2354_n5888# 0.01607f
C1340 source.n1132 a_n2354_n5888# 0.029906f
C1341 source.n1133 a_n2354_n5888# 0.029906f
C1342 source.n1134 a_n2354_n5888# 0.01607f
C1343 source.n1135 a_n2354_n5888# 0.016543f
C1344 source.n1136 a_n2354_n5888# 0.016543f
C1345 source.n1137 a_n2354_n5888# 0.037984f
C1346 source.n1138 a_n2354_n5888# 0.037984f
C1347 source.n1139 a_n2354_n5888# 0.017016f
C1348 source.n1140 a_n2354_n5888# 0.01607f
C1349 source.n1141 a_n2354_n5888# 0.029906f
C1350 source.n1142 a_n2354_n5888# 0.029906f
C1351 source.n1143 a_n2354_n5888# 0.01607f
C1352 source.n1144 a_n2354_n5888# 0.017016f
C1353 source.n1145 a_n2354_n5888# 0.037984f
C1354 source.n1146 a_n2354_n5888# 0.037984f
C1355 source.n1147 a_n2354_n5888# 0.017016f
C1356 source.n1148 a_n2354_n5888# 0.01607f
C1357 source.n1149 a_n2354_n5888# 0.029906f
C1358 source.n1150 a_n2354_n5888# 0.029906f
C1359 source.n1151 a_n2354_n5888# 0.01607f
C1360 source.n1152 a_n2354_n5888# 0.017016f
C1361 source.n1153 a_n2354_n5888# 0.037984f
C1362 source.n1154 a_n2354_n5888# 0.080802f
C1363 source.n1155 a_n2354_n5888# 0.017016f
C1364 source.n1156 a_n2354_n5888# 0.01607f
C1365 source.n1157 a_n2354_n5888# 0.065858f
C1366 source.n1158 a_n2354_n5888# 0.044963f
C1367 source.n1159 a_n2354_n5888# 0.290131f
C1368 source.n1160 a_n2354_n5888# 3.18804f
C1369 drain_left.t5 a_n2354_n5888# 0.683269f
C1370 drain_left.t8 a_n2354_n5888# 0.683269f
C1371 drain_left.n0 a_n2354_n5888# 6.30098f
C1372 drain_left.t22 a_n2354_n5888# 0.683269f
C1373 drain_left.t4 a_n2354_n5888# 0.683269f
C1374 drain_left.n1 a_n2354_n5888# 6.29706f
C1375 drain_left.n2 a_n2354_n5888# 0.836816f
C1376 drain_left.t23 a_n2354_n5888# 0.683269f
C1377 drain_left.t19 a_n2354_n5888# 0.683269f
C1378 drain_left.n3 a_n2354_n5888# 6.29706f
C1379 drain_left.n4 a_n2354_n5888# 0.380679f
C1380 drain_left.t9 a_n2354_n5888# 0.683269f
C1381 drain_left.t16 a_n2354_n5888# 0.683269f
C1382 drain_left.n5 a_n2354_n5888# 6.30098f
C1383 drain_left.t6 a_n2354_n5888# 0.683269f
C1384 drain_left.t15 a_n2354_n5888# 0.683269f
C1385 drain_left.n6 a_n2354_n5888# 6.29706f
C1386 drain_left.n7 a_n2354_n5888# 0.836816f
C1387 drain_left.t13 a_n2354_n5888# 0.683269f
C1388 drain_left.t20 a_n2354_n5888# 0.683269f
C1389 drain_left.n8 a_n2354_n5888# 6.29706f
C1390 drain_left.n9 a_n2354_n5888# 0.380679f
C1391 drain_left.n10 a_n2354_n5888# 3.00897f
C1392 drain_left.t0 a_n2354_n5888# 0.683269f
C1393 drain_left.t11 a_n2354_n5888# 0.683269f
C1394 drain_left.n11 a_n2354_n5888# 6.30098f
C1395 drain_left.t14 a_n2354_n5888# 0.683269f
C1396 drain_left.t17 a_n2354_n5888# 0.683269f
C1397 drain_left.n12 a_n2354_n5888# 6.29706f
C1398 drain_left.n13 a_n2354_n5888# 0.836812f
C1399 drain_left.t18 a_n2354_n5888# 0.683269f
C1400 drain_left.t7 a_n2354_n5888# 0.683269f
C1401 drain_left.n14 a_n2354_n5888# 6.29706f
C1402 drain_left.n15 a_n2354_n5888# 0.413399f
C1403 drain_left.t21 a_n2354_n5888# 0.683269f
C1404 drain_left.t1 a_n2354_n5888# 0.683269f
C1405 drain_left.n16 a_n2354_n5888# 6.29706f
C1406 drain_left.n17 a_n2354_n5888# 0.413399f
C1407 drain_left.t10 a_n2354_n5888# 0.683269f
C1408 drain_left.t12 a_n2354_n5888# 0.683269f
C1409 drain_left.n18 a_n2354_n5888# 6.29706f
C1410 drain_left.n19 a_n2354_n5888# 0.413399f
C1411 drain_left.t2 a_n2354_n5888# 0.683269f
C1412 drain_left.t3 a_n2354_n5888# 0.683269f
C1413 drain_left.n20 a_n2354_n5888# 6.29704f
C1414 drain_left.n21 a_n2354_n5888# 0.701294f
C1415 plus.n0 a_n2354_n5888# 0.049091f
C1416 plus.t0 a_n2354_n5888# 1.03595f
C1417 plus.t17 a_n2354_n5888# 1.03595f
C1418 plus.n1 a_n2354_n5888# 0.376961f
C1419 plus.n2 a_n2354_n5888# 0.049091f
C1420 plus.t10 a_n2354_n5888# 1.03595f
C1421 plus.t1 a_n2354_n5888# 1.03595f
C1422 plus.t20 a_n2354_n5888# 1.03595f
C1423 plus.n3 a_n2354_n5888# 0.376961f
C1424 plus.n4 a_n2354_n5888# 0.049091f
C1425 plus.t13 a_n2354_n5888# 1.03595f
C1426 plus.t8 a_n2354_n5888# 1.03595f
C1427 plus.n5 a_n2354_n5888# 0.376961f
C1428 plus.n6 a_n2354_n5888# 0.049091f
C1429 plus.t21 a_n2354_n5888# 1.03595f
C1430 plus.t15 a_n2354_n5888# 1.03595f
C1431 plus.n7 a_n2354_n5888# 0.018858f
C1432 plus.t2 a_n2354_n5888# 1.04148f
C1433 plus.t9 a_n2354_n5888# 1.03595f
C1434 plus.n8 a_n2354_n5888# 0.376961f
C1435 plus.n9 a_n2354_n5888# 0.392173f
C1436 plus.n10 a_n2354_n5888# 0.105078f
C1437 plus.n11 a_n2354_n5888# 0.049091f
C1438 plus.n12 a_n2354_n5888# 0.017647f
C1439 plus.n13 a_n2354_n5888# 0.376961f
C1440 plus.n14 a_n2354_n5888# 0.02022f
C1441 plus.n15 a_n2354_n5888# 0.376961f
C1442 plus.n16 a_n2354_n5888# 0.02022f
C1443 plus.n17 a_n2354_n5888# 0.049091f
C1444 plus.n18 a_n2354_n5888# 0.049091f
C1445 plus.n19 a_n2354_n5888# 0.02022f
C1446 plus.n20 a_n2354_n5888# 0.376961f
C1447 plus.n21 a_n2354_n5888# 0.018253f
C1448 plus.n22 a_n2354_n5888# 0.018253f
C1449 plus.n23 a_n2354_n5888# 0.049091f
C1450 plus.n24 a_n2354_n5888# 0.049091f
C1451 plus.n25 a_n2354_n5888# 0.02022f
C1452 plus.n26 a_n2354_n5888# 0.376961f
C1453 plus.n27 a_n2354_n5888# 0.02022f
C1454 plus.n28 a_n2354_n5888# 0.376961f
C1455 plus.n29 a_n2354_n5888# 0.02022f
C1456 plus.n30 a_n2354_n5888# 0.049091f
C1457 plus.n31 a_n2354_n5888# 0.049091f
C1458 plus.n32 a_n2354_n5888# 0.017647f
C1459 plus.n33 a_n2354_n5888# 0.018858f
C1460 plus.n34 a_n2354_n5888# 0.376961f
C1461 plus.t5 a_n2354_n5888# 1.04148f
C1462 plus.n35 a_n2354_n5888# 0.392107f
C1463 plus.n36 a_n2354_n5888# 0.873017f
C1464 plus.n37 a_n2354_n5888# 0.049091f
C1465 plus.t3 a_n2354_n5888# 1.04148f
C1466 plus.t12 a_n2354_n5888# 1.03595f
C1467 plus.t19 a_n2354_n5888# 1.03595f
C1468 plus.n38 a_n2354_n5888# 0.376961f
C1469 plus.n39 a_n2354_n5888# 0.049091f
C1470 plus.t4 a_n2354_n5888# 1.03595f
C1471 plus.t18 a_n2354_n5888# 1.03595f
C1472 plus.t7 a_n2354_n5888# 1.03595f
C1473 plus.n40 a_n2354_n5888# 0.376961f
C1474 plus.n41 a_n2354_n5888# 0.049091f
C1475 plus.t16 a_n2354_n5888# 1.03595f
C1476 plus.t6 a_n2354_n5888# 1.03595f
C1477 plus.n42 a_n2354_n5888# 0.376961f
C1478 plus.n43 a_n2354_n5888# 0.049091f
C1479 plus.t14 a_n2354_n5888# 1.03595f
C1480 plus.t23 a_n2354_n5888# 1.03595f
C1481 plus.n44 a_n2354_n5888# 0.018858f
C1482 plus.t11 a_n2354_n5888# 1.03595f
C1483 plus.n45 a_n2354_n5888# 0.376961f
C1484 plus.t22 a_n2354_n5888# 1.04148f
C1485 plus.n46 a_n2354_n5888# 0.392173f
C1486 plus.n47 a_n2354_n5888# 0.105078f
C1487 plus.n48 a_n2354_n5888# 0.049091f
C1488 plus.n49 a_n2354_n5888# 0.017647f
C1489 plus.n50 a_n2354_n5888# 0.376961f
C1490 plus.n51 a_n2354_n5888# 0.02022f
C1491 plus.n52 a_n2354_n5888# 0.376961f
C1492 plus.n53 a_n2354_n5888# 0.02022f
C1493 plus.n54 a_n2354_n5888# 0.049091f
C1494 plus.n55 a_n2354_n5888# 0.049091f
C1495 plus.n56 a_n2354_n5888# 0.02022f
C1496 plus.n57 a_n2354_n5888# 0.376961f
C1497 plus.n58 a_n2354_n5888# 0.018253f
C1498 plus.n59 a_n2354_n5888# 0.018253f
C1499 plus.n60 a_n2354_n5888# 0.049091f
C1500 plus.n61 a_n2354_n5888# 0.049091f
C1501 plus.n62 a_n2354_n5888# 0.02022f
C1502 plus.n63 a_n2354_n5888# 0.376961f
C1503 plus.n64 a_n2354_n5888# 0.02022f
C1504 plus.n65 a_n2354_n5888# 0.376961f
C1505 plus.n66 a_n2354_n5888# 0.02022f
C1506 plus.n67 a_n2354_n5888# 0.049091f
C1507 plus.n68 a_n2354_n5888# 0.049091f
C1508 plus.n69 a_n2354_n5888# 0.017647f
C1509 plus.n70 a_n2354_n5888# 0.018858f
C1510 plus.n71 a_n2354_n5888# 0.376961f
C1511 plus.n72 a_n2354_n5888# 0.392107f
C1512 plus.n73 a_n2354_n5888# 2.02293f
.ends

