* NGSPICE file created from diffpair620.ext - technology: sky130A

.subckt diffpair620 minus drain_right drain_left source plus
X0 drain_right minus source a_n1128_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.7
X1 a_n1128_n4892# a_n1128_n4892# a_n1128_n4892# a_n1128_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.7
X2 a_n1128_n4892# a_n1128_n4892# a_n1128_n4892# a_n1128_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X3 drain_left plus source a_n1128_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.7
X4 drain_left plus source a_n1128_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.7
X5 drain_right minus source a_n1128_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=7.8 ps=40.78 w=20 l=0.7
X6 a_n1128_n4892# a_n1128_n4892# a_n1128_n4892# a_n1128_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X7 a_n1128_n4892# a_n1128_n4892# a_n1128_n4892# a_n1128_n4892# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
.ends

