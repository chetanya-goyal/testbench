* NGSPICE file created from diffpair200.ext - technology: sky130A

.subckt diffpair200 minus drain_right drain_left source plus
X0 drain_right.t1 minus.t0 source.t2 a_n1048_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=0.5
X1 a_n1048_n1492# a_n1048_n1492# a_n1048_n1492# a_n1048_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.5
X2 drain_left.t1 plus.t0 source.t0 a_n1048_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=0.5
X3 a_n1048_n1492# a_n1048_n1492# a_n1048_n1492# a_n1048_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X4 a_n1048_n1492# a_n1048_n1492# a_n1048_n1492# a_n1048_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X5 drain_left.t0 plus.t1 source.t1 a_n1048_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=0.5
X6 a_n1048_n1492# a_n1048_n1492# a_n1048_n1492# a_n1048_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X7 drain_right.t0 minus.t1 source.t3 a_n1048_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=0.5
R0 minus.n0 minus.t0 410.757
R1 minus.n0 minus.t1 390.969
R2 minus minus.n0 0.188
R3 source.n0 source.t0 69.6943
R4 source.n1 source.t2 69.6943
R5 source.n3 source.t3 69.6942
R6 source.n2 source.t1 69.6942
R7 source.n2 source.n1 15.9157
R8 source.n4 source.n0 9.57952
R9 source.n4 source.n3 5.62119
R10 source.n1 source.n0 0.828086
R11 source.n3 source.n2 0.828086
R12 source source.n4 0.188
R13 drain_right drain_right.t0 107.401
R14 drain_right drain_right.t1 92.3836
R15 plus plus.t1 408.046
R16 plus plus.t0 393.204
R17 drain_left drain_left.t0 107.954
R18 drain_left drain_left.t1 92.7413
C0 drain_right plus 0.256691f
C1 source drain_left 2.47561f
C2 source minus 0.5553f
C3 drain_left minus 0.176817f
C4 source plus 0.569441f
C5 drain_right source 2.47199f
C6 drain_left plus 0.714988f
C7 drain_right drain_left 0.440057f
C8 minus plus 2.79144f
C9 drain_right minus 0.619484f
C10 drain_right a_n1048_n1492# 3.62077f
C11 drain_left a_n1048_n1492# 3.73301f
C12 source a_n1048_n1492# 2.554442f
C13 minus a_n1048_n1492# 3.210814f
C14 plus a_n1048_n1492# 5.30685f
C15 drain_left.t0 a_n1048_n1492# 0.475915f
C16 drain_left.t1 a_n1048_n1492# 0.39518f
C17 plus.t0 a_n1048_n1492# 0.246636f
C18 plus.t1 a_n1048_n1492# 0.290258f
C19 drain_right.t0 a_n1048_n1492# 0.47984f
C20 drain_right.t1 a_n1048_n1492# 0.405261f
C21 source.t0 a_n1048_n1492# 0.40839f
C22 source.n0 a_n1048_n1492# 0.585831f
C23 source.t2 a_n1048_n1492# 0.40839f
C24 source.n1 a_n1048_n1492# 0.853106f
C25 source.t1 a_n1048_n1492# 0.408388f
C26 source.n2 a_n1048_n1492# 0.853108f
C27 source.t3 a_n1048_n1492# 0.408388f
C28 source.n3 a_n1048_n1492# 0.431291f
C29 source.n4 a_n1048_n1492# 0.608189f
C30 minus.t0 a_n1048_n1492# 0.289719f
C31 minus.t1 a_n1048_n1492# 0.236493f
C32 minus.n0 a_n1048_n1492# 2.24643f
.ends

