* NGSPICE file created from diffpair450.ext - technology: sky130A

.subckt diffpair450 minus drain_right drain_left source plus
X0 drain_right minus source a_n1088_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.6
X1 drain_left plus source a_n1088_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.6
X2 drain_left plus source a_n1088_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.6
X3 a_n1088_n3292# a_n1088_n3292# a_n1088_n3292# a_n1088_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.6
X4 a_n1088_n3292# a_n1088_n3292# a_n1088_n3292# a_n1088_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.6
X5 a_n1088_n3292# a_n1088_n3292# a_n1088_n3292# a_n1088_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.6
X6 a_n1088_n3292# a_n1088_n3292# a_n1088_n3292# a_n1088_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.6
X7 drain_right minus source a_n1088_n3292# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=4.68 ps=24.78 w=12 l=0.6
.ends

