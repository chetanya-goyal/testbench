* NGSPICE file created from diffpair194.ext - technology: sky130A

.subckt diffpair194 minus drain_right drain_left source plus
X0 source.t15 minus.t0 drain_right.t4 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X1 drain_left.t9 plus.t0 source.t5 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X2 drain_right.t0 minus.t1 source.t14 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X3 a_n1472_n1488# a_n1472_n1488# a_n1472_n1488# a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.3
X4 drain_right.t8 minus.t2 source.t13 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X5 drain_left.t8 plus.t1 source.t1 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X6 a_n1472_n1488# a_n1472_n1488# a_n1472_n1488# a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X7 drain_left.t7 plus.t2 source.t3 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X8 a_n1472_n1488# a_n1472_n1488# a_n1472_n1488# a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X9 drain_right.t1 minus.t3 source.t12 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X10 drain_left.t6 plus.t3 source.t4 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X11 source.t0 plus.t4 drain_left.t5 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X12 source.t2 plus.t5 drain_left.t4 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X13 source.t11 minus.t4 drain_right.t6 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X14 source.t10 minus.t5 drain_right.t2 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X15 a_n1472_n1488# a_n1472_n1488# a_n1472_n1488# a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X16 drain_right.t3 minus.t6 source.t9 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X17 drain_left.t3 plus.t6 source.t16 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X18 drain_left.t2 plus.t7 source.t17 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X19 drain_right.t5 minus.t7 source.t8 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X20 source.t7 minus.t8 drain_right.t9 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X21 drain_right.t7 minus.t9 source.t6 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X22 source.t18 plus.t8 drain_left.t1 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
X23 source.t19 plus.t9 drain_left.t0 a_n1472_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.3
R0 minus.n9 minus.t7 383.409
R1 minus.n3 minus.t6 383.409
R2 minus.n20 minus.t2 383.409
R3 minus.n14 minus.t3 383.409
R4 minus.n6 minus.t1 345.433
R5 minus.n8 minus.t5 345.433
R6 minus.n2 minus.t8 345.433
R7 minus.n17 minus.t9 345.433
R8 minus.n19 minus.t4 345.433
R9 minus.n13 minus.t0 345.433
R10 minus.n4 minus.n3 161.489
R11 minus.n15 minus.n14 161.489
R12 minus.n10 minus.n9 161.3
R13 minus.n7 minus.n0 161.3
R14 minus.n6 minus.n5 161.3
R15 minus.n4 minus.n1 161.3
R16 minus.n21 minus.n20 161.3
R17 minus.n18 minus.n11 161.3
R18 minus.n17 minus.n16 161.3
R19 minus.n15 minus.n12 161.3
R20 minus.n7 minus.n6 73.0308
R21 minus.n6 minus.n1 73.0308
R22 minus.n17 minus.n12 73.0308
R23 minus.n18 minus.n17 73.0308
R24 minus.n9 minus.n8 54.0429
R25 minus.n3 minus.n2 54.0429
R26 minus.n14 minus.n13 54.0429
R27 minus.n20 minus.n19 54.0429
R28 minus.n22 minus.n10 27.866
R29 minus.n8 minus.n7 18.9884
R30 minus.n2 minus.n1 18.9884
R31 minus.n13 minus.n12 18.9884
R32 minus.n19 minus.n18 18.9884
R33 minus.n22 minus.n21 6.48724
R34 minus.n10 minus.n0 0.189894
R35 minus.n5 minus.n0 0.189894
R36 minus.n5 minus.n4 0.189894
R37 minus.n16 minus.n15 0.189894
R38 minus.n16 minus.n11 0.189894
R39 minus.n21 minus.n11 0.189894
R40 minus minus.n22 0.188
R41 drain_right.n1 drain_right.t1 86.9161
R42 drain_right.n7 drain_right.t5 86.3731
R43 drain_right.n6 drain_right.n4 80.3162
R44 drain_right.n3 drain_right.n2 80.125
R45 drain_right.n6 drain_right.n5 79.7731
R46 drain_right.n1 drain_right.n0 79.773
R47 drain_right drain_right.n3 22.3039
R48 drain_right.n2 drain_right.t6 6.6005
R49 drain_right.n2 drain_right.t8 6.6005
R50 drain_right.n0 drain_right.t4 6.6005
R51 drain_right.n0 drain_right.t7 6.6005
R52 drain_right.n4 drain_right.t9 6.6005
R53 drain_right.n4 drain_right.t3 6.6005
R54 drain_right.n5 drain_right.t2 6.6005
R55 drain_right.n5 drain_right.t0 6.6005
R56 drain_right drain_right.n7 5.92477
R57 drain_right.n7 drain_right.n6 0.543603
R58 drain_right.n3 drain_right.n1 0.0809298
R59 source.n0 source.t4 69.6943
R60 source.n5 source.t9 69.6943
R61 source.n19 source.t13 69.6942
R62 source.n14 source.t3 69.6942
R63 source.n2 source.n1 63.0943
R64 source.n4 source.n3 63.0943
R65 source.n7 source.n6 63.0943
R66 source.n9 source.n8 63.0943
R67 source.n18 source.n17 63.0942
R68 source.n16 source.n15 63.0942
R69 source.n13 source.n12 63.0942
R70 source.n11 source.n10 63.0942
R71 source.n11 source.n9 15.5558
R72 source.n20 source.n0 9.47816
R73 source.n17 source.t6 6.6005
R74 source.n17 source.t11 6.6005
R75 source.n15 source.t12 6.6005
R76 source.n15 source.t15 6.6005
R77 source.n12 source.t17 6.6005
R78 source.n12 source.t18 6.6005
R79 source.n10 source.t5 6.6005
R80 source.n10 source.t0 6.6005
R81 source.n1 source.t16 6.6005
R82 source.n1 source.t19 6.6005
R83 source.n3 source.t1 6.6005
R84 source.n3 source.t2 6.6005
R85 source.n6 source.t14 6.6005
R86 source.n6 source.t7 6.6005
R87 source.n8 source.t8 6.6005
R88 source.n8 source.t10 6.6005
R89 source.n20 source.n19 5.53498
R90 source.n5 source.n4 0.741879
R91 source.n16 source.n14 0.741879
R92 source.n9 source.n7 0.543603
R93 source.n7 source.n5 0.543603
R94 source.n4 source.n2 0.543603
R95 source.n2 source.n0 0.543603
R96 source.n13 source.n11 0.543603
R97 source.n14 source.n13 0.543603
R98 source.n18 source.n16 0.543603
R99 source.n19 source.n18 0.543603
R100 source source.n20 0.188
R101 plus.n3 plus.t1 383.409
R102 plus.n9 plus.t3 383.409
R103 plus.n14 plus.t2 383.409
R104 plus.n20 plus.t0 383.409
R105 plus.n6 plus.t6 345.433
R106 plus.n2 plus.t5 345.433
R107 plus.n8 plus.t9 345.433
R108 plus.n17 plus.t7 345.433
R109 plus.n13 plus.t8 345.433
R110 plus.n19 plus.t4 345.433
R111 plus.n4 plus.n3 161.489
R112 plus.n15 plus.n14 161.489
R113 plus.n4 plus.n1 161.3
R114 plus.n6 plus.n5 161.3
R115 plus.n7 plus.n0 161.3
R116 plus.n10 plus.n9 161.3
R117 plus.n15 plus.n12 161.3
R118 plus.n17 plus.n16 161.3
R119 plus.n18 plus.n11 161.3
R120 plus.n21 plus.n20 161.3
R121 plus.n6 plus.n1 73.0308
R122 plus.n7 plus.n6 73.0308
R123 plus.n18 plus.n17 73.0308
R124 plus.n17 plus.n12 73.0308
R125 plus.n3 plus.n2 54.0429
R126 plus.n9 plus.n8 54.0429
R127 plus.n20 plus.n19 54.0429
R128 plus.n14 plus.n13 54.0429
R129 plus plus.n21 25.1562
R130 plus.n2 plus.n1 18.9884
R131 plus.n8 plus.n7 18.9884
R132 plus.n19 plus.n18 18.9884
R133 plus.n13 plus.n12 18.9884
R134 plus plus.n10 8.72209
R135 plus.n5 plus.n4 0.189894
R136 plus.n5 plus.n0 0.189894
R137 plus.n10 plus.n0 0.189894
R138 plus.n21 plus.n11 0.189894
R139 plus.n16 plus.n11 0.189894
R140 plus.n16 plus.n15 0.189894
R141 drain_left.n5 drain_left.t8 86.9162
R142 drain_left.n1 drain_left.t9 86.9161
R143 drain_left.n3 drain_left.n2 80.125
R144 drain_left.n7 drain_left.n6 79.7731
R145 drain_left.n5 drain_left.n4 79.7731
R146 drain_left.n1 drain_left.n0 79.773
R147 drain_left drain_left.n3 22.8571
R148 drain_left.n2 drain_left.t1 6.6005
R149 drain_left.n2 drain_left.t7 6.6005
R150 drain_left.n0 drain_left.t5 6.6005
R151 drain_left.n0 drain_left.t2 6.6005
R152 drain_left.n6 drain_left.t0 6.6005
R153 drain_left.n6 drain_left.t6 6.6005
R154 drain_left.n4 drain_left.t4 6.6005
R155 drain_left.n4 drain_left.t3 6.6005
R156 drain_left drain_left.n7 6.19632
R157 drain_left.n7 drain_left.n5 0.543603
R158 drain_left.n3 drain_left.n1 0.0809298
C0 drain_right source 6.86985f
C1 plus drain_left 1.43365f
C2 drain_right minus 1.29397f
C3 source plus 1.36707f
C4 plus minus 3.32773f
C5 drain_right plus 0.300641f
C6 source drain_left 6.87358f
C7 minus drain_left 0.176413f
C8 drain_right drain_left 0.721115f
C9 source minus 1.3529f
C10 drain_right a_n1472_n1488# 3.83078f
C11 drain_left a_n1472_n1488# 4.04305f
C12 source a_n1472_n1488# 2.807247f
C13 minus a_n1472_n1488# 4.977016f
C14 plus a_n1472_n1488# 5.622816f
C15 drain_left.t9 a_n1472_n1488# 0.522919f
C16 drain_left.t5 a_n1472_n1488# 0.056306f
C17 drain_left.t2 a_n1472_n1488# 0.056306f
C18 drain_left.n0 a_n1472_n1488# 0.406071f
C19 drain_left.n1 a_n1472_n1488# 0.522651f
C20 drain_left.t1 a_n1472_n1488# 0.056306f
C21 drain_left.t7 a_n1472_n1488# 0.056306f
C22 drain_left.n2 a_n1472_n1488# 0.407256f
C23 drain_left.n3 a_n1472_n1488# 0.895828f
C24 drain_left.t8 a_n1472_n1488# 0.522921f
C25 drain_left.t4 a_n1472_n1488# 0.056306f
C26 drain_left.t3 a_n1472_n1488# 0.056306f
C27 drain_left.n4 a_n1472_n1488# 0.406073f
C28 drain_left.n5 a_n1472_n1488# 0.55121f
C29 drain_left.t0 a_n1472_n1488# 0.056306f
C30 drain_left.t6 a_n1472_n1488# 0.056306f
C31 drain_left.n6 a_n1472_n1488# 0.406073f
C32 drain_left.n7 a_n1472_n1488# 0.470939f
C33 plus.n0 a_n1472_n1488# 0.030003f
C34 plus.t9 a_n1472_n1488# 0.078197f
C35 plus.t6 a_n1472_n1488# 0.078197f
C36 plus.n1 a_n1472_n1488# 0.012358f
C37 plus.t1 a_n1472_n1488# 0.082804f
C38 plus.t5 a_n1472_n1488# 0.078197f
C39 plus.n2 a_n1472_n1488# 0.045405f
C40 plus.n3 a_n1472_n1488# 0.054307f
C41 plus.n4 a_n1472_n1488# 0.065884f
C42 plus.n5 a_n1472_n1488# 0.030003f
C43 plus.n6 a_n1472_n1488# 0.055358f
C44 plus.n7 a_n1472_n1488# 0.012358f
C45 plus.n8 a_n1472_n1488# 0.045405f
C46 plus.t3 a_n1472_n1488# 0.082804f
C47 plus.n9 a_n1472_n1488# 0.054265f
C48 plus.n10 a_n1472_n1488# 0.22317f
C49 plus.n11 a_n1472_n1488# 0.030003f
C50 plus.t0 a_n1472_n1488# 0.082804f
C51 plus.t4 a_n1472_n1488# 0.078197f
C52 plus.t7 a_n1472_n1488# 0.078197f
C53 plus.n12 a_n1472_n1488# 0.012358f
C54 plus.t8 a_n1472_n1488# 0.078197f
C55 plus.n13 a_n1472_n1488# 0.045405f
C56 plus.t2 a_n1472_n1488# 0.082804f
C57 plus.n14 a_n1472_n1488# 0.054307f
C58 plus.n15 a_n1472_n1488# 0.065884f
C59 plus.n16 a_n1472_n1488# 0.030003f
C60 plus.n17 a_n1472_n1488# 0.055358f
C61 plus.n18 a_n1472_n1488# 0.012358f
C62 plus.n19 a_n1472_n1488# 0.045405f
C63 plus.n20 a_n1472_n1488# 0.054265f
C64 plus.n21 a_n1472_n1488# 0.647256f
C65 source.t4 a_n1472_n1488# 0.551945f
C66 source.n0 a_n1472_n1488# 0.753038f
C67 source.t16 a_n1472_n1488# 0.066469f
C68 source.t19 a_n1472_n1488# 0.066469f
C69 source.n1 a_n1472_n1488# 0.42145f
C70 source.n2 a_n1472_n1488# 0.342377f
C71 source.t1 a_n1472_n1488# 0.066469f
C72 source.t2 a_n1472_n1488# 0.066469f
C73 source.n3 a_n1472_n1488# 0.42145f
C74 source.n4 a_n1472_n1488# 0.36029f
C75 source.t9 a_n1472_n1488# 0.551945f
C76 source.n5 a_n1472_n1488# 0.411074f
C77 source.t14 a_n1472_n1488# 0.066469f
C78 source.t7 a_n1472_n1488# 0.066469f
C79 source.n6 a_n1472_n1488# 0.42145f
C80 source.n7 a_n1472_n1488# 0.342377f
C81 source.t8 a_n1472_n1488# 0.066469f
C82 source.t10 a_n1472_n1488# 0.066469f
C83 source.n8 a_n1472_n1488# 0.42145f
C84 source.n9 a_n1472_n1488# 1.04358f
C85 source.t5 a_n1472_n1488# 0.066469f
C86 source.t0 a_n1472_n1488# 0.066469f
C87 source.n10 a_n1472_n1488# 0.421447f
C88 source.n11 a_n1472_n1488# 1.04358f
C89 source.t17 a_n1472_n1488# 0.066469f
C90 source.t18 a_n1472_n1488# 0.066469f
C91 source.n12 a_n1472_n1488# 0.421447f
C92 source.n13 a_n1472_n1488# 0.34238f
C93 source.t3 a_n1472_n1488# 0.551942f
C94 source.n14 a_n1472_n1488# 0.411077f
C95 source.t12 a_n1472_n1488# 0.066469f
C96 source.t15 a_n1472_n1488# 0.066469f
C97 source.n15 a_n1472_n1488# 0.421447f
C98 source.n16 a_n1472_n1488# 0.360293f
C99 source.t6 a_n1472_n1488# 0.066469f
C100 source.t11 a_n1472_n1488# 0.066469f
C101 source.n17 a_n1472_n1488# 0.421447f
C102 source.n18 a_n1472_n1488# 0.34238f
C103 source.t13 a_n1472_n1488# 0.551942f
C104 source.n19 a_n1472_n1488# 0.544816f
C105 source.n20 a_n1472_n1488# 0.812678f
C106 drain_right.t1 a_n1472_n1488# 0.530057f
C107 drain_right.t4 a_n1472_n1488# 0.057074f
C108 drain_right.t7 a_n1472_n1488# 0.057074f
C109 drain_right.n0 a_n1472_n1488# 0.411614f
C110 drain_right.n1 a_n1472_n1488# 0.529785f
C111 drain_right.t6 a_n1472_n1488# 0.057074f
C112 drain_right.t8 a_n1472_n1488# 0.057074f
C113 drain_right.n2 a_n1472_n1488# 0.412815f
C114 drain_right.n3 a_n1472_n1488# 0.860127f
C115 drain_right.t9 a_n1472_n1488# 0.057074f
C116 drain_right.t3 a_n1472_n1488# 0.057074f
C117 drain_right.n4 a_n1472_n1488# 0.413554f
C118 drain_right.t2 a_n1472_n1488# 0.057074f
C119 drain_right.t0 a_n1472_n1488# 0.057074f
C120 drain_right.n5 a_n1472_n1488# 0.411616f
C121 drain_right.n6 a_n1472_n1488# 0.561711f
C122 drain_right.t5 a_n1472_n1488# 0.528287f
C123 drain_right.n7 a_n1472_n1488# 0.484373f
C124 minus.n0 a_n1472_n1488# 0.029461f
C125 minus.t7 a_n1472_n1488# 0.081309f
C126 minus.t5 a_n1472_n1488# 0.076785f
C127 minus.t1 a_n1472_n1488# 0.076785f
C128 minus.n1 a_n1472_n1488# 0.012135f
C129 minus.t8 a_n1472_n1488# 0.076785f
C130 minus.n2 a_n1472_n1488# 0.044585f
C131 minus.t6 a_n1472_n1488# 0.081309f
C132 minus.n3 a_n1472_n1488# 0.053327f
C133 minus.n4 a_n1472_n1488# 0.064694f
C134 minus.n5 a_n1472_n1488# 0.029461f
C135 minus.n6 a_n1472_n1488# 0.054358f
C136 minus.n7 a_n1472_n1488# 0.012135f
C137 minus.n8 a_n1472_n1488# 0.044585f
C138 minus.n9 a_n1472_n1488# 0.053285f
C139 minus.n10 a_n1472_n1488# 0.673656f
C140 minus.n11 a_n1472_n1488# 0.029461f
C141 minus.t4 a_n1472_n1488# 0.076785f
C142 minus.t9 a_n1472_n1488# 0.076785f
C143 minus.n12 a_n1472_n1488# 0.012135f
C144 minus.t3 a_n1472_n1488# 0.081309f
C145 minus.t0 a_n1472_n1488# 0.076785f
C146 minus.n13 a_n1472_n1488# 0.044585f
C147 minus.n14 a_n1472_n1488# 0.053327f
C148 minus.n15 a_n1472_n1488# 0.064694f
C149 minus.n16 a_n1472_n1488# 0.029461f
C150 minus.n17 a_n1472_n1488# 0.054358f
C151 minus.n18 a_n1472_n1488# 0.012135f
C152 minus.n19 a_n1472_n1488# 0.044585f
C153 minus.t2 a_n1472_n1488# 0.081309f
C154 minus.n20 a_n1472_n1488# 0.053285f
C155 minus.n21 a_n1472_n1488# 0.191725f
C156 minus.n22 a_n1472_n1488# 0.833271f
.ends

