* NGSPICE file created from diffpair557.ext - technology: sky130A

.subckt diffpair557 minus drain_right drain_left source plus
X0 a_n2750_n3888# a_n2750_n3888# a_n2750_n3888# a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.8
X1 drain_left.t15 plus.t0 source.t24 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X2 source.t5 minus.t0 drain_right.t15 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X3 source.t8 minus.t1 drain_right.t14 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X4 source.t25 plus.t1 drain_left.t14 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X5 a_n2750_n3888# a_n2750_n3888# a_n2750_n3888# a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X6 drain_right.t13 minus.t2 source.t9 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X7 source.t18 plus.t2 drain_left.t13 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X8 drain_right.t12 minus.t3 source.t1 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X9 drain_right.t11 minus.t4 source.t2 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X10 drain_right.t10 minus.t5 source.t10 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X11 source.t29 plus.t3 drain_left.t12 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X12 source.t13 minus.t6 drain_right.t9 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X13 drain_right.t8 minus.t7 source.t6 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X14 source.t21 plus.t4 drain_left.t11 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X15 drain_right.t7 minus.t8 source.t12 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X16 source.t11 minus.t9 drain_right.t6 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X17 drain_right.t5 minus.t10 source.t4 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X18 drain_left.t10 plus.t5 source.t15 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X19 a_n2750_n3888# a_n2750_n3888# a_n2750_n3888# a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X20 drain_left.t9 plus.t6 source.t16 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X21 source.t31 minus.t11 drain_right.t4 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X22 drain_right.t3 minus.t12 source.t0 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X23 source.t19 plus.t7 drain_left.t8 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X24 drain_left.t7 plus.t8 source.t17 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X25 drain_left.t6 plus.t9 source.t28 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X26 source.t3 minus.t13 drain_right.t2 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X27 source.t26 plus.t10 drain_left.t5 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X28 drain_left.t4 plus.t11 source.t14 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X29 source.t22 plus.t12 drain_left.t3 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X30 drain_left.t2 plus.t13 source.t27 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X31 drain_left.t1 plus.t14 source.t23 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X32 a_n2750_n3888# a_n2750_n3888# a_n2750_n3888# a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X33 source.t7 minus.t14 drain_right.t1 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X34 source.t20 plus.t15 drain_left.t0 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X35 source.t30 minus.t15 drain_right.t0 a_n2750_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
R0 plus.n7 plus.t15 522.003
R1 plus.n29 plus.t0 522.003
R2 plus.n20 plus.t6 500.979
R3 plus.n18 plus.t7 500.979
R4 plus.n17 plus.t8 500.979
R5 plus.n3 plus.t12 500.979
R6 plus.n11 plus.t9 500.979
R7 plus.n5 plus.t10 500.979
R8 plus.n6 plus.t13 500.979
R9 plus.n42 plus.t2 500.979
R10 plus.n40 plus.t5 500.979
R11 plus.n39 plus.t1 500.979
R12 plus.n25 plus.t11 500.979
R13 plus.n33 plus.t3 500.979
R14 plus.n27 plus.t14 500.979
R15 plus.n28 plus.t4 500.979
R16 plus.n10 plus.n9 161.3
R17 plus.n11 plus.n4 161.3
R18 plus.n13 plus.n12 161.3
R19 plus.n14 plus.n3 161.3
R20 plus.n16 plus.n15 161.3
R21 plus.n19 plus.n0 161.3
R22 plus.n21 plus.n20 161.3
R23 plus.n32 plus.n31 161.3
R24 plus.n33 plus.n26 161.3
R25 plus.n35 plus.n34 161.3
R26 plus.n36 plus.n25 161.3
R27 plus.n38 plus.n37 161.3
R28 plus.n41 plus.n22 161.3
R29 plus.n43 plus.n42 161.3
R30 plus.n8 plus.n5 80.6037
R31 plus.n17 plus.n2 80.6037
R32 plus.n18 plus.n1 80.6037
R33 plus.n30 plus.n27 80.6037
R34 plus.n39 plus.n24 80.6037
R35 plus.n40 plus.n23 80.6037
R36 plus.n18 plus.n17 48.2005
R37 plus.n6 plus.n5 48.2005
R38 plus.n40 plus.n39 48.2005
R39 plus.n28 plus.n27 48.2005
R40 plus.n17 plus.n16 43.0884
R41 plus.n10 plus.n5 43.0884
R42 plus.n39 plus.n38 43.0884
R43 plus.n32 plus.n27 43.0884
R44 plus.n19 plus.n18 40.1672
R45 plus.n41 plus.n40 40.1672
R46 plus plus.n43 34.7111
R47 plus.n8 plus.n7 31.6481
R48 plus.n30 plus.n29 31.6481
R49 plus.n12 plus.n11 24.1005
R50 plus.n12 plus.n3 24.1005
R51 plus.n34 plus.n25 24.1005
R52 plus.n34 plus.n33 24.1005
R53 plus.n7 plus.n6 17.444
R54 plus.n29 plus.n28 17.444
R55 plus plus.n21 13.4361
R56 plus.n20 plus.n19 8.03383
R57 plus.n42 plus.n41 8.03383
R58 plus.n16 plus.n3 5.11262
R59 plus.n11 plus.n10 5.11262
R60 plus.n38 plus.n25 5.11262
R61 plus.n33 plus.n32 5.11262
R62 plus.n2 plus.n1 0.380177
R63 plus.n24 plus.n23 0.380177
R64 plus.n9 plus.n8 0.285035
R65 plus.n15 plus.n2 0.285035
R66 plus.n1 plus.n0 0.285035
R67 plus.n23 plus.n22 0.285035
R68 plus.n37 plus.n24 0.285035
R69 plus.n31 plus.n30 0.285035
R70 plus.n9 plus.n4 0.189894
R71 plus.n13 plus.n4 0.189894
R72 plus.n14 plus.n13 0.189894
R73 plus.n15 plus.n14 0.189894
R74 plus.n21 plus.n0 0.189894
R75 plus.n43 plus.n22 0.189894
R76 plus.n37 plus.n36 0.189894
R77 plus.n36 plus.n35 0.189894
R78 plus.n35 plus.n26 0.189894
R79 plus.n31 plus.n26 0.189894
R80 source.n7 source.t20 45.521
R81 source.n8 source.t12 45.521
R82 source.n15 source.t3 45.521
R83 source.n31 source.t9 45.5208
R84 source.n24 source.t8 45.5208
R85 source.n23 source.t24 45.5208
R86 source.n16 source.t18 45.5208
R87 source.n0 source.t16 45.5208
R88 source.n2 source.n1 44.201
R89 source.n4 source.n3 44.201
R90 source.n6 source.n5 44.201
R91 source.n10 source.n9 44.201
R92 source.n12 source.n11 44.201
R93 source.n14 source.n13 44.201
R94 source.n30 source.n29 44.2008
R95 source.n28 source.n27 44.2008
R96 source.n26 source.n25 44.2008
R97 source.n22 source.n21 44.2008
R98 source.n20 source.n19 44.2008
R99 source.n18 source.n17 44.2008
R100 source.n16 source.n15 24.5346
R101 source.n32 source.n0 18.7846
R102 source.n32 source.n31 5.7505
R103 source.n29 source.t1 1.3205
R104 source.n29 source.t7 1.3205
R105 source.n27 source.t10 1.3205
R106 source.n27 source.t5 1.3205
R107 source.n25 source.t4 1.3205
R108 source.n25 source.t30 1.3205
R109 source.n21 source.t23 1.3205
R110 source.n21 source.t21 1.3205
R111 source.n19 source.t14 1.3205
R112 source.n19 source.t29 1.3205
R113 source.n17 source.t15 1.3205
R114 source.n17 source.t25 1.3205
R115 source.n1 source.t17 1.3205
R116 source.n1 source.t19 1.3205
R117 source.n3 source.t28 1.3205
R118 source.n3 source.t22 1.3205
R119 source.n5 source.t27 1.3205
R120 source.n5 source.t26 1.3205
R121 source.n9 source.t2 1.3205
R122 source.n9 source.t13 1.3205
R123 source.n11 source.t0 1.3205
R124 source.n11 source.t31 1.3205
R125 source.n13 source.t6 1.3205
R126 source.n13 source.t11 1.3205
R127 source.n15 source.n14 0.974638
R128 source.n14 source.n12 0.974638
R129 source.n12 source.n10 0.974638
R130 source.n10 source.n8 0.974638
R131 source.n7 source.n6 0.974638
R132 source.n6 source.n4 0.974638
R133 source.n4 source.n2 0.974638
R134 source.n2 source.n0 0.974638
R135 source.n18 source.n16 0.974638
R136 source.n20 source.n18 0.974638
R137 source.n22 source.n20 0.974638
R138 source.n23 source.n22 0.974638
R139 source.n26 source.n24 0.974638
R140 source.n28 source.n26 0.974638
R141 source.n30 source.n28 0.974638
R142 source.n31 source.n30 0.974638
R143 source.n8 source.n7 0.470328
R144 source.n24 source.n23 0.470328
R145 source source.n32 0.188
R146 drain_left.n9 drain_left.n7 61.8539
R147 drain_left.n5 drain_left.n3 61.8537
R148 drain_left.n2 drain_left.n0 61.8537
R149 drain_left.n11 drain_left.n10 60.8798
R150 drain_left.n9 drain_left.n8 60.8798
R151 drain_left.n13 drain_left.n12 60.8796
R152 drain_left.n5 drain_left.n4 60.8796
R153 drain_left.n2 drain_left.n1 60.8796
R154 drain_left drain_left.n6 35.9717
R155 drain_left drain_left.n13 6.62735
R156 drain_left.n3 drain_left.t11 1.3205
R157 drain_left.n3 drain_left.t15 1.3205
R158 drain_left.n4 drain_left.t12 1.3205
R159 drain_left.n4 drain_left.t1 1.3205
R160 drain_left.n1 drain_left.t14 1.3205
R161 drain_left.n1 drain_left.t4 1.3205
R162 drain_left.n0 drain_left.t13 1.3205
R163 drain_left.n0 drain_left.t10 1.3205
R164 drain_left.n12 drain_left.t8 1.3205
R165 drain_left.n12 drain_left.t9 1.3205
R166 drain_left.n10 drain_left.t3 1.3205
R167 drain_left.n10 drain_left.t7 1.3205
R168 drain_left.n8 drain_left.t5 1.3205
R169 drain_left.n8 drain_left.t6 1.3205
R170 drain_left.n7 drain_left.t0 1.3205
R171 drain_left.n7 drain_left.t2 1.3205
R172 drain_left.n11 drain_left.n9 0.974638
R173 drain_left.n13 drain_left.n11 0.974638
R174 drain_left.n6 drain_left.n5 0.432223
R175 drain_left.n6 drain_left.n2 0.432223
R176 minus.n5 minus.t8 522.003
R177 minus.n27 minus.t1 522.003
R178 minus.n6 minus.t6 500.979
R179 minus.n7 minus.t4 500.979
R180 minus.n3 minus.t11 500.979
R181 minus.n13 minus.t12 500.979
R182 minus.n1 minus.t9 500.979
R183 minus.n18 minus.t7 500.979
R184 minus.n20 minus.t13 500.979
R185 minus.n28 minus.t10 500.979
R186 minus.n29 minus.t15 500.979
R187 minus.n25 minus.t5 500.979
R188 minus.n35 minus.t0 500.979
R189 minus.n23 minus.t3 500.979
R190 minus.n40 minus.t14 500.979
R191 minus.n42 minus.t2 500.979
R192 minus.n21 minus.n20 161.3
R193 minus.n19 minus.n0 161.3
R194 minus.n15 minus.n14 161.3
R195 minus.n13 minus.n2 161.3
R196 minus.n12 minus.n11 161.3
R197 minus.n10 minus.n3 161.3
R198 minus.n9 minus.n8 161.3
R199 minus.n43 minus.n42 161.3
R200 minus.n41 minus.n22 161.3
R201 minus.n37 minus.n36 161.3
R202 minus.n35 minus.n24 161.3
R203 minus.n34 minus.n33 161.3
R204 minus.n32 minus.n25 161.3
R205 minus.n31 minus.n30 161.3
R206 minus.n18 minus.n17 80.6037
R207 minus.n16 minus.n1 80.6037
R208 minus.n7 minus.n4 80.6037
R209 minus.n40 minus.n39 80.6037
R210 minus.n38 minus.n23 80.6037
R211 minus.n29 minus.n26 80.6037
R212 minus.n7 minus.n6 48.2005
R213 minus.n18 minus.n1 48.2005
R214 minus.n29 minus.n28 48.2005
R215 minus.n40 minus.n23 48.2005
R216 minus.n8 minus.n7 43.0884
R217 minus.n14 minus.n1 43.0884
R218 minus.n30 minus.n29 43.0884
R219 minus.n36 minus.n23 43.0884
R220 minus.n44 minus.n21 41.9664
R221 minus.n19 minus.n18 40.1672
R222 minus.n41 minus.n40 40.1672
R223 minus.n5 minus.n4 31.6481
R224 minus.n27 minus.n26 31.6481
R225 minus.n13 minus.n12 24.1005
R226 minus.n12 minus.n3 24.1005
R227 minus.n34 minus.n25 24.1005
R228 minus.n35 minus.n34 24.1005
R229 minus.n6 minus.n5 17.444
R230 minus.n28 minus.n27 17.444
R231 minus.n20 minus.n19 8.03383
R232 minus.n42 minus.n41 8.03383
R233 minus.n44 minus.n43 6.6558
R234 minus.n8 minus.n3 5.11262
R235 minus.n14 minus.n13 5.11262
R236 minus.n30 minus.n25 5.11262
R237 minus.n36 minus.n35 5.11262
R238 minus.n17 minus.n16 0.380177
R239 minus.n39 minus.n38 0.380177
R240 minus.n17 minus.n0 0.285035
R241 minus.n16 minus.n15 0.285035
R242 minus.n9 minus.n4 0.285035
R243 minus.n31 minus.n26 0.285035
R244 minus.n38 minus.n37 0.285035
R245 minus.n39 minus.n22 0.285035
R246 minus.n21 minus.n0 0.189894
R247 minus.n15 minus.n2 0.189894
R248 minus.n11 minus.n2 0.189894
R249 minus.n11 minus.n10 0.189894
R250 minus.n10 minus.n9 0.189894
R251 minus.n32 minus.n31 0.189894
R252 minus.n33 minus.n32 0.189894
R253 minus.n33 minus.n24 0.189894
R254 minus.n37 minus.n24 0.189894
R255 minus.n43 minus.n22 0.189894
R256 minus minus.n44 0.188
R257 drain_right.n9 drain_right.n7 61.8538
R258 drain_right.n5 drain_right.n3 61.8537
R259 drain_right.n2 drain_right.n0 61.8537
R260 drain_right.n9 drain_right.n8 60.8798
R261 drain_right.n11 drain_right.n10 60.8798
R262 drain_right.n13 drain_right.n12 60.8798
R263 drain_right.n5 drain_right.n4 60.8796
R264 drain_right.n2 drain_right.n1 60.8796
R265 drain_right drain_right.n6 35.4185
R266 drain_right drain_right.n13 6.62735
R267 drain_right.n3 drain_right.t1 1.3205
R268 drain_right.n3 drain_right.t13 1.3205
R269 drain_right.n4 drain_right.t15 1.3205
R270 drain_right.n4 drain_right.t12 1.3205
R271 drain_right.n1 drain_right.t0 1.3205
R272 drain_right.n1 drain_right.t10 1.3205
R273 drain_right.n0 drain_right.t14 1.3205
R274 drain_right.n0 drain_right.t5 1.3205
R275 drain_right.n7 drain_right.t9 1.3205
R276 drain_right.n7 drain_right.t7 1.3205
R277 drain_right.n8 drain_right.t4 1.3205
R278 drain_right.n8 drain_right.t11 1.3205
R279 drain_right.n10 drain_right.t6 1.3205
R280 drain_right.n10 drain_right.t3 1.3205
R281 drain_right.n12 drain_right.t2 1.3205
R282 drain_right.n12 drain_right.t8 1.3205
R283 drain_right.n13 drain_right.n11 0.974638
R284 drain_right.n11 drain_right.n9 0.974638
R285 drain_right.n6 drain_right.n5 0.432223
R286 drain_right.n6 drain_right.n2 0.432223
C0 drain_right plus 0.430381f
C1 minus plus 7.13158f
C2 drain_right minus 13.585401f
C3 plus drain_left 13.8587f
C4 plus source 13.5866f
C5 drain_right drain_left 1.44945f
C6 drain_right source 22.259901f
C7 minus drain_left 0.173489f
C8 minus source 13.5725f
C9 source drain_left 22.257101f
C10 drain_right a_n2750_n3888# 7.48085f
C11 drain_left a_n2750_n3888# 7.86813f
C12 source a_n2750_n3888# 11.084404f
C13 minus a_n2750_n3888# 11.217442f
C14 plus a_n2750_n3888# 13.057211f
C15 drain_right.t14 a_n2750_n3888# 0.314675f
C16 drain_right.t5 a_n2750_n3888# 0.314675f
C17 drain_right.n0 a_n2750_n3888# 2.85051f
C18 drain_right.t0 a_n2750_n3888# 0.314675f
C19 drain_right.t10 a_n2750_n3888# 0.314675f
C20 drain_right.n1 a_n2750_n3888# 2.8443f
C21 drain_right.n2 a_n2750_n3888# 0.727691f
C22 drain_right.t1 a_n2750_n3888# 0.314675f
C23 drain_right.t13 a_n2750_n3888# 0.314675f
C24 drain_right.n3 a_n2750_n3888# 2.85051f
C25 drain_right.t15 a_n2750_n3888# 0.314675f
C26 drain_right.t12 a_n2750_n3888# 0.314675f
C27 drain_right.n4 a_n2750_n3888# 2.8443f
C28 drain_right.n5 a_n2750_n3888# 0.727691f
C29 drain_right.n6 a_n2750_n3888# 1.71521f
C30 drain_right.t9 a_n2750_n3888# 0.314675f
C31 drain_right.t7 a_n2750_n3888# 0.314675f
C32 drain_right.n7 a_n2750_n3888# 2.85051f
C33 drain_right.t4 a_n2750_n3888# 0.314675f
C34 drain_right.t11 a_n2750_n3888# 0.314675f
C35 drain_right.n8 a_n2750_n3888# 2.8443f
C36 drain_right.n9 a_n2750_n3888# 0.772669f
C37 drain_right.t6 a_n2750_n3888# 0.314675f
C38 drain_right.t3 a_n2750_n3888# 0.314675f
C39 drain_right.n10 a_n2750_n3888# 2.8443f
C40 drain_right.n11 a_n2750_n3888# 0.384092f
C41 drain_right.t2 a_n2750_n3888# 0.314675f
C42 drain_right.t8 a_n2750_n3888# 0.314675f
C43 drain_right.n12 a_n2750_n3888# 2.8443f
C44 drain_right.n13 a_n2750_n3888# 0.622139f
C45 minus.n0 a_n2750_n3888# 0.051089f
C46 minus.t9 a_n2750_n3888# 1.3056f
C47 minus.n1 a_n2750_n3888# 0.511267f
C48 minus.t7 a_n2750_n3888# 1.3056f
C49 minus.n2 a_n2750_n3888# 0.038287f
C50 minus.t11 a_n2750_n3888# 1.3056f
C51 minus.n3 a_n2750_n3888# 0.500336f
C52 minus.n4 a_n2750_n3888# 0.219595f
C53 minus.t8 a_n2750_n3888# 1.32589f
C54 minus.n5 a_n2750_n3888# 0.486826f
C55 minus.t6 a_n2750_n3888# 1.3056f
C56 minus.n6 a_n2750_n3888# 0.511566f
C57 minus.t4 a_n2750_n3888# 1.3056f
C58 minus.n7 a_n2750_n3888# 0.511267f
C59 minus.n8 a_n2750_n3888# 0.008688f
C60 minus.n9 a_n2750_n3888# 0.051089f
C61 minus.n10 a_n2750_n3888# 0.038287f
C62 minus.n11 a_n2750_n3888# 0.038287f
C63 minus.n12 a_n2750_n3888# 0.008688f
C64 minus.t12 a_n2750_n3888# 1.3056f
C65 minus.n13 a_n2750_n3888# 0.500336f
C66 minus.n14 a_n2750_n3888# 0.008688f
C67 minus.n15 a_n2750_n3888# 0.051089f
C68 minus.n16 a_n2750_n3888# 0.063772f
C69 minus.n17 a_n2750_n3888# 0.063772f
C70 minus.n18 a_n2750_n3888# 0.510794f
C71 minus.n19 a_n2750_n3888# 0.008688f
C72 minus.t13 a_n2750_n3888# 1.3056f
C73 minus.n20 a_n2750_n3888# 0.496913f
C74 minus.n21 a_n2750_n3888# 1.69757f
C75 minus.n22 a_n2750_n3888# 0.051089f
C76 minus.t3 a_n2750_n3888# 1.3056f
C77 minus.n23 a_n2750_n3888# 0.511267f
C78 minus.n24 a_n2750_n3888# 0.038287f
C79 minus.t5 a_n2750_n3888# 1.3056f
C80 minus.n25 a_n2750_n3888# 0.500336f
C81 minus.n26 a_n2750_n3888# 0.219595f
C82 minus.t1 a_n2750_n3888# 1.32589f
C83 minus.n27 a_n2750_n3888# 0.486826f
C84 minus.t10 a_n2750_n3888# 1.3056f
C85 minus.n28 a_n2750_n3888# 0.511566f
C86 minus.t15 a_n2750_n3888# 1.3056f
C87 minus.n29 a_n2750_n3888# 0.511267f
C88 minus.n30 a_n2750_n3888# 0.008688f
C89 minus.n31 a_n2750_n3888# 0.051089f
C90 minus.n32 a_n2750_n3888# 0.038287f
C91 minus.n33 a_n2750_n3888# 0.038287f
C92 minus.n34 a_n2750_n3888# 0.008688f
C93 minus.t0 a_n2750_n3888# 1.3056f
C94 minus.n35 a_n2750_n3888# 0.500336f
C95 minus.n36 a_n2750_n3888# 0.008688f
C96 minus.n37 a_n2750_n3888# 0.051089f
C97 minus.n38 a_n2750_n3888# 0.063772f
C98 minus.n39 a_n2750_n3888# 0.063772f
C99 minus.t14 a_n2750_n3888# 1.3056f
C100 minus.n40 a_n2750_n3888# 0.510794f
C101 minus.n41 a_n2750_n3888# 0.008688f
C102 minus.t2 a_n2750_n3888# 1.3056f
C103 minus.n42 a_n2750_n3888# 0.496913f
C104 minus.n43 a_n2750_n3888# 0.264263f
C105 minus.n44 a_n2750_n3888# 2.02413f
C106 drain_left.t13 a_n2750_n3888# 0.31639f
C107 drain_left.t10 a_n2750_n3888# 0.31639f
C108 drain_left.n0 a_n2750_n3888# 2.86604f
C109 drain_left.t14 a_n2750_n3888# 0.31639f
C110 drain_left.t4 a_n2750_n3888# 0.31639f
C111 drain_left.n1 a_n2750_n3888# 2.85979f
C112 drain_left.n2 a_n2750_n3888# 0.731655f
C113 drain_left.t11 a_n2750_n3888# 0.31639f
C114 drain_left.t15 a_n2750_n3888# 0.31639f
C115 drain_left.n3 a_n2750_n3888# 2.86604f
C116 drain_left.t12 a_n2750_n3888# 0.31639f
C117 drain_left.t1 a_n2750_n3888# 0.31639f
C118 drain_left.n4 a_n2750_n3888# 2.85979f
C119 drain_left.n5 a_n2750_n3888# 0.731655f
C120 drain_left.n6 a_n2750_n3888# 1.77933f
C121 drain_left.t0 a_n2750_n3888# 0.31639f
C122 drain_left.t2 a_n2750_n3888# 0.31639f
C123 drain_left.n7 a_n2750_n3888# 2.86605f
C124 drain_left.t5 a_n2750_n3888# 0.31639f
C125 drain_left.t6 a_n2750_n3888# 0.31639f
C126 drain_left.n8 a_n2750_n3888# 2.8598f
C127 drain_left.n9 a_n2750_n3888# 0.776869f
C128 drain_left.t3 a_n2750_n3888# 0.31639f
C129 drain_left.t7 a_n2750_n3888# 0.31639f
C130 drain_left.n10 a_n2750_n3888# 2.8598f
C131 drain_left.n11 a_n2750_n3888# 0.386185f
C132 drain_left.t8 a_n2750_n3888# 0.31639f
C133 drain_left.t9 a_n2750_n3888# 0.31639f
C134 drain_left.n12 a_n2750_n3888# 2.85979f
C135 drain_left.n13 a_n2750_n3888# 0.625538f
C136 source.t16 a_n2750_n3888# 2.99103f
C137 source.n0 a_n2750_n3888# 1.43579f
C138 source.t17 a_n2750_n3888# 0.266899f
C139 source.t19 a_n2750_n3888# 0.266899f
C140 source.n1 a_n2750_n3888# 2.34448f
C141 source.n2 a_n2750_n3888# 0.363144f
C142 source.t28 a_n2750_n3888# 0.266899f
C143 source.t22 a_n2750_n3888# 0.266899f
C144 source.n3 a_n2750_n3888# 2.34448f
C145 source.n4 a_n2750_n3888# 0.363144f
C146 source.t27 a_n2750_n3888# 0.266899f
C147 source.t26 a_n2750_n3888# 0.266899f
C148 source.n5 a_n2750_n3888# 2.34448f
C149 source.n6 a_n2750_n3888# 0.363144f
C150 source.t20 a_n2750_n3888# 2.99103f
C151 source.n7 a_n2750_n3888# 0.407908f
C152 source.t12 a_n2750_n3888# 2.99103f
C153 source.n8 a_n2750_n3888# 0.407908f
C154 source.t2 a_n2750_n3888# 0.266899f
C155 source.t13 a_n2750_n3888# 0.266899f
C156 source.n9 a_n2750_n3888# 2.34448f
C157 source.n10 a_n2750_n3888# 0.363144f
C158 source.t0 a_n2750_n3888# 0.266899f
C159 source.t31 a_n2750_n3888# 0.266899f
C160 source.n11 a_n2750_n3888# 2.34448f
C161 source.n12 a_n2750_n3888# 0.363144f
C162 source.t6 a_n2750_n3888# 0.266899f
C163 source.t11 a_n2750_n3888# 0.266899f
C164 source.n13 a_n2750_n3888# 2.34448f
C165 source.n14 a_n2750_n3888# 0.363144f
C166 source.t3 a_n2750_n3888# 2.99103f
C167 source.n15 a_n2750_n3888# 1.82229f
C168 source.t18 a_n2750_n3888# 2.99103f
C169 source.n16 a_n2750_n3888# 1.82229f
C170 source.t15 a_n2750_n3888# 0.266899f
C171 source.t25 a_n2750_n3888# 0.266899f
C172 source.n17 a_n2750_n3888# 2.34448f
C173 source.n18 a_n2750_n3888# 0.363147f
C174 source.t14 a_n2750_n3888# 0.266899f
C175 source.t29 a_n2750_n3888# 0.266899f
C176 source.n19 a_n2750_n3888# 2.34448f
C177 source.n20 a_n2750_n3888# 0.363147f
C178 source.t23 a_n2750_n3888# 0.266899f
C179 source.t21 a_n2750_n3888# 0.266899f
C180 source.n21 a_n2750_n3888# 2.34448f
C181 source.n22 a_n2750_n3888# 0.363147f
C182 source.t24 a_n2750_n3888# 2.99103f
C183 source.n23 a_n2750_n3888# 0.407912f
C184 source.t8 a_n2750_n3888# 2.99103f
C185 source.n24 a_n2750_n3888# 0.407912f
C186 source.t4 a_n2750_n3888# 0.266899f
C187 source.t30 a_n2750_n3888# 0.266899f
C188 source.n25 a_n2750_n3888# 2.34448f
C189 source.n26 a_n2750_n3888# 0.363147f
C190 source.t10 a_n2750_n3888# 0.266899f
C191 source.t5 a_n2750_n3888# 0.266899f
C192 source.n27 a_n2750_n3888# 2.34448f
C193 source.n28 a_n2750_n3888# 0.363147f
C194 source.t1 a_n2750_n3888# 0.266899f
C195 source.t7 a_n2750_n3888# 0.266899f
C196 source.n29 a_n2750_n3888# 2.34448f
C197 source.n30 a_n2750_n3888# 0.363147f
C198 source.t9 a_n2750_n3888# 2.99103f
C199 source.n31 a_n2750_n3888# 0.559662f
C200 source.n32 a_n2750_n3888# 1.66515f
C201 plus.n0 a_n2750_n3888# 0.051653f
C202 plus.t6 a_n2750_n3888# 1.32f
C203 plus.t7 a_n2750_n3888# 1.32f
C204 plus.n1 a_n2750_n3888# 0.064475f
C205 plus.t8 a_n2750_n3888# 1.32f
C206 plus.n2 a_n2750_n3888# 0.064475f
C207 plus.t12 a_n2750_n3888# 1.32f
C208 plus.n3 a_n2750_n3888# 0.505854f
C209 plus.n4 a_n2750_n3888# 0.038709f
C210 plus.t9 a_n2750_n3888# 1.32f
C211 plus.t10 a_n2750_n3888# 1.32f
C212 plus.n5 a_n2750_n3888# 0.516905f
C213 plus.t13 a_n2750_n3888# 1.32f
C214 plus.n6 a_n2750_n3888# 0.517208f
C215 plus.t15 a_n2750_n3888# 1.34051f
C216 plus.n7 a_n2750_n3888# 0.492195f
C217 plus.n8 a_n2750_n3888# 0.222017f
C218 plus.n9 a_n2750_n3888# 0.051653f
C219 plus.n10 a_n2750_n3888# 0.008784f
C220 plus.n11 a_n2750_n3888# 0.505854f
C221 plus.n12 a_n2750_n3888# 0.008784f
C222 plus.n13 a_n2750_n3888# 0.038709f
C223 plus.n14 a_n2750_n3888# 0.038709f
C224 plus.n15 a_n2750_n3888# 0.051653f
C225 plus.n16 a_n2750_n3888# 0.008784f
C226 plus.n17 a_n2750_n3888# 0.516905f
C227 plus.n18 a_n2750_n3888# 0.516428f
C228 plus.n19 a_n2750_n3888# 0.008784f
C229 plus.n20 a_n2750_n3888# 0.502393f
C230 plus.n21 a_n2750_n3888# 0.50332f
C231 plus.n22 a_n2750_n3888# 0.051653f
C232 plus.t2 a_n2750_n3888# 1.32f
C233 plus.n23 a_n2750_n3888# 0.064475f
C234 plus.t5 a_n2750_n3888# 1.32f
C235 plus.n24 a_n2750_n3888# 0.064475f
C236 plus.t1 a_n2750_n3888# 1.32f
C237 plus.t11 a_n2750_n3888# 1.32f
C238 plus.n25 a_n2750_n3888# 0.505854f
C239 plus.n26 a_n2750_n3888# 0.038709f
C240 plus.t3 a_n2750_n3888# 1.32f
C241 plus.t14 a_n2750_n3888# 1.32f
C242 plus.n27 a_n2750_n3888# 0.516905f
C243 plus.t4 a_n2750_n3888# 1.32f
C244 plus.n28 a_n2750_n3888# 0.517208f
C245 plus.t0 a_n2750_n3888# 1.34051f
C246 plus.n29 a_n2750_n3888# 0.492195f
C247 plus.n30 a_n2750_n3888# 0.222017f
C248 plus.n31 a_n2750_n3888# 0.051653f
C249 plus.n32 a_n2750_n3888# 0.008784f
C250 plus.n33 a_n2750_n3888# 0.505854f
C251 plus.n34 a_n2750_n3888# 0.008784f
C252 plus.n35 a_n2750_n3888# 0.038709f
C253 plus.n36 a_n2750_n3888# 0.038709f
C254 plus.n37 a_n2750_n3888# 0.051653f
C255 plus.n38 a_n2750_n3888# 0.008784f
C256 plus.n39 a_n2750_n3888# 0.516905f
C257 plus.n40 a_n2750_n3888# 0.516428f
C258 plus.n41 a_n2750_n3888# 0.008784f
C259 plus.n42 a_n2750_n3888# 0.502393f
C260 plus.n43 a_n2750_n3888# 1.42943f
.ends

