* NGSPICE file created from diffpair558.ext - technology: sky130A

.subckt diffpair558 minus drain_right drain_left source plus
X0 source.t38 plus.t0 drain_left.t4 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X1 a_n3202_n3888# a_n3202_n3888# a_n3202_n3888# a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.8
X2 drain_left.t3 plus.t1 source.t37 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X3 source.t18 minus.t0 drain_right.t19 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X4 a_n3202_n3888# a_n3202_n3888# a_n3202_n3888# a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X5 source.t5 minus.t1 drain_right.t18 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X6 source.t36 plus.t2 drain_left.t2 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X7 drain_right.t17 minus.t2 source.t9 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X8 drain_right.t16 minus.t3 source.t17 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X9 source.t35 plus.t3 drain_left.t17 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X10 drain_right.t15 minus.t4 source.t4 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X11 source.t8 minus.t5 drain_right.t14 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X12 drain_right.t13 minus.t6 source.t10 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X13 drain_right.t12 minus.t7 source.t12 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X14 source.t34 plus.t4 drain_left.t16 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X15 drain_left.t6 plus.t5 source.t33 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X16 source.t15 minus.t8 drain_right.t11 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X17 a_n3202_n3888# a_n3202_n3888# a_n3202_n3888# a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X18 drain_right.t10 minus.t9 source.t16 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X19 source.t32 plus.t6 drain_left.t5 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X20 drain_left.t12 plus.t7 source.t31 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X21 drain_right.t9 minus.t10 source.t39 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X22 source.t30 plus.t8 drain_left.t11 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X23 source.t3 minus.t11 drain_right.t8 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X24 drain_right.t7 minus.t12 source.t11 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X25 drain_left.t19 plus.t9 source.t29 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X26 drain_left.t18 plus.t10 source.t28 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X27 source.t13 minus.t13 drain_right.t6 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X28 drain_right.t5 minus.t14 source.t14 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X29 drain_right.t4 minus.t15 source.t0 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X30 a_n3202_n3888# a_n3202_n3888# a_n3202_n3888# a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X31 source.t27 plus.t11 drain_left.t14 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X32 drain_left.t13 plus.t12 source.t26 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X33 drain_left.t1 plus.t13 source.t25 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X34 source.t2 minus.t16 drain_right.t3 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X35 source.t24 plus.t14 drain_left.t0 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X36 drain_left.t8 plus.t15 source.t23 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X37 source.t22 plus.t16 drain_left.t7 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X38 drain_left.t10 plus.t17 source.t21 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X39 drain_left.t9 plus.t18 source.t20 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X40 source.t1 minus.t17 drain_right.t2 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X41 source.t19 plus.t19 drain_left.t15 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X42 source.t6 minus.t18 drain_right.t1 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X43 source.t7 minus.t19 drain_right.t0 a_n3202_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
R0 plus.n9 plus.t19 522.769
R1 plus.n39 plus.t1 522.769
R2 plus.n28 plus.t5 500.979
R3 plus.n26 plus.t8 500.979
R4 plus.n2 plus.t10 500.979
R5 plus.n21 plus.t11 500.979
R6 plus.n19 plus.t12 500.979
R7 plus.n5 plus.t16 500.979
R8 plus.n13 plus.t13 500.979
R9 plus.n12 plus.t14 500.979
R10 plus.n8 plus.t17 500.979
R11 plus.n58 plus.t0 500.979
R12 plus.n56 plus.t7 500.979
R13 plus.n32 plus.t3 500.979
R14 plus.n51 plus.t9 500.979
R15 plus.n49 plus.t2 500.979
R16 plus.n35 plus.t15 500.979
R17 plus.n43 plus.t4 500.979
R18 plus.n42 plus.t18 500.979
R19 plus.n38 plus.t6 500.979
R20 plus.n11 plus.n10 161.3
R21 plus.n15 plus.n14 161.3
R22 plus.n16 plus.n5 161.3
R23 plus.n18 plus.n17 161.3
R24 plus.n19 plus.n4 161.3
R25 plus.n20 plus.n3 161.3
R26 plus.n25 plus.n24 161.3
R27 plus.n26 plus.n1 161.3
R28 plus.n27 plus.n0 161.3
R29 plus.n29 plus.n28 161.3
R30 plus.n41 plus.n40 161.3
R31 plus.n45 plus.n44 161.3
R32 plus.n46 plus.n35 161.3
R33 plus.n48 plus.n47 161.3
R34 plus.n49 plus.n34 161.3
R35 plus.n50 plus.n33 161.3
R36 plus.n55 plus.n54 161.3
R37 plus.n56 plus.n31 161.3
R38 plus.n57 plus.n30 161.3
R39 plus.n59 plus.n58 161.3
R40 plus.n12 plus.n7 80.6037
R41 plus.n13 plus.n6 80.6037
R42 plus.n22 plus.n21 80.6037
R43 plus.n23 plus.n2 80.6037
R44 plus.n42 plus.n37 80.6037
R45 plus.n43 plus.n36 80.6037
R46 plus.n52 plus.n51 80.6037
R47 plus.n53 plus.n32 80.6037
R48 plus.n21 plus.n2 48.2005
R49 plus.n13 plus.n12 48.2005
R50 plus.n51 plus.n32 48.2005
R51 plus.n43 plus.n42 48.2005
R52 plus.n40 plus.n39 44.8565
R53 plus.n10 plus.n9 44.8565
R54 plus.n21 plus.n20 43.0884
R55 plus.n14 plus.n13 43.0884
R56 plus.n51 plus.n50 43.0884
R57 plus.n44 plus.n43 43.0884
R58 plus.n25 plus.n2 40.1672
R59 plus.n12 plus.n11 40.1672
R60 plus.n55 plus.n32 40.1672
R61 plus.n42 plus.n41 40.1672
R62 plus plus.n59 36.4725
R63 plus.n28 plus.n27 27.0217
R64 plus.n58 plus.n57 27.0217
R65 plus.n18 plus.n5 24.1005
R66 plus.n19 plus.n18 24.1005
R67 plus.n49 plus.n48 24.1005
R68 plus.n48 plus.n35 24.1005
R69 plus.n27 plus.n26 21.1793
R70 plus.n57 plus.n56 21.1793
R71 plus.n39 plus.n38 20.1275
R72 plus.n9 plus.n8 20.1275
R73 plus plus.n29 13.4853
R74 plus.n26 plus.n25 8.03383
R75 plus.n11 plus.n8 8.03383
R76 plus.n56 plus.n55 8.03383
R77 plus.n41 plus.n38 8.03383
R78 plus.n20 plus.n19 5.11262
R79 plus.n14 plus.n5 5.11262
R80 plus.n50 plus.n49 5.11262
R81 plus.n44 plus.n35 5.11262
R82 plus.n7 plus.n6 0.380177
R83 plus.n23 plus.n22 0.380177
R84 plus.n53 plus.n52 0.380177
R85 plus.n37 plus.n36 0.380177
R86 plus.n10 plus.n7 0.285035
R87 plus.n15 plus.n6 0.285035
R88 plus.n22 plus.n3 0.285035
R89 plus.n24 plus.n23 0.285035
R90 plus.n54 plus.n53 0.285035
R91 plus.n52 plus.n33 0.285035
R92 plus.n45 plus.n36 0.285035
R93 plus.n40 plus.n37 0.285035
R94 plus.n16 plus.n15 0.189894
R95 plus.n17 plus.n16 0.189894
R96 plus.n17 plus.n4 0.189894
R97 plus.n4 plus.n3 0.189894
R98 plus.n24 plus.n1 0.189894
R99 plus.n1 plus.n0 0.189894
R100 plus.n29 plus.n0 0.189894
R101 plus.n59 plus.n30 0.189894
R102 plus.n31 plus.n30 0.189894
R103 plus.n54 plus.n31 0.189894
R104 plus.n34 plus.n33 0.189894
R105 plus.n47 plus.n34 0.189894
R106 plus.n47 plus.n46 0.189894
R107 plus.n46 plus.n45 0.189894
R108 drain_left.n10 drain_left.n8 61.8539
R109 drain_left.n6 drain_left.n4 61.8537
R110 drain_left.n2 drain_left.n0 61.8537
R111 drain_left.n14 drain_left.n13 60.8798
R112 drain_left.n12 drain_left.n11 60.8798
R113 drain_left.n10 drain_left.n9 60.8798
R114 drain_left.n16 drain_left.n15 60.8796
R115 drain_left.n7 drain_left.n3 60.8796
R116 drain_left.n6 drain_left.n5 60.8796
R117 drain_left.n2 drain_left.n1 60.8796
R118 drain_left drain_left.n7 37.4329
R119 drain_left drain_left.n16 6.62735
R120 drain_left.n3 drain_left.t2 1.3205
R121 drain_left.n3 drain_left.t8 1.3205
R122 drain_left.n4 drain_left.t5 1.3205
R123 drain_left.n4 drain_left.t3 1.3205
R124 drain_left.n5 drain_left.t16 1.3205
R125 drain_left.n5 drain_left.t9 1.3205
R126 drain_left.n1 drain_left.t17 1.3205
R127 drain_left.n1 drain_left.t19 1.3205
R128 drain_left.n0 drain_left.t4 1.3205
R129 drain_left.n0 drain_left.t12 1.3205
R130 drain_left.n15 drain_left.t11 1.3205
R131 drain_left.n15 drain_left.t6 1.3205
R132 drain_left.n13 drain_left.t14 1.3205
R133 drain_left.n13 drain_left.t18 1.3205
R134 drain_left.n11 drain_left.t7 1.3205
R135 drain_left.n11 drain_left.t13 1.3205
R136 drain_left.n9 drain_left.t0 1.3205
R137 drain_left.n9 drain_left.t1 1.3205
R138 drain_left.n8 drain_left.t15 1.3205
R139 drain_left.n8 drain_left.t10 1.3205
R140 drain_left.n12 drain_left.n10 0.974638
R141 drain_left.n14 drain_left.n12 0.974638
R142 drain_left.n16 drain_left.n14 0.974638
R143 drain_left.n7 drain_left.n6 0.919292
R144 drain_left.n7 drain_left.n2 0.919292
R145 source.n9 source.t19 45.521
R146 source.n10 source.t39 45.521
R147 source.n19 source.t8 45.521
R148 source.n39 source.t17 45.5208
R149 source.n30 source.t5 45.5208
R150 source.n29 source.t37 45.5208
R151 source.n20 source.t38 45.5208
R152 source.n0 source.t33 45.5208
R153 source.n2 source.n1 44.201
R154 source.n4 source.n3 44.201
R155 source.n6 source.n5 44.201
R156 source.n8 source.n7 44.201
R157 source.n12 source.n11 44.201
R158 source.n14 source.n13 44.201
R159 source.n16 source.n15 44.201
R160 source.n18 source.n17 44.201
R161 source.n38 source.n37 44.2008
R162 source.n36 source.n35 44.2008
R163 source.n34 source.n33 44.2008
R164 source.n32 source.n31 44.2008
R165 source.n28 source.n27 44.2008
R166 source.n26 source.n25 44.2008
R167 source.n24 source.n23 44.2008
R168 source.n22 source.n21 44.2008
R169 source.n20 source.n19 24.5346
R170 source.n40 source.n0 18.7846
R171 source.n40 source.n39 5.7505
R172 source.n37 source.t9 1.3205
R173 source.n37 source.t7 1.3205
R174 source.n35 source.t4 1.3205
R175 source.n35 source.t1 1.3205
R176 source.n33 source.t12 1.3205
R177 source.n33 source.t18 1.3205
R178 source.n31 source.t11 1.3205
R179 source.n31 source.t6 1.3205
R180 source.n27 source.t20 1.3205
R181 source.n27 source.t32 1.3205
R182 source.n25 source.t23 1.3205
R183 source.n25 source.t34 1.3205
R184 source.n23 source.t29 1.3205
R185 source.n23 source.t36 1.3205
R186 source.n21 source.t31 1.3205
R187 source.n21 source.t35 1.3205
R188 source.n1 source.t28 1.3205
R189 source.n1 source.t30 1.3205
R190 source.n3 source.t26 1.3205
R191 source.n3 source.t27 1.3205
R192 source.n5 source.t25 1.3205
R193 source.n5 source.t22 1.3205
R194 source.n7 source.t21 1.3205
R195 source.n7 source.t24 1.3205
R196 source.n11 source.t10 1.3205
R197 source.n11 source.t15 1.3205
R198 source.n13 source.t0 1.3205
R199 source.n13 source.t13 1.3205
R200 source.n15 source.t16 1.3205
R201 source.n15 source.t3 1.3205
R202 source.n17 source.t14 1.3205
R203 source.n17 source.t2 1.3205
R204 source.n19 source.n18 0.974638
R205 source.n18 source.n16 0.974638
R206 source.n16 source.n14 0.974638
R207 source.n14 source.n12 0.974638
R208 source.n12 source.n10 0.974638
R209 source.n9 source.n8 0.974638
R210 source.n8 source.n6 0.974638
R211 source.n6 source.n4 0.974638
R212 source.n4 source.n2 0.974638
R213 source.n2 source.n0 0.974638
R214 source.n22 source.n20 0.974638
R215 source.n24 source.n22 0.974638
R216 source.n26 source.n24 0.974638
R217 source.n28 source.n26 0.974638
R218 source.n29 source.n28 0.974638
R219 source.n32 source.n30 0.974638
R220 source.n34 source.n32 0.974638
R221 source.n36 source.n34 0.974638
R222 source.n38 source.n36 0.974638
R223 source.n39 source.n38 0.974638
R224 source.n10 source.n9 0.470328
R225 source.n30 source.n29 0.470328
R226 source source.n40 0.188
R227 minus.n7 minus.t10 522.769
R228 minus.n37 minus.t1 522.769
R229 minus.n8 minus.t8 500.979
R230 minus.n10 minus.t6 500.979
R231 minus.n5 minus.t13 500.979
R232 minus.n15 minus.t15 500.979
R233 minus.n3 minus.t11 500.979
R234 minus.n21 minus.t9 500.979
R235 minus.n22 minus.t16 500.979
R236 minus.n26 minus.t14 500.979
R237 minus.n28 minus.t5 500.979
R238 minus.n38 minus.t12 500.979
R239 minus.n40 minus.t18 500.979
R240 minus.n35 minus.t7 500.979
R241 minus.n45 minus.t0 500.979
R242 minus.n33 minus.t4 500.979
R243 minus.n51 minus.t17 500.979
R244 minus.n52 minus.t2 500.979
R245 minus.n56 minus.t19 500.979
R246 minus.n58 minus.t3 500.979
R247 minus.n29 minus.n28 161.3
R248 minus.n27 minus.n0 161.3
R249 minus.n26 minus.n25 161.3
R250 minus.n24 minus.n1 161.3
R251 minus.n20 minus.n19 161.3
R252 minus.n18 minus.n3 161.3
R253 minus.n17 minus.n16 161.3
R254 minus.n15 minus.n4 161.3
R255 minus.n14 minus.n13 161.3
R256 minus.n9 minus.n6 161.3
R257 minus.n59 minus.n58 161.3
R258 minus.n57 minus.n30 161.3
R259 minus.n56 minus.n55 161.3
R260 minus.n54 minus.n31 161.3
R261 minus.n50 minus.n49 161.3
R262 minus.n48 minus.n33 161.3
R263 minus.n47 minus.n46 161.3
R264 minus.n45 minus.n34 161.3
R265 minus.n44 minus.n43 161.3
R266 minus.n39 minus.n36 161.3
R267 minus.n23 minus.n22 80.6037
R268 minus.n21 minus.n2 80.6037
R269 minus.n12 minus.n5 80.6037
R270 minus.n11 minus.n10 80.6037
R271 minus.n53 minus.n52 80.6037
R272 minus.n51 minus.n32 80.6037
R273 minus.n42 minus.n35 80.6037
R274 minus.n41 minus.n40 80.6037
R275 minus.n10 minus.n5 48.2005
R276 minus.n22 minus.n21 48.2005
R277 minus.n40 minus.n35 48.2005
R278 minus.n52 minus.n51 48.2005
R279 minus.n7 minus.n6 44.8565
R280 minus.n37 minus.n36 44.8565
R281 minus.n60 minus.n29 43.7278
R282 minus.n14 minus.n5 43.0884
R283 minus.n21 minus.n20 43.0884
R284 minus.n44 minus.n35 43.0884
R285 minus.n51 minus.n50 43.0884
R286 minus.n10 minus.n9 40.1672
R287 minus.n22 minus.n1 40.1672
R288 minus.n40 minus.n39 40.1672
R289 minus.n52 minus.n31 40.1672
R290 minus.n28 minus.n27 27.0217
R291 minus.n58 minus.n57 27.0217
R292 minus.n16 minus.n3 24.1005
R293 minus.n16 minus.n15 24.1005
R294 minus.n46 minus.n45 24.1005
R295 minus.n46 minus.n33 24.1005
R296 minus.n27 minus.n26 21.1793
R297 minus.n57 minus.n56 21.1793
R298 minus.n8 minus.n7 20.1275
R299 minus.n38 minus.n37 20.1275
R300 minus.n9 minus.n8 8.03383
R301 minus.n26 minus.n1 8.03383
R302 minus.n39 minus.n38 8.03383
R303 minus.n56 minus.n31 8.03383
R304 minus.n60 minus.n59 6.70505
R305 minus.n15 minus.n14 5.11262
R306 minus.n20 minus.n3 5.11262
R307 minus.n45 minus.n44 5.11262
R308 minus.n50 minus.n33 5.11262
R309 minus.n23 minus.n2 0.380177
R310 minus.n12 minus.n11 0.380177
R311 minus.n42 minus.n41 0.380177
R312 minus.n53 minus.n32 0.380177
R313 minus.n24 minus.n23 0.285035
R314 minus.n19 minus.n2 0.285035
R315 minus.n13 minus.n12 0.285035
R316 minus.n11 minus.n6 0.285035
R317 minus.n41 minus.n36 0.285035
R318 minus.n43 minus.n42 0.285035
R319 minus.n49 minus.n32 0.285035
R320 minus.n54 minus.n53 0.285035
R321 minus.n29 minus.n0 0.189894
R322 minus.n25 minus.n0 0.189894
R323 minus.n25 minus.n24 0.189894
R324 minus.n19 minus.n18 0.189894
R325 minus.n18 minus.n17 0.189894
R326 minus.n17 minus.n4 0.189894
R327 minus.n13 minus.n4 0.189894
R328 minus.n43 minus.n34 0.189894
R329 minus.n47 minus.n34 0.189894
R330 minus.n48 minus.n47 0.189894
R331 minus.n49 minus.n48 0.189894
R332 minus.n55 minus.n54 0.189894
R333 minus.n55 minus.n30 0.189894
R334 minus.n59 minus.n30 0.189894
R335 minus minus.n60 0.188
R336 drain_right.n10 drain_right.n8 61.8538
R337 drain_right.n6 drain_right.n4 61.8537
R338 drain_right.n2 drain_right.n0 61.8537
R339 drain_right.n10 drain_right.n9 60.8798
R340 drain_right.n12 drain_right.n11 60.8798
R341 drain_right.n14 drain_right.n13 60.8798
R342 drain_right.n16 drain_right.n15 60.8798
R343 drain_right.n7 drain_right.n3 60.8796
R344 drain_right.n6 drain_right.n5 60.8796
R345 drain_right.n2 drain_right.n1 60.8796
R346 drain_right drain_right.n7 36.8797
R347 drain_right drain_right.n16 6.62735
R348 drain_right.n3 drain_right.t19 1.3205
R349 drain_right.n3 drain_right.t15 1.3205
R350 drain_right.n4 drain_right.t0 1.3205
R351 drain_right.n4 drain_right.t16 1.3205
R352 drain_right.n5 drain_right.t2 1.3205
R353 drain_right.n5 drain_right.t17 1.3205
R354 drain_right.n1 drain_right.t1 1.3205
R355 drain_right.n1 drain_right.t12 1.3205
R356 drain_right.n0 drain_right.t18 1.3205
R357 drain_right.n0 drain_right.t7 1.3205
R358 drain_right.n8 drain_right.t11 1.3205
R359 drain_right.n8 drain_right.t9 1.3205
R360 drain_right.n9 drain_right.t6 1.3205
R361 drain_right.n9 drain_right.t13 1.3205
R362 drain_right.n11 drain_right.t8 1.3205
R363 drain_right.n11 drain_right.t4 1.3205
R364 drain_right.n13 drain_right.t3 1.3205
R365 drain_right.n13 drain_right.t10 1.3205
R366 drain_right.n15 drain_right.t14 1.3205
R367 drain_right.n15 drain_right.t5 1.3205
R368 drain_right.n16 drain_right.n14 0.974638
R369 drain_right.n14 drain_right.n12 0.974638
R370 drain_right.n12 drain_right.n10 0.974638
R371 drain_right.n7 drain_right.n6 0.919292
R372 drain_right.n7 drain_right.n2 0.919292
C0 plus drain_left 17.0667f
C1 source plus 16.8861f
C2 minus plus 7.69386f
C3 drain_right drain_left 1.72917f
C4 drain_right source 27.0357f
C5 drain_right minus 16.7463f
C6 source drain_left 27.0328f
C7 minus drain_left 0.17405f
C8 source minus 16.8721f
C9 drain_right plus 0.478206f
C10 drain_right a_n3202_n3888# 8.047379f
C11 drain_left a_n3202_n3888# 8.495999f
C12 source a_n3202_n3888# 11.254059f
C13 minus a_n3202_n3888# 13.137457f
C14 plus a_n3202_n3888# 15.047881f
C15 drain_right.t18 a_n3202_n3888# 0.313488f
C16 drain_right.t7 a_n3202_n3888# 0.313488f
C17 drain_right.n0 a_n3202_n3888# 2.83976f
C18 drain_right.t1 a_n3202_n3888# 0.313488f
C19 drain_right.t12 a_n3202_n3888# 0.313488f
C20 drain_right.n1 a_n3202_n3888# 2.83357f
C21 drain_right.n2 a_n3202_n3888# 0.7657f
C22 drain_right.t19 a_n3202_n3888# 0.313488f
C23 drain_right.t15 a_n3202_n3888# 0.313488f
C24 drain_right.n3 a_n3202_n3888# 2.83357f
C25 drain_right.t0 a_n3202_n3888# 0.313488f
C26 drain_right.t16 a_n3202_n3888# 0.313488f
C27 drain_right.n4 a_n3202_n3888# 2.83976f
C28 drain_right.t2 a_n3202_n3888# 0.313488f
C29 drain_right.t17 a_n3202_n3888# 0.313488f
C30 drain_right.n5 a_n3202_n3888# 2.83357f
C31 drain_right.n6 a_n3202_n3888# 0.7657f
C32 drain_right.n7 a_n3202_n3888# 2.13468f
C33 drain_right.t11 a_n3202_n3888# 0.313488f
C34 drain_right.t9 a_n3202_n3888# 0.313488f
C35 drain_right.n8 a_n3202_n3888# 2.83975f
C36 drain_right.t6 a_n3202_n3888# 0.313488f
C37 drain_right.t13 a_n3202_n3888# 0.313488f
C38 drain_right.n9 a_n3202_n3888# 2.83357f
C39 drain_right.n10 a_n3202_n3888# 0.769754f
C40 drain_right.t8 a_n3202_n3888# 0.313488f
C41 drain_right.t4 a_n3202_n3888# 0.313488f
C42 drain_right.n11 a_n3202_n3888# 2.83357f
C43 drain_right.n12 a_n3202_n3888# 0.382643f
C44 drain_right.t3 a_n3202_n3888# 0.313488f
C45 drain_right.t10 a_n3202_n3888# 0.313488f
C46 drain_right.n13 a_n3202_n3888# 2.83357f
C47 drain_right.n14 a_n3202_n3888# 0.382643f
C48 drain_right.t14 a_n3202_n3888# 0.313488f
C49 drain_right.t5 a_n3202_n3888# 0.313488f
C50 drain_right.n15 a_n3202_n3888# 2.83357f
C51 drain_right.n16 a_n3202_n3888# 0.619792f
C52 minus.n0 a_n3202_n3888# 0.037546f
C53 minus.n1 a_n3202_n3888# 0.00852f
C54 minus.t14 a_n3202_n3888# 1.28034f
C55 minus.n2 a_n3202_n3888# 0.062538f
C56 minus.t11 a_n3202_n3888# 1.28034f
C57 minus.n3 a_n3202_n3888# 0.490653f
C58 minus.n4 a_n3202_n3888# 0.037546f
C59 minus.t13 a_n3202_n3888# 1.28034f
C60 minus.n5 a_n3202_n3888# 0.501372f
C61 minus.n6 a_n3202_n3888# 0.172824f
C62 minus.t10 a_n3202_n3888# 1.30088f
C63 minus.n7 a_n3202_n3888# 0.475926f
C64 minus.t8 a_n3202_n3888# 1.28034f
C65 minus.n8 a_n3202_n3888# 0.493809f
C66 minus.n9 a_n3202_n3888# 0.00852f
C67 minus.t6 a_n3202_n3888# 1.28034f
C68 minus.n10 a_n3202_n3888# 0.500909f
C69 minus.n11 a_n3202_n3888# 0.062538f
C70 minus.n12 a_n3202_n3888# 0.062538f
C71 minus.n13 a_n3202_n3888# 0.050101f
C72 minus.n14 a_n3202_n3888# 0.00852f
C73 minus.t15 a_n3202_n3888# 1.28034f
C74 minus.n15 a_n3202_n3888# 0.490653f
C75 minus.n16 a_n3202_n3888# 0.00852f
C76 minus.n17 a_n3202_n3888# 0.037546f
C77 minus.n18 a_n3202_n3888# 0.037546f
C78 minus.n19 a_n3202_n3888# 0.050101f
C79 minus.n20 a_n3202_n3888# 0.00852f
C80 minus.t9 a_n3202_n3888# 1.28034f
C81 minus.n21 a_n3202_n3888# 0.501372f
C82 minus.t16 a_n3202_n3888# 1.28034f
C83 minus.n22 a_n3202_n3888# 0.500909f
C84 minus.n23 a_n3202_n3888# 0.062538f
C85 minus.n24 a_n3202_n3888# 0.050101f
C86 minus.n25 a_n3202_n3888# 0.037546f
C87 minus.n26 a_n3202_n3888# 0.490653f
C88 minus.n27 a_n3202_n3888# 0.00852f
C89 minus.t5 a_n3202_n3888# 1.28034f
C90 minus.n28 a_n3202_n3888# 0.490306f
C91 minus.n29 a_n3202_n3888# 1.76861f
C92 minus.n30 a_n3202_n3888# 0.037546f
C93 minus.n31 a_n3202_n3888# 0.00852f
C94 minus.n32 a_n3202_n3888# 0.062538f
C95 minus.t4 a_n3202_n3888# 1.28034f
C96 minus.n33 a_n3202_n3888# 0.490653f
C97 minus.n34 a_n3202_n3888# 0.037546f
C98 minus.t7 a_n3202_n3888# 1.28034f
C99 minus.n35 a_n3202_n3888# 0.501372f
C100 minus.n36 a_n3202_n3888# 0.172824f
C101 minus.t1 a_n3202_n3888# 1.30088f
C102 minus.n37 a_n3202_n3888# 0.475926f
C103 minus.t12 a_n3202_n3888# 1.28034f
C104 minus.n38 a_n3202_n3888# 0.493809f
C105 minus.n39 a_n3202_n3888# 0.00852f
C106 minus.t18 a_n3202_n3888# 1.28034f
C107 minus.n40 a_n3202_n3888# 0.500909f
C108 minus.n41 a_n3202_n3888# 0.062538f
C109 minus.n42 a_n3202_n3888# 0.062538f
C110 minus.n43 a_n3202_n3888# 0.050101f
C111 minus.n44 a_n3202_n3888# 0.00852f
C112 minus.t0 a_n3202_n3888# 1.28034f
C113 minus.n45 a_n3202_n3888# 0.490653f
C114 minus.n46 a_n3202_n3888# 0.00852f
C115 minus.n47 a_n3202_n3888# 0.037546f
C116 minus.n48 a_n3202_n3888# 0.037546f
C117 minus.n49 a_n3202_n3888# 0.050101f
C118 minus.n50 a_n3202_n3888# 0.00852f
C119 minus.t17 a_n3202_n3888# 1.28034f
C120 minus.n51 a_n3202_n3888# 0.501372f
C121 minus.t2 a_n3202_n3888# 1.28034f
C122 minus.n52 a_n3202_n3888# 0.500909f
C123 minus.n53 a_n3202_n3888# 0.062538f
C124 minus.n54 a_n3202_n3888# 0.050101f
C125 minus.n55 a_n3202_n3888# 0.037546f
C126 minus.t19 a_n3202_n3888# 1.28034f
C127 minus.n56 a_n3202_n3888# 0.490653f
C128 minus.n57 a_n3202_n3888# 0.00852f
C129 minus.t3 a_n3202_n3888# 1.28034f
C130 minus.n58 a_n3202_n3888# 0.490306f
C131 minus.n59 a_n3202_n3888# 0.263432f
C132 minus.n60 a_n3202_n3888# 2.09807f
C133 source.t33 a_n3202_n3888# 3.0981f
C134 source.n0 a_n3202_n3888# 1.48718f
C135 source.t28 a_n3202_n3888# 0.276453f
C136 source.t30 a_n3202_n3888# 0.276453f
C137 source.n1 a_n3202_n3888# 2.4284f
C138 source.n2 a_n3202_n3888# 0.376144f
C139 source.t26 a_n3202_n3888# 0.276453f
C140 source.t27 a_n3202_n3888# 0.276453f
C141 source.n3 a_n3202_n3888# 2.4284f
C142 source.n4 a_n3202_n3888# 0.376144f
C143 source.t25 a_n3202_n3888# 0.276453f
C144 source.t22 a_n3202_n3888# 0.276453f
C145 source.n5 a_n3202_n3888# 2.4284f
C146 source.n6 a_n3202_n3888# 0.376144f
C147 source.t21 a_n3202_n3888# 0.276453f
C148 source.t24 a_n3202_n3888# 0.276453f
C149 source.n7 a_n3202_n3888# 2.4284f
C150 source.n8 a_n3202_n3888# 0.376144f
C151 source.t19 a_n3202_n3888# 3.0981f
C152 source.n9 a_n3202_n3888# 0.42251f
C153 source.t39 a_n3202_n3888# 3.0981f
C154 source.n10 a_n3202_n3888# 0.42251f
C155 source.t10 a_n3202_n3888# 0.276453f
C156 source.t15 a_n3202_n3888# 0.276453f
C157 source.n11 a_n3202_n3888# 2.4284f
C158 source.n12 a_n3202_n3888# 0.376144f
C159 source.t0 a_n3202_n3888# 0.276453f
C160 source.t13 a_n3202_n3888# 0.276453f
C161 source.n13 a_n3202_n3888# 2.4284f
C162 source.n14 a_n3202_n3888# 0.376144f
C163 source.t16 a_n3202_n3888# 0.276453f
C164 source.t3 a_n3202_n3888# 0.276453f
C165 source.n15 a_n3202_n3888# 2.4284f
C166 source.n16 a_n3202_n3888# 0.376144f
C167 source.t14 a_n3202_n3888# 0.276453f
C168 source.t2 a_n3202_n3888# 0.276453f
C169 source.n17 a_n3202_n3888# 2.4284f
C170 source.n18 a_n3202_n3888# 0.376144f
C171 source.t8 a_n3202_n3888# 3.0981f
C172 source.n19 a_n3202_n3888# 1.88752f
C173 source.t38 a_n3202_n3888# 3.0981f
C174 source.n20 a_n3202_n3888# 1.88752f
C175 source.t31 a_n3202_n3888# 0.276453f
C176 source.t35 a_n3202_n3888# 0.276453f
C177 source.n21 a_n3202_n3888# 2.4284f
C178 source.n22 a_n3202_n3888# 0.376147f
C179 source.t29 a_n3202_n3888# 0.276453f
C180 source.t36 a_n3202_n3888# 0.276453f
C181 source.n23 a_n3202_n3888# 2.4284f
C182 source.n24 a_n3202_n3888# 0.376147f
C183 source.t23 a_n3202_n3888# 0.276453f
C184 source.t34 a_n3202_n3888# 0.276453f
C185 source.n25 a_n3202_n3888# 2.4284f
C186 source.n26 a_n3202_n3888# 0.376147f
C187 source.t20 a_n3202_n3888# 0.276453f
C188 source.t32 a_n3202_n3888# 0.276453f
C189 source.n27 a_n3202_n3888# 2.4284f
C190 source.n28 a_n3202_n3888# 0.376147f
C191 source.t37 a_n3202_n3888# 3.0981f
C192 source.n29 a_n3202_n3888# 0.422513f
C193 source.t5 a_n3202_n3888# 3.0981f
C194 source.n30 a_n3202_n3888# 0.422513f
C195 source.t11 a_n3202_n3888# 0.276453f
C196 source.t6 a_n3202_n3888# 0.276453f
C197 source.n31 a_n3202_n3888# 2.4284f
C198 source.n32 a_n3202_n3888# 0.376147f
C199 source.t12 a_n3202_n3888# 0.276453f
C200 source.t18 a_n3202_n3888# 0.276453f
C201 source.n33 a_n3202_n3888# 2.4284f
C202 source.n34 a_n3202_n3888# 0.376147f
C203 source.t4 a_n3202_n3888# 0.276453f
C204 source.t1 a_n3202_n3888# 0.276453f
C205 source.n35 a_n3202_n3888# 2.4284f
C206 source.n36 a_n3202_n3888# 0.376147f
C207 source.t9 a_n3202_n3888# 0.276453f
C208 source.t7 a_n3202_n3888# 0.276453f
C209 source.n37 a_n3202_n3888# 2.4284f
C210 source.n38 a_n3202_n3888# 0.376147f
C211 source.t17 a_n3202_n3888# 3.0981f
C212 source.n39 a_n3202_n3888# 0.579696f
C213 source.n40 a_n3202_n3888# 1.72475f
C214 drain_left.t4 a_n3202_n3888# 0.315611f
C215 drain_left.t12 a_n3202_n3888# 0.315611f
C216 drain_left.n0 a_n3202_n3888# 2.85899f
C217 drain_left.t17 a_n3202_n3888# 0.315611f
C218 drain_left.t19 a_n3202_n3888# 0.315611f
C219 drain_left.n1 a_n3202_n3888# 2.85275f
C220 drain_left.n2 a_n3202_n3888# 0.770884f
C221 drain_left.t2 a_n3202_n3888# 0.315611f
C222 drain_left.t8 a_n3202_n3888# 0.315611f
C223 drain_left.n3 a_n3202_n3888# 2.85275f
C224 drain_left.t5 a_n3202_n3888# 0.315611f
C225 drain_left.t3 a_n3202_n3888# 0.315611f
C226 drain_left.n4 a_n3202_n3888# 2.85899f
C227 drain_left.t16 a_n3202_n3888# 0.315611f
C228 drain_left.t9 a_n3202_n3888# 0.315611f
C229 drain_left.n5 a_n3202_n3888# 2.85275f
C230 drain_left.n6 a_n3202_n3888# 0.770884f
C231 drain_left.n7 a_n3202_n3888# 2.20343f
C232 drain_left.t15 a_n3202_n3888# 0.315611f
C233 drain_left.t10 a_n3202_n3888# 0.315611f
C234 drain_left.n8 a_n3202_n3888# 2.85899f
C235 drain_left.t0 a_n3202_n3888# 0.315611f
C236 drain_left.t1 a_n3202_n3888# 0.315611f
C237 drain_left.n9 a_n3202_n3888# 2.85275f
C238 drain_left.n10 a_n3202_n3888# 0.774956f
C239 drain_left.t7 a_n3202_n3888# 0.315611f
C240 drain_left.t13 a_n3202_n3888# 0.315611f
C241 drain_left.n11 a_n3202_n3888# 2.85275f
C242 drain_left.n12 a_n3202_n3888# 0.385234f
C243 drain_left.t14 a_n3202_n3888# 0.315611f
C244 drain_left.t18 a_n3202_n3888# 0.315611f
C245 drain_left.n13 a_n3202_n3888# 2.85275f
C246 drain_left.n14 a_n3202_n3888# 0.385234f
C247 drain_left.t11 a_n3202_n3888# 0.315611f
C248 drain_left.t6 a_n3202_n3888# 0.315611f
C249 drain_left.n15 a_n3202_n3888# 2.85274f
C250 drain_left.n16 a_n3202_n3888# 0.623998f
C251 plus.n0 a_n3202_n3888# 0.03798f
C252 plus.t5 a_n3202_n3888# 1.29512f
C253 plus.t8 a_n3202_n3888# 1.29512f
C254 plus.n1 a_n3202_n3888# 0.03798f
C255 plus.t10 a_n3202_n3888# 1.29512f
C256 plus.n2 a_n3202_n3888# 0.506692f
C257 plus.n3 a_n3202_n3888# 0.050679f
C258 plus.t11 a_n3202_n3888# 1.29512f
C259 plus.t12 a_n3202_n3888# 1.29512f
C260 plus.n4 a_n3202_n3888# 0.03798f
C261 plus.t16 a_n3202_n3888# 1.29512f
C262 plus.n5 a_n3202_n3888# 0.496318f
C263 plus.n6 a_n3202_n3888# 0.06326f
C264 plus.t13 a_n3202_n3888# 1.29512f
C265 plus.t14 a_n3202_n3888# 1.29512f
C266 plus.n7 a_n3202_n3888# 0.06326f
C267 plus.t17 a_n3202_n3888# 1.29512f
C268 plus.n8 a_n3202_n3888# 0.49951f
C269 plus.t19 a_n3202_n3888# 1.3159f
C270 plus.n9 a_n3202_n3888# 0.481421f
C271 plus.n10 a_n3202_n3888# 0.174819f
C272 plus.n11 a_n3202_n3888# 0.008618f
C273 plus.n12 a_n3202_n3888# 0.506692f
C274 plus.n13 a_n3202_n3888# 0.507161f
C275 plus.n14 a_n3202_n3888# 0.008618f
C276 plus.n15 a_n3202_n3888# 0.050679f
C277 plus.n16 a_n3202_n3888# 0.03798f
C278 plus.n17 a_n3202_n3888# 0.03798f
C279 plus.n18 a_n3202_n3888# 0.008618f
C280 plus.n19 a_n3202_n3888# 0.496318f
C281 plus.n20 a_n3202_n3888# 0.008618f
C282 plus.n21 a_n3202_n3888# 0.507161f
C283 plus.n22 a_n3202_n3888# 0.06326f
C284 plus.n23 a_n3202_n3888# 0.06326f
C285 plus.n24 a_n3202_n3888# 0.050679f
C286 plus.n25 a_n3202_n3888# 0.008618f
C287 plus.n26 a_n3202_n3888# 0.496318f
C288 plus.n27 a_n3202_n3888# 0.008618f
C289 plus.n28 a_n3202_n3888# 0.495966f
C290 plus.n29 a_n3202_n3888# 0.498202f
C291 plus.n30 a_n3202_n3888# 0.03798f
C292 plus.t0 a_n3202_n3888# 1.29512f
C293 plus.n31 a_n3202_n3888# 0.03798f
C294 plus.t7 a_n3202_n3888# 1.29512f
C295 plus.t3 a_n3202_n3888# 1.29512f
C296 plus.n32 a_n3202_n3888# 0.506692f
C297 plus.n33 a_n3202_n3888# 0.050679f
C298 plus.t9 a_n3202_n3888# 1.29512f
C299 plus.n34 a_n3202_n3888# 0.03798f
C300 plus.t2 a_n3202_n3888# 1.29512f
C301 plus.t15 a_n3202_n3888# 1.29512f
C302 plus.n35 a_n3202_n3888# 0.496318f
C303 plus.n36 a_n3202_n3888# 0.06326f
C304 plus.t4 a_n3202_n3888# 1.29512f
C305 plus.n37 a_n3202_n3888# 0.06326f
C306 plus.t18 a_n3202_n3888# 1.29512f
C307 plus.t6 a_n3202_n3888# 1.29512f
C308 plus.n38 a_n3202_n3888# 0.49951f
C309 plus.t1 a_n3202_n3888# 1.3159f
C310 plus.n39 a_n3202_n3888# 0.481421f
C311 plus.n40 a_n3202_n3888# 0.174819f
C312 plus.n41 a_n3202_n3888# 0.008618f
C313 plus.n42 a_n3202_n3888# 0.506692f
C314 plus.n43 a_n3202_n3888# 0.507161f
C315 plus.n44 a_n3202_n3888# 0.008618f
C316 plus.n45 a_n3202_n3888# 0.050679f
C317 plus.n46 a_n3202_n3888# 0.03798f
C318 plus.n47 a_n3202_n3888# 0.03798f
C319 plus.n48 a_n3202_n3888# 0.008618f
C320 plus.n49 a_n3202_n3888# 0.496318f
C321 plus.n50 a_n3202_n3888# 0.008618f
C322 plus.n51 a_n3202_n3888# 0.507161f
C323 plus.n52 a_n3202_n3888# 0.06326f
C324 plus.n53 a_n3202_n3888# 0.06326f
C325 plus.n54 a_n3202_n3888# 0.050679f
C326 plus.n55 a_n3202_n3888# 0.008618f
C327 plus.n56 a_n3202_n3888# 0.496318f
C328 plus.n57 a_n3202_n3888# 0.008618f
C329 plus.n58 a_n3202_n3888# 0.495966f
C330 plus.n59 a_n3202_n3888# 1.49876f
.ends

