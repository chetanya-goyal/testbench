* NGSPICE file created from diffpair478.ext - technology: sky130A

.subckt diffpair478 minus drain_right drain_left source plus
X0 drain_right.t19 minus.t0 source.t38 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X1 a_n3202_n3288# a_n3202_n3288# a_n3202_n3288# a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.8
X2 drain_right.t18 minus.t1 source.t22 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X3 source.t9 plus.t0 drain_left.t19 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X4 a_n3202_n3288# a_n3202_n3288# a_n3202_n3288# a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.8
X5 drain_right.t17 minus.t2 source.t25 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X6 drain_right.t16 minus.t3 source.t29 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X7 source.t6 plus.t1 drain_left.t18 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X8 a_n3202_n3288# a_n3202_n3288# a_n3202_n3288# a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.8
X9 source.t15 plus.t2 drain_left.t17 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X10 drain_left.t16 plus.t3 source.t7 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X11 source.t34 minus.t4 drain_right.t15 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
X12 drain_right.t14 minus.t5 source.t23 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X13 drain_left.t15 plus.t4 source.t1 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X14 drain_right.t13 minus.t6 source.t26 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X15 a_n3202_n3288# a_n3202_n3288# a_n3202_n3288# a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.8
X16 drain_left.t14 plus.t5 source.t17 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X17 source.t19 minus.t7 drain_right.t12 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X18 drain_right.t11 minus.t8 source.t32 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X19 drain_right.t10 minus.t9 source.t30 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X20 source.t8 plus.t6 drain_left.t13 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X21 source.t36 minus.t10 drain_right.t9 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X22 drain_left.t12 plus.t7 source.t0 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X23 drain_left.t11 plus.t8 source.t11 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X24 source.t35 minus.t11 drain_right.t8 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X25 drain_right.t7 minus.t12 source.t24 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X26 drain_left.t10 plus.t9 source.t18 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X27 drain_right.t6 minus.t13 source.t27 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X28 source.t21 minus.t14 drain_right.t5 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X29 source.t10 plus.t10 drain_left.t9 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X30 source.t20 minus.t15 drain_right.t4 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X31 source.t33 minus.t16 drain_right.t3 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X32 drain_left.t8 plus.t11 source.t14 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X33 drain_left.t7 plus.t12 source.t3 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X34 source.t31 minus.t17 drain_right.t2 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X35 source.t16 plus.t13 drain_left.t6 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X36 source.t13 plus.t14 drain_left.t5 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
X37 drain_left.t4 plus.t15 source.t39 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.8
X38 source.t4 plus.t16 drain_left.t3 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X39 drain_left.t2 plus.t17 source.t2 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X40 source.t37 minus.t18 drain_right.t1 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
X41 source.t12 plus.t18 drain_left.t1 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
X42 source.t28 minus.t19 drain_right.t0 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.8
X43 source.t5 plus.t19 drain_left.t0 a_n3202_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.8
R0 minus.n7 minus.t9 432.394
R1 minus.n37 minus.t19 432.394
R2 minus.n8 minus.t7 410.604
R3 minus.n10 minus.t6 410.604
R4 minus.n5 minus.t11 410.604
R5 minus.n15 minus.t13 410.604
R6 minus.n3 minus.t10 410.604
R7 minus.n21 minus.t8 410.604
R8 minus.n22 minus.t17 410.604
R9 minus.n26 minus.t12 410.604
R10 minus.n28 minus.t4 410.604
R11 minus.n38 minus.t5 410.604
R12 minus.n40 minus.t16 410.604
R13 minus.n35 minus.t3 410.604
R14 minus.n45 minus.t18 410.604
R15 minus.n33 minus.t2 410.604
R16 minus.n51 minus.t14 410.604
R17 minus.n52 minus.t0 410.604
R18 minus.n56 minus.t15 410.604
R19 minus.n58 minus.t1 410.604
R20 minus.n29 minus.n28 161.3
R21 minus.n27 minus.n0 161.3
R22 minus.n26 minus.n25 161.3
R23 minus.n24 minus.n1 161.3
R24 minus.n20 minus.n19 161.3
R25 minus.n18 minus.n3 161.3
R26 minus.n17 minus.n16 161.3
R27 minus.n15 minus.n4 161.3
R28 minus.n14 minus.n13 161.3
R29 minus.n9 minus.n6 161.3
R30 minus.n59 minus.n58 161.3
R31 minus.n57 minus.n30 161.3
R32 minus.n56 minus.n55 161.3
R33 minus.n54 minus.n31 161.3
R34 minus.n50 minus.n49 161.3
R35 minus.n48 minus.n33 161.3
R36 minus.n47 minus.n46 161.3
R37 minus.n45 minus.n34 161.3
R38 minus.n44 minus.n43 161.3
R39 minus.n39 minus.n36 161.3
R40 minus.n23 minus.n22 80.6037
R41 minus.n21 minus.n2 80.6037
R42 minus.n12 minus.n5 80.6037
R43 minus.n11 minus.n10 80.6037
R44 minus.n53 minus.n52 80.6037
R45 minus.n51 minus.n32 80.6037
R46 minus.n42 minus.n35 80.6037
R47 minus.n41 minus.n40 80.6037
R48 minus.n10 minus.n5 48.2005
R49 minus.n22 minus.n21 48.2005
R50 minus.n40 minus.n35 48.2005
R51 minus.n52 minus.n51 48.2005
R52 minus.n7 minus.n6 44.8565
R53 minus.n37 minus.n36 44.8565
R54 minus.n14 minus.n5 43.0884
R55 minus.n21 minus.n20 43.0884
R56 minus.n44 minus.n35 43.0884
R57 minus.n51 minus.n50 43.0884
R58 minus.n60 minus.n29 41.455
R59 minus.n10 minus.n9 40.1672
R60 minus.n22 minus.n1 40.1672
R61 minus.n40 minus.n39 40.1672
R62 minus.n52 minus.n31 40.1672
R63 minus.n28 minus.n27 27.0217
R64 minus.n58 minus.n57 27.0217
R65 minus.n16 minus.n3 24.1005
R66 minus.n16 minus.n15 24.1005
R67 minus.n46 minus.n45 24.1005
R68 minus.n46 minus.n33 24.1005
R69 minus.n27 minus.n26 21.1793
R70 minus.n57 minus.n56 21.1793
R71 minus.n8 minus.n7 20.1275
R72 minus.n38 minus.n37 20.1275
R73 minus.n9 minus.n8 8.03383
R74 minus.n26 minus.n1 8.03383
R75 minus.n39 minus.n38 8.03383
R76 minus.n56 minus.n31 8.03383
R77 minus.n60 minus.n59 6.70505
R78 minus.n15 minus.n14 5.11262
R79 minus.n20 minus.n3 5.11262
R80 minus.n45 minus.n44 5.11262
R81 minus.n50 minus.n33 5.11262
R82 minus.n23 minus.n2 0.380177
R83 minus.n12 minus.n11 0.380177
R84 minus.n42 minus.n41 0.380177
R85 minus.n53 minus.n32 0.380177
R86 minus.n24 minus.n23 0.285035
R87 minus.n19 minus.n2 0.285035
R88 minus.n13 minus.n12 0.285035
R89 minus.n11 minus.n6 0.285035
R90 minus.n41 minus.n36 0.285035
R91 minus.n43 minus.n42 0.285035
R92 minus.n49 minus.n32 0.285035
R93 minus.n54 minus.n53 0.285035
R94 minus.n29 minus.n0 0.189894
R95 minus.n25 minus.n0 0.189894
R96 minus.n25 minus.n24 0.189894
R97 minus.n19 minus.n18 0.189894
R98 minus.n18 minus.n17 0.189894
R99 minus.n17 minus.n4 0.189894
R100 minus.n13 minus.n4 0.189894
R101 minus.n43 minus.n34 0.189894
R102 minus.n47 minus.n34 0.189894
R103 minus.n48 minus.n47 0.189894
R104 minus.n49 minus.n48 0.189894
R105 minus.n55 minus.n54 0.189894
R106 minus.n55 minus.n30 0.189894
R107 minus.n59 minus.n30 0.189894
R108 minus minus.n60 0.188
R109 source.n554 source.n494 289.615
R110 source.n480 source.n420 289.615
R111 source.n414 source.n354 289.615
R112 source.n340 source.n280 289.615
R113 source.n60 source.n0 289.615
R114 source.n134 source.n74 289.615
R115 source.n200 source.n140 289.615
R116 source.n274 source.n214 289.615
R117 source.n514 source.n513 185
R118 source.n519 source.n518 185
R119 source.n521 source.n520 185
R120 source.n510 source.n509 185
R121 source.n527 source.n526 185
R122 source.n529 source.n528 185
R123 source.n506 source.n505 185
R124 source.n536 source.n535 185
R125 source.n537 source.n504 185
R126 source.n539 source.n538 185
R127 source.n502 source.n501 185
R128 source.n545 source.n544 185
R129 source.n547 source.n546 185
R130 source.n498 source.n497 185
R131 source.n553 source.n552 185
R132 source.n555 source.n554 185
R133 source.n440 source.n439 185
R134 source.n445 source.n444 185
R135 source.n447 source.n446 185
R136 source.n436 source.n435 185
R137 source.n453 source.n452 185
R138 source.n455 source.n454 185
R139 source.n432 source.n431 185
R140 source.n462 source.n461 185
R141 source.n463 source.n430 185
R142 source.n465 source.n464 185
R143 source.n428 source.n427 185
R144 source.n471 source.n470 185
R145 source.n473 source.n472 185
R146 source.n424 source.n423 185
R147 source.n479 source.n478 185
R148 source.n481 source.n480 185
R149 source.n374 source.n373 185
R150 source.n379 source.n378 185
R151 source.n381 source.n380 185
R152 source.n370 source.n369 185
R153 source.n387 source.n386 185
R154 source.n389 source.n388 185
R155 source.n366 source.n365 185
R156 source.n396 source.n395 185
R157 source.n397 source.n364 185
R158 source.n399 source.n398 185
R159 source.n362 source.n361 185
R160 source.n405 source.n404 185
R161 source.n407 source.n406 185
R162 source.n358 source.n357 185
R163 source.n413 source.n412 185
R164 source.n415 source.n414 185
R165 source.n300 source.n299 185
R166 source.n305 source.n304 185
R167 source.n307 source.n306 185
R168 source.n296 source.n295 185
R169 source.n313 source.n312 185
R170 source.n315 source.n314 185
R171 source.n292 source.n291 185
R172 source.n322 source.n321 185
R173 source.n323 source.n290 185
R174 source.n325 source.n324 185
R175 source.n288 source.n287 185
R176 source.n331 source.n330 185
R177 source.n333 source.n332 185
R178 source.n284 source.n283 185
R179 source.n339 source.n338 185
R180 source.n341 source.n340 185
R181 source.n61 source.n60 185
R182 source.n59 source.n58 185
R183 source.n4 source.n3 185
R184 source.n53 source.n52 185
R185 source.n51 source.n50 185
R186 source.n8 source.n7 185
R187 source.n45 source.n44 185
R188 source.n43 source.n10 185
R189 source.n42 source.n41 185
R190 source.n13 source.n11 185
R191 source.n36 source.n35 185
R192 source.n34 source.n33 185
R193 source.n17 source.n16 185
R194 source.n28 source.n27 185
R195 source.n26 source.n25 185
R196 source.n21 source.n20 185
R197 source.n135 source.n134 185
R198 source.n133 source.n132 185
R199 source.n78 source.n77 185
R200 source.n127 source.n126 185
R201 source.n125 source.n124 185
R202 source.n82 source.n81 185
R203 source.n119 source.n118 185
R204 source.n117 source.n84 185
R205 source.n116 source.n115 185
R206 source.n87 source.n85 185
R207 source.n110 source.n109 185
R208 source.n108 source.n107 185
R209 source.n91 source.n90 185
R210 source.n102 source.n101 185
R211 source.n100 source.n99 185
R212 source.n95 source.n94 185
R213 source.n201 source.n200 185
R214 source.n199 source.n198 185
R215 source.n144 source.n143 185
R216 source.n193 source.n192 185
R217 source.n191 source.n190 185
R218 source.n148 source.n147 185
R219 source.n185 source.n184 185
R220 source.n183 source.n150 185
R221 source.n182 source.n181 185
R222 source.n153 source.n151 185
R223 source.n176 source.n175 185
R224 source.n174 source.n173 185
R225 source.n157 source.n156 185
R226 source.n168 source.n167 185
R227 source.n166 source.n165 185
R228 source.n161 source.n160 185
R229 source.n275 source.n274 185
R230 source.n273 source.n272 185
R231 source.n218 source.n217 185
R232 source.n267 source.n266 185
R233 source.n265 source.n264 185
R234 source.n222 source.n221 185
R235 source.n259 source.n258 185
R236 source.n257 source.n224 185
R237 source.n256 source.n255 185
R238 source.n227 source.n225 185
R239 source.n250 source.n249 185
R240 source.n248 source.n247 185
R241 source.n231 source.n230 185
R242 source.n242 source.n241 185
R243 source.n240 source.n239 185
R244 source.n235 source.n234 185
R245 source.n515 source.t22 149.524
R246 source.n441 source.t28 149.524
R247 source.n375 source.t39 149.524
R248 source.n301 source.t13 149.524
R249 source.n22 source.t17 149.524
R250 source.n96 source.t12 149.524
R251 source.n162 source.t30 149.524
R252 source.n236 source.t34 149.524
R253 source.n519 source.n513 104.615
R254 source.n520 source.n519 104.615
R255 source.n520 source.n509 104.615
R256 source.n527 source.n509 104.615
R257 source.n528 source.n527 104.615
R258 source.n528 source.n505 104.615
R259 source.n536 source.n505 104.615
R260 source.n537 source.n536 104.615
R261 source.n538 source.n537 104.615
R262 source.n538 source.n501 104.615
R263 source.n545 source.n501 104.615
R264 source.n546 source.n545 104.615
R265 source.n546 source.n497 104.615
R266 source.n553 source.n497 104.615
R267 source.n554 source.n553 104.615
R268 source.n445 source.n439 104.615
R269 source.n446 source.n445 104.615
R270 source.n446 source.n435 104.615
R271 source.n453 source.n435 104.615
R272 source.n454 source.n453 104.615
R273 source.n454 source.n431 104.615
R274 source.n462 source.n431 104.615
R275 source.n463 source.n462 104.615
R276 source.n464 source.n463 104.615
R277 source.n464 source.n427 104.615
R278 source.n471 source.n427 104.615
R279 source.n472 source.n471 104.615
R280 source.n472 source.n423 104.615
R281 source.n479 source.n423 104.615
R282 source.n480 source.n479 104.615
R283 source.n379 source.n373 104.615
R284 source.n380 source.n379 104.615
R285 source.n380 source.n369 104.615
R286 source.n387 source.n369 104.615
R287 source.n388 source.n387 104.615
R288 source.n388 source.n365 104.615
R289 source.n396 source.n365 104.615
R290 source.n397 source.n396 104.615
R291 source.n398 source.n397 104.615
R292 source.n398 source.n361 104.615
R293 source.n405 source.n361 104.615
R294 source.n406 source.n405 104.615
R295 source.n406 source.n357 104.615
R296 source.n413 source.n357 104.615
R297 source.n414 source.n413 104.615
R298 source.n305 source.n299 104.615
R299 source.n306 source.n305 104.615
R300 source.n306 source.n295 104.615
R301 source.n313 source.n295 104.615
R302 source.n314 source.n313 104.615
R303 source.n314 source.n291 104.615
R304 source.n322 source.n291 104.615
R305 source.n323 source.n322 104.615
R306 source.n324 source.n323 104.615
R307 source.n324 source.n287 104.615
R308 source.n331 source.n287 104.615
R309 source.n332 source.n331 104.615
R310 source.n332 source.n283 104.615
R311 source.n339 source.n283 104.615
R312 source.n340 source.n339 104.615
R313 source.n60 source.n59 104.615
R314 source.n59 source.n3 104.615
R315 source.n52 source.n3 104.615
R316 source.n52 source.n51 104.615
R317 source.n51 source.n7 104.615
R318 source.n44 source.n7 104.615
R319 source.n44 source.n43 104.615
R320 source.n43 source.n42 104.615
R321 source.n42 source.n11 104.615
R322 source.n35 source.n11 104.615
R323 source.n35 source.n34 104.615
R324 source.n34 source.n16 104.615
R325 source.n27 source.n16 104.615
R326 source.n27 source.n26 104.615
R327 source.n26 source.n20 104.615
R328 source.n134 source.n133 104.615
R329 source.n133 source.n77 104.615
R330 source.n126 source.n77 104.615
R331 source.n126 source.n125 104.615
R332 source.n125 source.n81 104.615
R333 source.n118 source.n81 104.615
R334 source.n118 source.n117 104.615
R335 source.n117 source.n116 104.615
R336 source.n116 source.n85 104.615
R337 source.n109 source.n85 104.615
R338 source.n109 source.n108 104.615
R339 source.n108 source.n90 104.615
R340 source.n101 source.n90 104.615
R341 source.n101 source.n100 104.615
R342 source.n100 source.n94 104.615
R343 source.n200 source.n199 104.615
R344 source.n199 source.n143 104.615
R345 source.n192 source.n143 104.615
R346 source.n192 source.n191 104.615
R347 source.n191 source.n147 104.615
R348 source.n184 source.n147 104.615
R349 source.n184 source.n183 104.615
R350 source.n183 source.n182 104.615
R351 source.n182 source.n151 104.615
R352 source.n175 source.n151 104.615
R353 source.n175 source.n174 104.615
R354 source.n174 source.n156 104.615
R355 source.n167 source.n156 104.615
R356 source.n167 source.n166 104.615
R357 source.n166 source.n160 104.615
R358 source.n274 source.n273 104.615
R359 source.n273 source.n217 104.615
R360 source.n266 source.n217 104.615
R361 source.n266 source.n265 104.615
R362 source.n265 source.n221 104.615
R363 source.n258 source.n221 104.615
R364 source.n258 source.n257 104.615
R365 source.n257 source.n256 104.615
R366 source.n256 source.n225 104.615
R367 source.n249 source.n225 104.615
R368 source.n249 source.n248 104.615
R369 source.n248 source.n230 104.615
R370 source.n241 source.n230 104.615
R371 source.n241 source.n240 104.615
R372 source.n240 source.n234 104.615
R373 source.t22 source.n513 52.3082
R374 source.t28 source.n439 52.3082
R375 source.t39 source.n373 52.3082
R376 source.t13 source.n299 52.3082
R377 source.t17 source.n20 52.3082
R378 source.t12 source.n94 52.3082
R379 source.t30 source.n160 52.3082
R380 source.t34 source.n234 52.3082
R381 source.n67 source.n66 42.8739
R382 source.n69 source.n68 42.8739
R383 source.n71 source.n70 42.8739
R384 source.n73 source.n72 42.8739
R385 source.n207 source.n206 42.8739
R386 source.n209 source.n208 42.8739
R387 source.n211 source.n210 42.8739
R388 source.n213 source.n212 42.8739
R389 source.n493 source.n492 42.8737
R390 source.n491 source.n490 42.8737
R391 source.n489 source.n488 42.8737
R392 source.n487 source.n486 42.8737
R393 source.n353 source.n352 42.8737
R394 source.n351 source.n350 42.8737
R395 source.n349 source.n348 42.8737
R396 source.n347 source.n346 42.8737
R397 source.n559 source.n558 29.8581
R398 source.n485 source.n484 29.8581
R399 source.n419 source.n418 29.8581
R400 source.n345 source.n344 29.8581
R401 source.n65 source.n64 29.8581
R402 source.n139 source.n138 29.8581
R403 source.n205 source.n204 29.8581
R404 source.n279 source.n278 29.8581
R405 source.n345 source.n279 22.2619
R406 source.n560 source.n65 16.5119
R407 source.n539 source.n504 13.1884
R408 source.n465 source.n430 13.1884
R409 source.n399 source.n364 13.1884
R410 source.n325 source.n290 13.1884
R411 source.n45 source.n10 13.1884
R412 source.n119 source.n84 13.1884
R413 source.n185 source.n150 13.1884
R414 source.n259 source.n224 13.1884
R415 source.n535 source.n534 12.8005
R416 source.n540 source.n502 12.8005
R417 source.n461 source.n460 12.8005
R418 source.n466 source.n428 12.8005
R419 source.n395 source.n394 12.8005
R420 source.n400 source.n362 12.8005
R421 source.n321 source.n320 12.8005
R422 source.n326 source.n288 12.8005
R423 source.n46 source.n8 12.8005
R424 source.n41 source.n12 12.8005
R425 source.n120 source.n82 12.8005
R426 source.n115 source.n86 12.8005
R427 source.n186 source.n148 12.8005
R428 source.n181 source.n152 12.8005
R429 source.n260 source.n222 12.8005
R430 source.n255 source.n226 12.8005
R431 source.n533 source.n506 12.0247
R432 source.n544 source.n543 12.0247
R433 source.n459 source.n432 12.0247
R434 source.n470 source.n469 12.0247
R435 source.n393 source.n366 12.0247
R436 source.n404 source.n403 12.0247
R437 source.n319 source.n292 12.0247
R438 source.n330 source.n329 12.0247
R439 source.n50 source.n49 12.0247
R440 source.n40 source.n13 12.0247
R441 source.n124 source.n123 12.0247
R442 source.n114 source.n87 12.0247
R443 source.n190 source.n189 12.0247
R444 source.n180 source.n153 12.0247
R445 source.n264 source.n263 12.0247
R446 source.n254 source.n227 12.0247
R447 source.n530 source.n529 11.249
R448 source.n547 source.n500 11.249
R449 source.n456 source.n455 11.249
R450 source.n473 source.n426 11.249
R451 source.n390 source.n389 11.249
R452 source.n407 source.n360 11.249
R453 source.n316 source.n315 11.249
R454 source.n333 source.n286 11.249
R455 source.n53 source.n6 11.249
R456 source.n37 source.n36 11.249
R457 source.n127 source.n80 11.249
R458 source.n111 source.n110 11.249
R459 source.n193 source.n146 11.249
R460 source.n177 source.n176 11.249
R461 source.n267 source.n220 11.249
R462 source.n251 source.n250 11.249
R463 source.n526 source.n508 10.4732
R464 source.n548 source.n498 10.4732
R465 source.n452 source.n434 10.4732
R466 source.n474 source.n424 10.4732
R467 source.n386 source.n368 10.4732
R468 source.n408 source.n358 10.4732
R469 source.n312 source.n294 10.4732
R470 source.n334 source.n284 10.4732
R471 source.n54 source.n4 10.4732
R472 source.n33 source.n15 10.4732
R473 source.n128 source.n78 10.4732
R474 source.n107 source.n89 10.4732
R475 source.n194 source.n144 10.4732
R476 source.n173 source.n155 10.4732
R477 source.n268 source.n218 10.4732
R478 source.n247 source.n229 10.4732
R479 source.n515 source.n514 10.2747
R480 source.n441 source.n440 10.2747
R481 source.n375 source.n374 10.2747
R482 source.n301 source.n300 10.2747
R483 source.n22 source.n21 10.2747
R484 source.n96 source.n95 10.2747
R485 source.n162 source.n161 10.2747
R486 source.n236 source.n235 10.2747
R487 source.n525 source.n510 9.69747
R488 source.n552 source.n551 9.69747
R489 source.n451 source.n436 9.69747
R490 source.n478 source.n477 9.69747
R491 source.n385 source.n370 9.69747
R492 source.n412 source.n411 9.69747
R493 source.n311 source.n296 9.69747
R494 source.n338 source.n337 9.69747
R495 source.n58 source.n57 9.69747
R496 source.n32 source.n17 9.69747
R497 source.n132 source.n131 9.69747
R498 source.n106 source.n91 9.69747
R499 source.n198 source.n197 9.69747
R500 source.n172 source.n157 9.69747
R501 source.n272 source.n271 9.69747
R502 source.n246 source.n231 9.69747
R503 source.n558 source.n557 9.45567
R504 source.n484 source.n483 9.45567
R505 source.n418 source.n417 9.45567
R506 source.n344 source.n343 9.45567
R507 source.n64 source.n63 9.45567
R508 source.n138 source.n137 9.45567
R509 source.n204 source.n203 9.45567
R510 source.n278 source.n277 9.45567
R511 source.n557 source.n556 9.3005
R512 source.n496 source.n495 9.3005
R513 source.n551 source.n550 9.3005
R514 source.n549 source.n548 9.3005
R515 source.n500 source.n499 9.3005
R516 source.n543 source.n542 9.3005
R517 source.n541 source.n540 9.3005
R518 source.n517 source.n516 9.3005
R519 source.n512 source.n511 9.3005
R520 source.n523 source.n522 9.3005
R521 source.n525 source.n524 9.3005
R522 source.n508 source.n507 9.3005
R523 source.n531 source.n530 9.3005
R524 source.n533 source.n532 9.3005
R525 source.n534 source.n503 9.3005
R526 source.n483 source.n482 9.3005
R527 source.n422 source.n421 9.3005
R528 source.n477 source.n476 9.3005
R529 source.n475 source.n474 9.3005
R530 source.n426 source.n425 9.3005
R531 source.n469 source.n468 9.3005
R532 source.n467 source.n466 9.3005
R533 source.n443 source.n442 9.3005
R534 source.n438 source.n437 9.3005
R535 source.n449 source.n448 9.3005
R536 source.n451 source.n450 9.3005
R537 source.n434 source.n433 9.3005
R538 source.n457 source.n456 9.3005
R539 source.n459 source.n458 9.3005
R540 source.n460 source.n429 9.3005
R541 source.n417 source.n416 9.3005
R542 source.n356 source.n355 9.3005
R543 source.n411 source.n410 9.3005
R544 source.n409 source.n408 9.3005
R545 source.n360 source.n359 9.3005
R546 source.n403 source.n402 9.3005
R547 source.n401 source.n400 9.3005
R548 source.n377 source.n376 9.3005
R549 source.n372 source.n371 9.3005
R550 source.n383 source.n382 9.3005
R551 source.n385 source.n384 9.3005
R552 source.n368 source.n367 9.3005
R553 source.n391 source.n390 9.3005
R554 source.n393 source.n392 9.3005
R555 source.n394 source.n363 9.3005
R556 source.n343 source.n342 9.3005
R557 source.n282 source.n281 9.3005
R558 source.n337 source.n336 9.3005
R559 source.n335 source.n334 9.3005
R560 source.n286 source.n285 9.3005
R561 source.n329 source.n328 9.3005
R562 source.n327 source.n326 9.3005
R563 source.n303 source.n302 9.3005
R564 source.n298 source.n297 9.3005
R565 source.n309 source.n308 9.3005
R566 source.n311 source.n310 9.3005
R567 source.n294 source.n293 9.3005
R568 source.n317 source.n316 9.3005
R569 source.n319 source.n318 9.3005
R570 source.n320 source.n289 9.3005
R571 source.n24 source.n23 9.3005
R572 source.n19 source.n18 9.3005
R573 source.n30 source.n29 9.3005
R574 source.n32 source.n31 9.3005
R575 source.n15 source.n14 9.3005
R576 source.n38 source.n37 9.3005
R577 source.n40 source.n39 9.3005
R578 source.n12 source.n9 9.3005
R579 source.n63 source.n62 9.3005
R580 source.n2 source.n1 9.3005
R581 source.n57 source.n56 9.3005
R582 source.n55 source.n54 9.3005
R583 source.n6 source.n5 9.3005
R584 source.n49 source.n48 9.3005
R585 source.n47 source.n46 9.3005
R586 source.n98 source.n97 9.3005
R587 source.n93 source.n92 9.3005
R588 source.n104 source.n103 9.3005
R589 source.n106 source.n105 9.3005
R590 source.n89 source.n88 9.3005
R591 source.n112 source.n111 9.3005
R592 source.n114 source.n113 9.3005
R593 source.n86 source.n83 9.3005
R594 source.n137 source.n136 9.3005
R595 source.n76 source.n75 9.3005
R596 source.n131 source.n130 9.3005
R597 source.n129 source.n128 9.3005
R598 source.n80 source.n79 9.3005
R599 source.n123 source.n122 9.3005
R600 source.n121 source.n120 9.3005
R601 source.n164 source.n163 9.3005
R602 source.n159 source.n158 9.3005
R603 source.n170 source.n169 9.3005
R604 source.n172 source.n171 9.3005
R605 source.n155 source.n154 9.3005
R606 source.n178 source.n177 9.3005
R607 source.n180 source.n179 9.3005
R608 source.n152 source.n149 9.3005
R609 source.n203 source.n202 9.3005
R610 source.n142 source.n141 9.3005
R611 source.n197 source.n196 9.3005
R612 source.n195 source.n194 9.3005
R613 source.n146 source.n145 9.3005
R614 source.n189 source.n188 9.3005
R615 source.n187 source.n186 9.3005
R616 source.n238 source.n237 9.3005
R617 source.n233 source.n232 9.3005
R618 source.n244 source.n243 9.3005
R619 source.n246 source.n245 9.3005
R620 source.n229 source.n228 9.3005
R621 source.n252 source.n251 9.3005
R622 source.n254 source.n253 9.3005
R623 source.n226 source.n223 9.3005
R624 source.n277 source.n276 9.3005
R625 source.n216 source.n215 9.3005
R626 source.n271 source.n270 9.3005
R627 source.n269 source.n268 9.3005
R628 source.n220 source.n219 9.3005
R629 source.n263 source.n262 9.3005
R630 source.n261 source.n260 9.3005
R631 source.n522 source.n521 8.92171
R632 source.n555 source.n496 8.92171
R633 source.n448 source.n447 8.92171
R634 source.n481 source.n422 8.92171
R635 source.n382 source.n381 8.92171
R636 source.n415 source.n356 8.92171
R637 source.n308 source.n307 8.92171
R638 source.n341 source.n282 8.92171
R639 source.n61 source.n2 8.92171
R640 source.n29 source.n28 8.92171
R641 source.n135 source.n76 8.92171
R642 source.n103 source.n102 8.92171
R643 source.n201 source.n142 8.92171
R644 source.n169 source.n168 8.92171
R645 source.n275 source.n216 8.92171
R646 source.n243 source.n242 8.92171
R647 source.n518 source.n512 8.14595
R648 source.n556 source.n494 8.14595
R649 source.n444 source.n438 8.14595
R650 source.n482 source.n420 8.14595
R651 source.n378 source.n372 8.14595
R652 source.n416 source.n354 8.14595
R653 source.n304 source.n298 8.14595
R654 source.n342 source.n280 8.14595
R655 source.n62 source.n0 8.14595
R656 source.n25 source.n19 8.14595
R657 source.n136 source.n74 8.14595
R658 source.n99 source.n93 8.14595
R659 source.n202 source.n140 8.14595
R660 source.n165 source.n159 8.14595
R661 source.n276 source.n214 8.14595
R662 source.n239 source.n233 8.14595
R663 source.n517 source.n514 7.3702
R664 source.n443 source.n440 7.3702
R665 source.n377 source.n374 7.3702
R666 source.n303 source.n300 7.3702
R667 source.n24 source.n21 7.3702
R668 source.n98 source.n95 7.3702
R669 source.n164 source.n161 7.3702
R670 source.n238 source.n235 7.3702
R671 source.n518 source.n517 5.81868
R672 source.n558 source.n494 5.81868
R673 source.n444 source.n443 5.81868
R674 source.n484 source.n420 5.81868
R675 source.n378 source.n377 5.81868
R676 source.n418 source.n354 5.81868
R677 source.n304 source.n303 5.81868
R678 source.n344 source.n280 5.81868
R679 source.n64 source.n0 5.81868
R680 source.n25 source.n24 5.81868
R681 source.n138 source.n74 5.81868
R682 source.n99 source.n98 5.81868
R683 source.n204 source.n140 5.81868
R684 source.n165 source.n164 5.81868
R685 source.n278 source.n214 5.81868
R686 source.n239 source.n238 5.81868
R687 source.n560 source.n559 5.7505
R688 source.n521 source.n512 5.04292
R689 source.n556 source.n555 5.04292
R690 source.n447 source.n438 5.04292
R691 source.n482 source.n481 5.04292
R692 source.n381 source.n372 5.04292
R693 source.n416 source.n415 5.04292
R694 source.n307 source.n298 5.04292
R695 source.n342 source.n341 5.04292
R696 source.n62 source.n61 5.04292
R697 source.n28 source.n19 5.04292
R698 source.n136 source.n135 5.04292
R699 source.n102 source.n93 5.04292
R700 source.n202 source.n201 5.04292
R701 source.n168 source.n159 5.04292
R702 source.n276 source.n275 5.04292
R703 source.n242 source.n233 5.04292
R704 source.n522 source.n510 4.26717
R705 source.n552 source.n496 4.26717
R706 source.n448 source.n436 4.26717
R707 source.n478 source.n422 4.26717
R708 source.n382 source.n370 4.26717
R709 source.n412 source.n356 4.26717
R710 source.n308 source.n296 4.26717
R711 source.n338 source.n282 4.26717
R712 source.n58 source.n2 4.26717
R713 source.n29 source.n17 4.26717
R714 source.n132 source.n76 4.26717
R715 source.n103 source.n91 4.26717
R716 source.n198 source.n142 4.26717
R717 source.n169 source.n157 4.26717
R718 source.n272 source.n216 4.26717
R719 source.n243 source.n231 4.26717
R720 source.n526 source.n525 3.49141
R721 source.n551 source.n498 3.49141
R722 source.n452 source.n451 3.49141
R723 source.n477 source.n424 3.49141
R724 source.n386 source.n385 3.49141
R725 source.n411 source.n358 3.49141
R726 source.n312 source.n311 3.49141
R727 source.n337 source.n284 3.49141
R728 source.n57 source.n4 3.49141
R729 source.n33 source.n32 3.49141
R730 source.n131 source.n78 3.49141
R731 source.n107 source.n106 3.49141
R732 source.n197 source.n144 3.49141
R733 source.n173 source.n172 3.49141
R734 source.n271 source.n218 3.49141
R735 source.n247 source.n246 3.49141
R736 source.n516 source.n515 2.84303
R737 source.n442 source.n441 2.84303
R738 source.n376 source.n375 2.84303
R739 source.n302 source.n301 2.84303
R740 source.n23 source.n22 2.84303
R741 source.n97 source.n96 2.84303
R742 source.n163 source.n162 2.84303
R743 source.n237 source.n236 2.84303
R744 source.n529 source.n508 2.71565
R745 source.n548 source.n547 2.71565
R746 source.n455 source.n434 2.71565
R747 source.n474 source.n473 2.71565
R748 source.n389 source.n368 2.71565
R749 source.n408 source.n407 2.71565
R750 source.n315 source.n294 2.71565
R751 source.n334 source.n333 2.71565
R752 source.n54 source.n53 2.71565
R753 source.n36 source.n15 2.71565
R754 source.n128 source.n127 2.71565
R755 source.n110 source.n89 2.71565
R756 source.n194 source.n193 2.71565
R757 source.n176 source.n155 2.71565
R758 source.n268 source.n267 2.71565
R759 source.n250 source.n229 2.71565
R760 source.n530 source.n506 1.93989
R761 source.n544 source.n500 1.93989
R762 source.n456 source.n432 1.93989
R763 source.n470 source.n426 1.93989
R764 source.n390 source.n366 1.93989
R765 source.n404 source.n360 1.93989
R766 source.n316 source.n292 1.93989
R767 source.n330 source.n286 1.93989
R768 source.n50 source.n6 1.93989
R769 source.n37 source.n13 1.93989
R770 source.n124 source.n80 1.93989
R771 source.n111 source.n87 1.93989
R772 source.n190 source.n146 1.93989
R773 source.n177 source.n153 1.93989
R774 source.n264 source.n220 1.93989
R775 source.n251 source.n227 1.93989
R776 source.n492 source.t38 1.6505
R777 source.n492 source.t20 1.6505
R778 source.n490 source.t25 1.6505
R779 source.n490 source.t21 1.6505
R780 source.n488 source.t29 1.6505
R781 source.n488 source.t37 1.6505
R782 source.n486 source.t23 1.6505
R783 source.n486 source.t33 1.6505
R784 source.n352 source.t18 1.6505
R785 source.n352 source.t15 1.6505
R786 source.n350 source.t0 1.6505
R787 source.n350 source.t6 1.6505
R788 source.n348 source.t1 1.6505
R789 source.n348 source.t5 1.6505
R790 source.n346 source.t7 1.6505
R791 source.n346 source.t9 1.6505
R792 source.n66 source.t11 1.6505
R793 source.n66 source.t8 1.6505
R794 source.n68 source.t14 1.6505
R795 source.n68 source.t10 1.6505
R796 source.n70 source.t3 1.6505
R797 source.n70 source.t4 1.6505
R798 source.n72 source.t2 1.6505
R799 source.n72 source.t16 1.6505
R800 source.n206 source.t26 1.6505
R801 source.n206 source.t19 1.6505
R802 source.n208 source.t27 1.6505
R803 source.n208 source.t35 1.6505
R804 source.n210 source.t32 1.6505
R805 source.n210 source.t36 1.6505
R806 source.n212 source.t24 1.6505
R807 source.n212 source.t31 1.6505
R808 source.n535 source.n533 1.16414
R809 source.n543 source.n502 1.16414
R810 source.n461 source.n459 1.16414
R811 source.n469 source.n428 1.16414
R812 source.n395 source.n393 1.16414
R813 source.n403 source.n362 1.16414
R814 source.n321 source.n319 1.16414
R815 source.n329 source.n288 1.16414
R816 source.n49 source.n8 1.16414
R817 source.n41 source.n40 1.16414
R818 source.n123 source.n82 1.16414
R819 source.n115 source.n114 1.16414
R820 source.n189 source.n148 1.16414
R821 source.n181 source.n180 1.16414
R822 source.n263 source.n222 1.16414
R823 source.n255 source.n254 1.16414
R824 source.n279 source.n213 0.974638
R825 source.n213 source.n211 0.974638
R826 source.n211 source.n209 0.974638
R827 source.n209 source.n207 0.974638
R828 source.n207 source.n205 0.974638
R829 source.n139 source.n73 0.974638
R830 source.n73 source.n71 0.974638
R831 source.n71 source.n69 0.974638
R832 source.n69 source.n67 0.974638
R833 source.n67 source.n65 0.974638
R834 source.n347 source.n345 0.974638
R835 source.n349 source.n347 0.974638
R836 source.n351 source.n349 0.974638
R837 source.n353 source.n351 0.974638
R838 source.n419 source.n353 0.974638
R839 source.n487 source.n485 0.974638
R840 source.n489 source.n487 0.974638
R841 source.n491 source.n489 0.974638
R842 source.n493 source.n491 0.974638
R843 source.n559 source.n493 0.974638
R844 source.n205 source.n139 0.470328
R845 source.n485 source.n419 0.470328
R846 source.n534 source.n504 0.388379
R847 source.n540 source.n539 0.388379
R848 source.n460 source.n430 0.388379
R849 source.n466 source.n465 0.388379
R850 source.n394 source.n364 0.388379
R851 source.n400 source.n399 0.388379
R852 source.n320 source.n290 0.388379
R853 source.n326 source.n325 0.388379
R854 source.n46 source.n45 0.388379
R855 source.n12 source.n10 0.388379
R856 source.n120 source.n119 0.388379
R857 source.n86 source.n84 0.388379
R858 source.n186 source.n185 0.388379
R859 source.n152 source.n150 0.388379
R860 source.n260 source.n259 0.388379
R861 source.n226 source.n224 0.388379
R862 source source.n560 0.188
R863 source.n516 source.n511 0.155672
R864 source.n523 source.n511 0.155672
R865 source.n524 source.n523 0.155672
R866 source.n524 source.n507 0.155672
R867 source.n531 source.n507 0.155672
R868 source.n532 source.n531 0.155672
R869 source.n532 source.n503 0.155672
R870 source.n541 source.n503 0.155672
R871 source.n542 source.n541 0.155672
R872 source.n542 source.n499 0.155672
R873 source.n549 source.n499 0.155672
R874 source.n550 source.n549 0.155672
R875 source.n550 source.n495 0.155672
R876 source.n557 source.n495 0.155672
R877 source.n442 source.n437 0.155672
R878 source.n449 source.n437 0.155672
R879 source.n450 source.n449 0.155672
R880 source.n450 source.n433 0.155672
R881 source.n457 source.n433 0.155672
R882 source.n458 source.n457 0.155672
R883 source.n458 source.n429 0.155672
R884 source.n467 source.n429 0.155672
R885 source.n468 source.n467 0.155672
R886 source.n468 source.n425 0.155672
R887 source.n475 source.n425 0.155672
R888 source.n476 source.n475 0.155672
R889 source.n476 source.n421 0.155672
R890 source.n483 source.n421 0.155672
R891 source.n376 source.n371 0.155672
R892 source.n383 source.n371 0.155672
R893 source.n384 source.n383 0.155672
R894 source.n384 source.n367 0.155672
R895 source.n391 source.n367 0.155672
R896 source.n392 source.n391 0.155672
R897 source.n392 source.n363 0.155672
R898 source.n401 source.n363 0.155672
R899 source.n402 source.n401 0.155672
R900 source.n402 source.n359 0.155672
R901 source.n409 source.n359 0.155672
R902 source.n410 source.n409 0.155672
R903 source.n410 source.n355 0.155672
R904 source.n417 source.n355 0.155672
R905 source.n302 source.n297 0.155672
R906 source.n309 source.n297 0.155672
R907 source.n310 source.n309 0.155672
R908 source.n310 source.n293 0.155672
R909 source.n317 source.n293 0.155672
R910 source.n318 source.n317 0.155672
R911 source.n318 source.n289 0.155672
R912 source.n327 source.n289 0.155672
R913 source.n328 source.n327 0.155672
R914 source.n328 source.n285 0.155672
R915 source.n335 source.n285 0.155672
R916 source.n336 source.n335 0.155672
R917 source.n336 source.n281 0.155672
R918 source.n343 source.n281 0.155672
R919 source.n63 source.n1 0.155672
R920 source.n56 source.n1 0.155672
R921 source.n56 source.n55 0.155672
R922 source.n55 source.n5 0.155672
R923 source.n48 source.n5 0.155672
R924 source.n48 source.n47 0.155672
R925 source.n47 source.n9 0.155672
R926 source.n39 source.n9 0.155672
R927 source.n39 source.n38 0.155672
R928 source.n38 source.n14 0.155672
R929 source.n31 source.n14 0.155672
R930 source.n31 source.n30 0.155672
R931 source.n30 source.n18 0.155672
R932 source.n23 source.n18 0.155672
R933 source.n137 source.n75 0.155672
R934 source.n130 source.n75 0.155672
R935 source.n130 source.n129 0.155672
R936 source.n129 source.n79 0.155672
R937 source.n122 source.n79 0.155672
R938 source.n122 source.n121 0.155672
R939 source.n121 source.n83 0.155672
R940 source.n113 source.n83 0.155672
R941 source.n113 source.n112 0.155672
R942 source.n112 source.n88 0.155672
R943 source.n105 source.n88 0.155672
R944 source.n105 source.n104 0.155672
R945 source.n104 source.n92 0.155672
R946 source.n97 source.n92 0.155672
R947 source.n203 source.n141 0.155672
R948 source.n196 source.n141 0.155672
R949 source.n196 source.n195 0.155672
R950 source.n195 source.n145 0.155672
R951 source.n188 source.n145 0.155672
R952 source.n188 source.n187 0.155672
R953 source.n187 source.n149 0.155672
R954 source.n179 source.n149 0.155672
R955 source.n179 source.n178 0.155672
R956 source.n178 source.n154 0.155672
R957 source.n171 source.n154 0.155672
R958 source.n171 source.n170 0.155672
R959 source.n170 source.n158 0.155672
R960 source.n163 source.n158 0.155672
R961 source.n277 source.n215 0.155672
R962 source.n270 source.n215 0.155672
R963 source.n270 source.n269 0.155672
R964 source.n269 source.n219 0.155672
R965 source.n262 source.n219 0.155672
R966 source.n262 source.n261 0.155672
R967 source.n261 source.n223 0.155672
R968 source.n253 source.n223 0.155672
R969 source.n253 source.n252 0.155672
R970 source.n252 source.n228 0.155672
R971 source.n245 source.n228 0.155672
R972 source.n245 source.n244 0.155672
R973 source.n244 source.n232 0.155672
R974 source.n237 source.n232 0.155672
R975 drain_right.n6 drain_right.n4 60.5266
R976 drain_right.n2 drain_right.n0 60.5266
R977 drain_right.n10 drain_right.n8 60.5266
R978 drain_right.n10 drain_right.n9 59.5527
R979 drain_right.n12 drain_right.n11 59.5527
R980 drain_right.n14 drain_right.n13 59.5527
R981 drain_right.n16 drain_right.n15 59.5527
R982 drain_right.n7 drain_right.n3 59.5525
R983 drain_right.n6 drain_right.n5 59.5525
R984 drain_right.n2 drain_right.n1 59.5525
R985 drain_right drain_right.n7 34.6069
R986 drain_right drain_right.n16 6.62735
R987 drain_right.n3 drain_right.t1 1.6505
R988 drain_right.n3 drain_right.t17 1.6505
R989 drain_right.n4 drain_right.t4 1.6505
R990 drain_right.n4 drain_right.t18 1.6505
R991 drain_right.n5 drain_right.t5 1.6505
R992 drain_right.n5 drain_right.t19 1.6505
R993 drain_right.n1 drain_right.t3 1.6505
R994 drain_right.n1 drain_right.t16 1.6505
R995 drain_right.n0 drain_right.t0 1.6505
R996 drain_right.n0 drain_right.t14 1.6505
R997 drain_right.n8 drain_right.t12 1.6505
R998 drain_right.n8 drain_right.t10 1.6505
R999 drain_right.n9 drain_right.t8 1.6505
R1000 drain_right.n9 drain_right.t13 1.6505
R1001 drain_right.n11 drain_right.t9 1.6505
R1002 drain_right.n11 drain_right.t6 1.6505
R1003 drain_right.n13 drain_right.t2 1.6505
R1004 drain_right.n13 drain_right.t11 1.6505
R1005 drain_right.n15 drain_right.t15 1.6505
R1006 drain_right.n15 drain_right.t7 1.6505
R1007 drain_right.n16 drain_right.n14 0.974638
R1008 drain_right.n14 drain_right.n12 0.974638
R1009 drain_right.n12 drain_right.n10 0.974638
R1010 drain_right.n7 drain_right.n6 0.919292
R1011 drain_right.n7 drain_right.n2 0.919292
R1012 plus.n9 plus.t18 432.394
R1013 plus.n39 plus.t15 432.394
R1014 plus.n28 plus.t5 410.604
R1015 plus.n26 plus.t6 410.604
R1016 plus.n2 plus.t8 410.604
R1017 plus.n21 plus.t10 410.604
R1018 plus.n19 plus.t11 410.604
R1019 plus.n5 plus.t16 410.604
R1020 plus.n13 plus.t12 410.604
R1021 plus.n12 plus.t13 410.604
R1022 plus.n8 plus.t17 410.604
R1023 plus.n58 plus.t14 410.604
R1024 plus.n56 plus.t3 410.604
R1025 plus.n32 plus.t0 410.604
R1026 plus.n51 plus.t4 410.604
R1027 plus.n49 plus.t19 410.604
R1028 plus.n35 plus.t7 410.604
R1029 plus.n43 plus.t1 410.604
R1030 plus.n42 plus.t9 410.604
R1031 plus.n38 plus.t2 410.604
R1032 plus.n11 plus.n10 161.3
R1033 plus.n15 plus.n14 161.3
R1034 plus.n16 plus.n5 161.3
R1035 plus.n18 plus.n17 161.3
R1036 plus.n19 plus.n4 161.3
R1037 plus.n20 plus.n3 161.3
R1038 plus.n25 plus.n24 161.3
R1039 plus.n26 plus.n1 161.3
R1040 plus.n27 plus.n0 161.3
R1041 plus.n29 plus.n28 161.3
R1042 plus.n41 plus.n40 161.3
R1043 plus.n45 plus.n44 161.3
R1044 plus.n46 plus.n35 161.3
R1045 plus.n48 plus.n47 161.3
R1046 plus.n49 plus.n34 161.3
R1047 plus.n50 plus.n33 161.3
R1048 plus.n55 plus.n54 161.3
R1049 plus.n56 plus.n31 161.3
R1050 plus.n57 plus.n30 161.3
R1051 plus.n59 plus.n58 161.3
R1052 plus.n12 plus.n7 80.6037
R1053 plus.n13 plus.n6 80.6037
R1054 plus.n22 plus.n21 80.6037
R1055 plus.n23 plus.n2 80.6037
R1056 plus.n42 plus.n37 80.6037
R1057 plus.n43 plus.n36 80.6037
R1058 plus.n52 plus.n51 80.6037
R1059 plus.n53 plus.n32 80.6037
R1060 plus.n21 plus.n2 48.2005
R1061 plus.n13 plus.n12 48.2005
R1062 plus.n51 plus.n32 48.2005
R1063 plus.n43 plus.n42 48.2005
R1064 plus.n40 plus.n39 44.8565
R1065 plus.n10 plus.n9 44.8565
R1066 plus.n21 plus.n20 43.0884
R1067 plus.n14 plus.n13 43.0884
R1068 plus.n51 plus.n50 43.0884
R1069 plus.n44 plus.n43 43.0884
R1070 plus.n25 plus.n2 40.1672
R1071 plus.n12 plus.n11 40.1672
R1072 plus.n55 plus.n32 40.1672
R1073 plus.n42 plus.n41 40.1672
R1074 plus plus.n59 35.3361
R1075 plus.n28 plus.n27 27.0217
R1076 plus.n58 plus.n57 27.0217
R1077 plus.n18 plus.n5 24.1005
R1078 plus.n19 plus.n18 24.1005
R1079 plus.n49 plus.n48 24.1005
R1080 plus.n48 plus.n35 24.1005
R1081 plus.n27 plus.n26 21.1793
R1082 plus.n57 plus.n56 21.1793
R1083 plus.n39 plus.n38 20.1275
R1084 plus.n9 plus.n8 20.1275
R1085 plus plus.n29 12.349
R1086 plus.n26 plus.n25 8.03383
R1087 plus.n11 plus.n8 8.03383
R1088 plus.n56 plus.n55 8.03383
R1089 plus.n41 plus.n38 8.03383
R1090 plus.n20 plus.n19 5.11262
R1091 plus.n14 plus.n5 5.11262
R1092 plus.n50 plus.n49 5.11262
R1093 plus.n44 plus.n35 5.11262
R1094 plus.n7 plus.n6 0.380177
R1095 plus.n23 plus.n22 0.380177
R1096 plus.n53 plus.n52 0.380177
R1097 plus.n37 plus.n36 0.380177
R1098 plus.n10 plus.n7 0.285035
R1099 plus.n15 plus.n6 0.285035
R1100 plus.n22 plus.n3 0.285035
R1101 plus.n24 plus.n23 0.285035
R1102 plus.n54 plus.n53 0.285035
R1103 plus.n52 plus.n33 0.285035
R1104 plus.n45 plus.n36 0.285035
R1105 plus.n40 plus.n37 0.285035
R1106 plus.n16 plus.n15 0.189894
R1107 plus.n17 plus.n16 0.189894
R1108 plus.n17 plus.n4 0.189894
R1109 plus.n4 plus.n3 0.189894
R1110 plus.n24 plus.n1 0.189894
R1111 plus.n1 plus.n0 0.189894
R1112 plus.n29 plus.n0 0.189894
R1113 plus.n59 plus.n30 0.189894
R1114 plus.n31 plus.n30 0.189894
R1115 plus.n54 plus.n31 0.189894
R1116 plus.n34 plus.n33 0.189894
R1117 plus.n47 plus.n34 0.189894
R1118 plus.n47 plus.n46 0.189894
R1119 plus.n46 plus.n45 0.189894
R1120 drain_left.n10 drain_left.n8 60.5268
R1121 drain_left.n6 drain_left.n4 60.5266
R1122 drain_left.n2 drain_left.n0 60.5266
R1123 drain_left.n14 drain_left.n13 59.5527
R1124 drain_left.n12 drain_left.n11 59.5527
R1125 drain_left.n10 drain_left.n9 59.5527
R1126 drain_left.n7 drain_left.n3 59.5525
R1127 drain_left.n6 drain_left.n5 59.5525
R1128 drain_left.n2 drain_left.n1 59.5525
R1129 drain_left.n16 drain_left.n15 59.5525
R1130 drain_left drain_left.n7 35.1602
R1131 drain_left drain_left.n16 6.62735
R1132 drain_left.n3 drain_left.t0 1.6505
R1133 drain_left.n3 drain_left.t12 1.6505
R1134 drain_left.n4 drain_left.t17 1.6505
R1135 drain_left.n4 drain_left.t4 1.6505
R1136 drain_left.n5 drain_left.t18 1.6505
R1137 drain_left.n5 drain_left.t10 1.6505
R1138 drain_left.n1 drain_left.t19 1.6505
R1139 drain_left.n1 drain_left.t15 1.6505
R1140 drain_left.n0 drain_left.t5 1.6505
R1141 drain_left.n0 drain_left.t16 1.6505
R1142 drain_left.n15 drain_left.t13 1.6505
R1143 drain_left.n15 drain_left.t14 1.6505
R1144 drain_left.n13 drain_left.t9 1.6505
R1145 drain_left.n13 drain_left.t11 1.6505
R1146 drain_left.n11 drain_left.t3 1.6505
R1147 drain_left.n11 drain_left.t8 1.6505
R1148 drain_left.n9 drain_left.t6 1.6505
R1149 drain_left.n9 drain_left.t7 1.6505
R1150 drain_left.n8 drain_left.t1 1.6505
R1151 drain_left.n8 drain_left.t2 1.6505
R1152 drain_left.n12 drain_left.n10 0.974638
R1153 drain_left.n14 drain_left.n12 0.974638
R1154 drain_left.n16 drain_left.n14 0.974638
R1155 drain_left.n7 drain_left.n6 0.919292
R1156 drain_left.n7 drain_left.n2 0.919292
C0 drain_right drain_left 1.72917f
C1 minus source 13.7795f
C2 plus source 13.793599f
C3 minus drain_left 0.17405f
C4 minus drain_right 13.5374f
C5 plus drain_left 13.8578f
C6 plus drain_right 0.478206f
C7 plus minus 7.1383f
C8 source drain_left 22.4917f
C9 source drain_right 22.4945f
C10 drain_right a_n3202_n3288# 7.51032f
C11 drain_left a_n3202_n3288# 7.96142f
C12 source a_n3202_n3288# 9.567579f
C13 minus a_n3202_n3288# 12.935336f
C14 plus a_n3202_n3288# 14.70884f
C15 drain_left.t5 a_n3202_n3288# 0.253f
C16 drain_left.t16 a_n3202_n3288# 0.253f
C17 drain_left.n0 a_n3202_n3288# 2.25778f
C18 drain_left.t19 a_n3202_n3288# 0.253f
C19 drain_left.t15 a_n3202_n3288# 0.253f
C20 drain_left.n1 a_n3202_n3288# 2.25131f
C21 drain_left.n2 a_n3202_n3288# 0.782998f
C22 drain_left.t0 a_n3202_n3288# 0.253f
C23 drain_left.t12 a_n3202_n3288# 0.253f
C24 drain_left.n3 a_n3202_n3288# 2.25131f
C25 drain_left.t17 a_n3202_n3288# 0.253f
C26 drain_left.t4 a_n3202_n3288# 0.253f
C27 drain_left.n4 a_n3202_n3288# 2.25778f
C28 drain_left.t18 a_n3202_n3288# 0.253f
C29 drain_left.t10 a_n3202_n3288# 0.253f
C30 drain_left.n5 a_n3202_n3288# 2.25131f
C31 drain_left.n6 a_n3202_n3288# 0.782998f
C32 drain_left.n7 a_n3202_n3288# 2.02246f
C33 drain_left.t1 a_n3202_n3288# 0.253f
C34 drain_left.t2 a_n3202_n3288# 0.253f
C35 drain_left.n8 a_n3202_n3288# 2.25779f
C36 drain_left.t6 a_n3202_n3288# 0.253f
C37 drain_left.t7 a_n3202_n3288# 0.253f
C38 drain_left.n9 a_n3202_n3288# 2.25132f
C39 drain_left.n10 a_n3202_n3288# 0.787064f
C40 drain_left.t3 a_n3202_n3288# 0.253f
C41 drain_left.t8 a_n3202_n3288# 0.253f
C42 drain_left.n11 a_n3202_n3288# 2.25132f
C43 drain_left.n12 a_n3202_n3288# 0.391395f
C44 drain_left.t9 a_n3202_n3288# 0.253f
C45 drain_left.t11 a_n3202_n3288# 0.253f
C46 drain_left.n13 a_n3202_n3288# 2.25132f
C47 drain_left.n14 a_n3202_n3288# 0.391395f
C48 drain_left.t13 a_n3202_n3288# 0.253f
C49 drain_left.t14 a_n3202_n3288# 0.253f
C50 drain_left.n15 a_n3202_n3288# 2.25131f
C51 drain_left.n16 a_n3202_n3288# 0.630642f
C52 plus.n0 a_n3202_n3288# 0.038191f
C53 plus.t5 a_n3202_n3288# 1.04547f
C54 plus.t6 a_n3202_n3288# 1.04547f
C55 plus.n1 a_n3202_n3288# 0.038191f
C56 plus.t8 a_n3202_n3288# 1.04547f
C57 plus.n2 a_n3202_n3288# 0.423893f
C58 plus.n3 a_n3202_n3288# 0.050961f
C59 plus.t10 a_n3202_n3288# 1.04547f
C60 plus.t11 a_n3202_n3288# 1.04547f
C61 plus.n4 a_n3202_n3288# 0.038191f
C62 plus.t16 a_n3202_n3288# 1.04547f
C63 plus.n5 a_n3202_n3288# 0.413461f
C64 plus.n6 a_n3202_n3288# 0.063612f
C65 plus.t12 a_n3202_n3288# 1.04547f
C66 plus.t13 a_n3202_n3288# 1.04547f
C67 plus.n7 a_n3202_n3288# 0.063612f
C68 plus.t17 a_n3202_n3288# 1.04547f
C69 plus.n8 a_n3202_n3288# 0.416671f
C70 plus.t18 a_n3202_n3288# 1.06641f
C71 plus.n9 a_n3202_n3288# 0.398429f
C72 plus.n10 a_n3202_n3288# 0.175793f
C73 plus.n11 a_n3202_n3288# 0.008666f
C74 plus.n12 a_n3202_n3288# 0.423893f
C75 plus.n13 a_n3202_n3288# 0.424364f
C76 plus.n14 a_n3202_n3288# 0.008666f
C77 plus.n15 a_n3202_n3288# 0.050961f
C78 plus.n16 a_n3202_n3288# 0.038191f
C79 plus.n17 a_n3202_n3288# 0.038191f
C80 plus.n18 a_n3202_n3288# 0.008666f
C81 plus.n19 a_n3202_n3288# 0.413461f
C82 plus.n20 a_n3202_n3288# 0.008666f
C83 plus.n21 a_n3202_n3288# 0.424364f
C84 plus.n22 a_n3202_n3288# 0.063612f
C85 plus.n23 a_n3202_n3288# 0.063612f
C86 plus.n24 a_n3202_n3288# 0.050961f
C87 plus.n25 a_n3202_n3288# 0.008666f
C88 plus.n26 a_n3202_n3288# 0.413461f
C89 plus.n27 a_n3202_n3288# 0.008666f
C90 plus.n28 a_n3202_n3288# 0.413107f
C91 plus.n29 a_n3202_n3288# 0.445927f
C92 plus.n30 a_n3202_n3288# 0.038191f
C93 plus.t14 a_n3202_n3288# 1.04547f
C94 plus.n31 a_n3202_n3288# 0.038191f
C95 plus.t3 a_n3202_n3288# 1.04547f
C96 plus.t0 a_n3202_n3288# 1.04547f
C97 plus.n32 a_n3202_n3288# 0.423893f
C98 plus.n33 a_n3202_n3288# 0.050961f
C99 plus.t4 a_n3202_n3288# 1.04547f
C100 plus.n34 a_n3202_n3288# 0.038191f
C101 plus.t19 a_n3202_n3288# 1.04547f
C102 plus.t7 a_n3202_n3288# 1.04547f
C103 plus.n35 a_n3202_n3288# 0.413461f
C104 plus.n36 a_n3202_n3288# 0.063612f
C105 plus.t1 a_n3202_n3288# 1.04547f
C106 plus.n37 a_n3202_n3288# 0.063612f
C107 plus.t9 a_n3202_n3288# 1.04547f
C108 plus.t2 a_n3202_n3288# 1.04547f
C109 plus.n38 a_n3202_n3288# 0.416671f
C110 plus.t15 a_n3202_n3288# 1.06641f
C111 plus.n39 a_n3202_n3288# 0.398429f
C112 plus.n40 a_n3202_n3288# 0.175793f
C113 plus.n41 a_n3202_n3288# 0.008666f
C114 plus.n42 a_n3202_n3288# 0.423893f
C115 plus.n43 a_n3202_n3288# 0.424364f
C116 plus.n44 a_n3202_n3288# 0.008666f
C117 plus.n45 a_n3202_n3288# 0.050961f
C118 plus.n46 a_n3202_n3288# 0.038191f
C119 plus.n47 a_n3202_n3288# 0.038191f
C120 plus.n48 a_n3202_n3288# 0.008666f
C121 plus.n49 a_n3202_n3288# 0.413461f
C122 plus.n50 a_n3202_n3288# 0.008666f
C123 plus.n51 a_n3202_n3288# 0.424364f
C124 plus.n52 a_n3202_n3288# 0.063612f
C125 plus.n53 a_n3202_n3288# 0.063612f
C126 plus.n54 a_n3202_n3288# 0.050961f
C127 plus.n55 a_n3202_n3288# 0.008666f
C128 plus.n56 a_n3202_n3288# 0.413461f
C129 plus.n57 a_n3202_n3288# 0.008666f
C130 plus.n58 a_n3202_n3288# 0.413107f
C131 plus.n59 a_n3202_n3288# 1.42832f
C132 drain_right.t0 a_n3202_n3288# 0.250939f
C133 drain_right.t14 a_n3202_n3288# 0.250939f
C134 drain_right.n0 a_n3202_n3288# 2.23939f
C135 drain_right.t3 a_n3202_n3288# 0.250939f
C136 drain_right.t16 a_n3202_n3288# 0.250939f
C137 drain_right.n1 a_n3202_n3288# 2.23297f
C138 drain_right.n2 a_n3202_n3288# 0.77662f
C139 drain_right.t1 a_n3202_n3288# 0.250939f
C140 drain_right.t17 a_n3202_n3288# 0.250939f
C141 drain_right.n3 a_n3202_n3288# 2.23297f
C142 drain_right.t4 a_n3202_n3288# 0.250939f
C143 drain_right.t18 a_n3202_n3288# 0.250939f
C144 drain_right.n4 a_n3202_n3288# 2.23939f
C145 drain_right.t5 a_n3202_n3288# 0.250939f
C146 drain_right.t19 a_n3202_n3288# 0.250939f
C147 drain_right.n5 a_n3202_n3288# 2.23297f
C148 drain_right.n6 a_n3202_n3288# 0.77662f
C149 drain_right.n7 a_n3202_n3288# 1.95226f
C150 drain_right.t12 a_n3202_n3288# 0.250939f
C151 drain_right.t10 a_n3202_n3288# 0.250939f
C152 drain_right.n8 a_n3202_n3288# 2.23939f
C153 drain_right.t8 a_n3202_n3288# 0.250939f
C154 drain_right.t13 a_n3202_n3288# 0.250939f
C155 drain_right.n9 a_n3202_n3288# 2.23298f
C156 drain_right.n10 a_n3202_n3288# 0.780662f
C157 drain_right.t9 a_n3202_n3288# 0.250939f
C158 drain_right.t6 a_n3202_n3288# 0.250939f
C159 drain_right.n11 a_n3202_n3288# 2.23298f
C160 drain_right.n12 a_n3202_n3288# 0.388207f
C161 drain_right.t2 a_n3202_n3288# 0.250939f
C162 drain_right.t11 a_n3202_n3288# 0.250939f
C163 drain_right.n13 a_n3202_n3288# 2.23298f
C164 drain_right.n14 a_n3202_n3288# 0.388207f
C165 drain_right.t15 a_n3202_n3288# 0.250939f
C166 drain_right.t7 a_n3202_n3288# 0.250939f
C167 drain_right.n15 a_n3202_n3288# 2.23298f
C168 drain_right.n16 a_n3202_n3288# 0.625496f
C169 source.n0 a_n3202_n3288# 0.031451f
C170 source.n1 a_n3202_n3288# 0.023743f
C171 source.n2 a_n3202_n3288# 0.012759f
C172 source.n3 a_n3202_n3288# 0.030157f
C173 source.n4 a_n3202_n3288# 0.013509f
C174 source.n5 a_n3202_n3288# 0.023743f
C175 source.n6 a_n3202_n3288# 0.012759f
C176 source.n7 a_n3202_n3288# 0.030157f
C177 source.n8 a_n3202_n3288# 0.013509f
C178 source.n9 a_n3202_n3288# 0.023743f
C179 source.n10 a_n3202_n3288# 0.013134f
C180 source.n11 a_n3202_n3288# 0.030157f
C181 source.n12 a_n3202_n3288# 0.012759f
C182 source.n13 a_n3202_n3288# 0.013509f
C183 source.n14 a_n3202_n3288# 0.023743f
C184 source.n15 a_n3202_n3288# 0.012759f
C185 source.n16 a_n3202_n3288# 0.030157f
C186 source.n17 a_n3202_n3288# 0.013509f
C187 source.n18 a_n3202_n3288# 0.023743f
C188 source.n19 a_n3202_n3288# 0.012759f
C189 source.n20 a_n3202_n3288# 0.022618f
C190 source.n21 a_n3202_n3288# 0.021319f
C191 source.t17 a_n3202_n3288# 0.050933f
C192 source.n22 a_n3202_n3288# 0.171186f
C193 source.n23 a_n3202_n3288# 1.19781f
C194 source.n24 a_n3202_n3288# 0.012759f
C195 source.n25 a_n3202_n3288# 0.013509f
C196 source.n26 a_n3202_n3288# 0.030157f
C197 source.n27 a_n3202_n3288# 0.030157f
C198 source.n28 a_n3202_n3288# 0.013509f
C199 source.n29 a_n3202_n3288# 0.012759f
C200 source.n30 a_n3202_n3288# 0.023743f
C201 source.n31 a_n3202_n3288# 0.023743f
C202 source.n32 a_n3202_n3288# 0.012759f
C203 source.n33 a_n3202_n3288# 0.013509f
C204 source.n34 a_n3202_n3288# 0.030157f
C205 source.n35 a_n3202_n3288# 0.030157f
C206 source.n36 a_n3202_n3288# 0.013509f
C207 source.n37 a_n3202_n3288# 0.012759f
C208 source.n38 a_n3202_n3288# 0.023743f
C209 source.n39 a_n3202_n3288# 0.023743f
C210 source.n40 a_n3202_n3288# 0.012759f
C211 source.n41 a_n3202_n3288# 0.013509f
C212 source.n42 a_n3202_n3288# 0.030157f
C213 source.n43 a_n3202_n3288# 0.030157f
C214 source.n44 a_n3202_n3288# 0.030157f
C215 source.n45 a_n3202_n3288# 0.013134f
C216 source.n46 a_n3202_n3288# 0.012759f
C217 source.n47 a_n3202_n3288# 0.023743f
C218 source.n48 a_n3202_n3288# 0.023743f
C219 source.n49 a_n3202_n3288# 0.012759f
C220 source.n50 a_n3202_n3288# 0.013509f
C221 source.n51 a_n3202_n3288# 0.030157f
C222 source.n52 a_n3202_n3288# 0.030157f
C223 source.n53 a_n3202_n3288# 0.013509f
C224 source.n54 a_n3202_n3288# 0.012759f
C225 source.n55 a_n3202_n3288# 0.023743f
C226 source.n56 a_n3202_n3288# 0.023743f
C227 source.n57 a_n3202_n3288# 0.012759f
C228 source.n58 a_n3202_n3288# 0.013509f
C229 source.n59 a_n3202_n3288# 0.030157f
C230 source.n60 a_n3202_n3288# 0.061885f
C231 source.n61 a_n3202_n3288# 0.013509f
C232 source.n62 a_n3202_n3288# 0.012759f
C233 source.n63 a_n3202_n3288# 0.050989f
C234 source.n64 a_n3202_n3288# 0.034154f
C235 source.n65 a_n3202_n3288# 1.00959f
C236 source.t11 a_n3202_n3288# 0.225152f
C237 source.t8 a_n3202_n3288# 0.225152f
C238 source.n66 a_n3202_n3288# 1.92776f
C239 source.n67 a_n3202_n3288# 0.3918f
C240 source.t14 a_n3202_n3288# 0.225152f
C241 source.t10 a_n3202_n3288# 0.225152f
C242 source.n68 a_n3202_n3288# 1.92776f
C243 source.n69 a_n3202_n3288# 0.3918f
C244 source.t3 a_n3202_n3288# 0.225152f
C245 source.t4 a_n3202_n3288# 0.225152f
C246 source.n70 a_n3202_n3288# 1.92776f
C247 source.n71 a_n3202_n3288# 0.3918f
C248 source.t2 a_n3202_n3288# 0.225152f
C249 source.t16 a_n3202_n3288# 0.225152f
C250 source.n72 a_n3202_n3288# 1.92776f
C251 source.n73 a_n3202_n3288# 0.3918f
C252 source.n74 a_n3202_n3288# 0.031451f
C253 source.n75 a_n3202_n3288# 0.023743f
C254 source.n76 a_n3202_n3288# 0.012759f
C255 source.n77 a_n3202_n3288# 0.030157f
C256 source.n78 a_n3202_n3288# 0.013509f
C257 source.n79 a_n3202_n3288# 0.023743f
C258 source.n80 a_n3202_n3288# 0.012759f
C259 source.n81 a_n3202_n3288# 0.030157f
C260 source.n82 a_n3202_n3288# 0.013509f
C261 source.n83 a_n3202_n3288# 0.023743f
C262 source.n84 a_n3202_n3288# 0.013134f
C263 source.n85 a_n3202_n3288# 0.030157f
C264 source.n86 a_n3202_n3288# 0.012759f
C265 source.n87 a_n3202_n3288# 0.013509f
C266 source.n88 a_n3202_n3288# 0.023743f
C267 source.n89 a_n3202_n3288# 0.012759f
C268 source.n90 a_n3202_n3288# 0.030157f
C269 source.n91 a_n3202_n3288# 0.013509f
C270 source.n92 a_n3202_n3288# 0.023743f
C271 source.n93 a_n3202_n3288# 0.012759f
C272 source.n94 a_n3202_n3288# 0.022618f
C273 source.n95 a_n3202_n3288# 0.021319f
C274 source.t12 a_n3202_n3288# 0.050933f
C275 source.n96 a_n3202_n3288# 0.171186f
C276 source.n97 a_n3202_n3288# 1.19781f
C277 source.n98 a_n3202_n3288# 0.012759f
C278 source.n99 a_n3202_n3288# 0.013509f
C279 source.n100 a_n3202_n3288# 0.030157f
C280 source.n101 a_n3202_n3288# 0.030157f
C281 source.n102 a_n3202_n3288# 0.013509f
C282 source.n103 a_n3202_n3288# 0.012759f
C283 source.n104 a_n3202_n3288# 0.023743f
C284 source.n105 a_n3202_n3288# 0.023743f
C285 source.n106 a_n3202_n3288# 0.012759f
C286 source.n107 a_n3202_n3288# 0.013509f
C287 source.n108 a_n3202_n3288# 0.030157f
C288 source.n109 a_n3202_n3288# 0.030157f
C289 source.n110 a_n3202_n3288# 0.013509f
C290 source.n111 a_n3202_n3288# 0.012759f
C291 source.n112 a_n3202_n3288# 0.023743f
C292 source.n113 a_n3202_n3288# 0.023743f
C293 source.n114 a_n3202_n3288# 0.012759f
C294 source.n115 a_n3202_n3288# 0.013509f
C295 source.n116 a_n3202_n3288# 0.030157f
C296 source.n117 a_n3202_n3288# 0.030157f
C297 source.n118 a_n3202_n3288# 0.030157f
C298 source.n119 a_n3202_n3288# 0.013134f
C299 source.n120 a_n3202_n3288# 0.012759f
C300 source.n121 a_n3202_n3288# 0.023743f
C301 source.n122 a_n3202_n3288# 0.023743f
C302 source.n123 a_n3202_n3288# 0.012759f
C303 source.n124 a_n3202_n3288# 0.013509f
C304 source.n125 a_n3202_n3288# 0.030157f
C305 source.n126 a_n3202_n3288# 0.030157f
C306 source.n127 a_n3202_n3288# 0.013509f
C307 source.n128 a_n3202_n3288# 0.012759f
C308 source.n129 a_n3202_n3288# 0.023743f
C309 source.n130 a_n3202_n3288# 0.023743f
C310 source.n131 a_n3202_n3288# 0.012759f
C311 source.n132 a_n3202_n3288# 0.013509f
C312 source.n133 a_n3202_n3288# 0.030157f
C313 source.n134 a_n3202_n3288# 0.061885f
C314 source.n135 a_n3202_n3288# 0.013509f
C315 source.n136 a_n3202_n3288# 0.012759f
C316 source.n137 a_n3202_n3288# 0.050989f
C317 source.n138 a_n3202_n3288# 0.034154f
C318 source.n139 a_n3202_n3288# 0.128558f
C319 source.n140 a_n3202_n3288# 0.031451f
C320 source.n141 a_n3202_n3288# 0.023743f
C321 source.n142 a_n3202_n3288# 0.012759f
C322 source.n143 a_n3202_n3288# 0.030157f
C323 source.n144 a_n3202_n3288# 0.013509f
C324 source.n145 a_n3202_n3288# 0.023743f
C325 source.n146 a_n3202_n3288# 0.012759f
C326 source.n147 a_n3202_n3288# 0.030157f
C327 source.n148 a_n3202_n3288# 0.013509f
C328 source.n149 a_n3202_n3288# 0.023743f
C329 source.n150 a_n3202_n3288# 0.013134f
C330 source.n151 a_n3202_n3288# 0.030157f
C331 source.n152 a_n3202_n3288# 0.012759f
C332 source.n153 a_n3202_n3288# 0.013509f
C333 source.n154 a_n3202_n3288# 0.023743f
C334 source.n155 a_n3202_n3288# 0.012759f
C335 source.n156 a_n3202_n3288# 0.030157f
C336 source.n157 a_n3202_n3288# 0.013509f
C337 source.n158 a_n3202_n3288# 0.023743f
C338 source.n159 a_n3202_n3288# 0.012759f
C339 source.n160 a_n3202_n3288# 0.022618f
C340 source.n161 a_n3202_n3288# 0.021319f
C341 source.t30 a_n3202_n3288# 0.050933f
C342 source.n162 a_n3202_n3288# 0.171186f
C343 source.n163 a_n3202_n3288# 1.19781f
C344 source.n164 a_n3202_n3288# 0.012759f
C345 source.n165 a_n3202_n3288# 0.013509f
C346 source.n166 a_n3202_n3288# 0.030157f
C347 source.n167 a_n3202_n3288# 0.030157f
C348 source.n168 a_n3202_n3288# 0.013509f
C349 source.n169 a_n3202_n3288# 0.012759f
C350 source.n170 a_n3202_n3288# 0.023743f
C351 source.n171 a_n3202_n3288# 0.023743f
C352 source.n172 a_n3202_n3288# 0.012759f
C353 source.n173 a_n3202_n3288# 0.013509f
C354 source.n174 a_n3202_n3288# 0.030157f
C355 source.n175 a_n3202_n3288# 0.030157f
C356 source.n176 a_n3202_n3288# 0.013509f
C357 source.n177 a_n3202_n3288# 0.012759f
C358 source.n178 a_n3202_n3288# 0.023743f
C359 source.n179 a_n3202_n3288# 0.023743f
C360 source.n180 a_n3202_n3288# 0.012759f
C361 source.n181 a_n3202_n3288# 0.013509f
C362 source.n182 a_n3202_n3288# 0.030157f
C363 source.n183 a_n3202_n3288# 0.030157f
C364 source.n184 a_n3202_n3288# 0.030157f
C365 source.n185 a_n3202_n3288# 0.013134f
C366 source.n186 a_n3202_n3288# 0.012759f
C367 source.n187 a_n3202_n3288# 0.023743f
C368 source.n188 a_n3202_n3288# 0.023743f
C369 source.n189 a_n3202_n3288# 0.012759f
C370 source.n190 a_n3202_n3288# 0.013509f
C371 source.n191 a_n3202_n3288# 0.030157f
C372 source.n192 a_n3202_n3288# 0.030157f
C373 source.n193 a_n3202_n3288# 0.013509f
C374 source.n194 a_n3202_n3288# 0.012759f
C375 source.n195 a_n3202_n3288# 0.023743f
C376 source.n196 a_n3202_n3288# 0.023743f
C377 source.n197 a_n3202_n3288# 0.012759f
C378 source.n198 a_n3202_n3288# 0.013509f
C379 source.n199 a_n3202_n3288# 0.030157f
C380 source.n200 a_n3202_n3288# 0.061885f
C381 source.n201 a_n3202_n3288# 0.013509f
C382 source.n202 a_n3202_n3288# 0.012759f
C383 source.n203 a_n3202_n3288# 0.050989f
C384 source.n204 a_n3202_n3288# 0.034154f
C385 source.n205 a_n3202_n3288# 0.128558f
C386 source.t26 a_n3202_n3288# 0.225152f
C387 source.t19 a_n3202_n3288# 0.225152f
C388 source.n206 a_n3202_n3288# 1.92776f
C389 source.n207 a_n3202_n3288# 0.3918f
C390 source.t27 a_n3202_n3288# 0.225152f
C391 source.t35 a_n3202_n3288# 0.225152f
C392 source.n208 a_n3202_n3288# 1.92776f
C393 source.n209 a_n3202_n3288# 0.3918f
C394 source.t32 a_n3202_n3288# 0.225152f
C395 source.t36 a_n3202_n3288# 0.225152f
C396 source.n210 a_n3202_n3288# 1.92776f
C397 source.n211 a_n3202_n3288# 0.3918f
C398 source.t24 a_n3202_n3288# 0.225152f
C399 source.t31 a_n3202_n3288# 0.225152f
C400 source.n212 a_n3202_n3288# 1.92776f
C401 source.n213 a_n3202_n3288# 0.3918f
C402 source.n214 a_n3202_n3288# 0.031451f
C403 source.n215 a_n3202_n3288# 0.023743f
C404 source.n216 a_n3202_n3288# 0.012759f
C405 source.n217 a_n3202_n3288# 0.030157f
C406 source.n218 a_n3202_n3288# 0.013509f
C407 source.n219 a_n3202_n3288# 0.023743f
C408 source.n220 a_n3202_n3288# 0.012759f
C409 source.n221 a_n3202_n3288# 0.030157f
C410 source.n222 a_n3202_n3288# 0.013509f
C411 source.n223 a_n3202_n3288# 0.023743f
C412 source.n224 a_n3202_n3288# 0.013134f
C413 source.n225 a_n3202_n3288# 0.030157f
C414 source.n226 a_n3202_n3288# 0.012759f
C415 source.n227 a_n3202_n3288# 0.013509f
C416 source.n228 a_n3202_n3288# 0.023743f
C417 source.n229 a_n3202_n3288# 0.012759f
C418 source.n230 a_n3202_n3288# 0.030157f
C419 source.n231 a_n3202_n3288# 0.013509f
C420 source.n232 a_n3202_n3288# 0.023743f
C421 source.n233 a_n3202_n3288# 0.012759f
C422 source.n234 a_n3202_n3288# 0.022618f
C423 source.n235 a_n3202_n3288# 0.021319f
C424 source.t34 a_n3202_n3288# 0.050933f
C425 source.n236 a_n3202_n3288# 0.171186f
C426 source.n237 a_n3202_n3288# 1.19781f
C427 source.n238 a_n3202_n3288# 0.012759f
C428 source.n239 a_n3202_n3288# 0.013509f
C429 source.n240 a_n3202_n3288# 0.030157f
C430 source.n241 a_n3202_n3288# 0.030157f
C431 source.n242 a_n3202_n3288# 0.013509f
C432 source.n243 a_n3202_n3288# 0.012759f
C433 source.n244 a_n3202_n3288# 0.023743f
C434 source.n245 a_n3202_n3288# 0.023743f
C435 source.n246 a_n3202_n3288# 0.012759f
C436 source.n247 a_n3202_n3288# 0.013509f
C437 source.n248 a_n3202_n3288# 0.030157f
C438 source.n249 a_n3202_n3288# 0.030157f
C439 source.n250 a_n3202_n3288# 0.013509f
C440 source.n251 a_n3202_n3288# 0.012759f
C441 source.n252 a_n3202_n3288# 0.023743f
C442 source.n253 a_n3202_n3288# 0.023743f
C443 source.n254 a_n3202_n3288# 0.012759f
C444 source.n255 a_n3202_n3288# 0.013509f
C445 source.n256 a_n3202_n3288# 0.030157f
C446 source.n257 a_n3202_n3288# 0.030157f
C447 source.n258 a_n3202_n3288# 0.030157f
C448 source.n259 a_n3202_n3288# 0.013134f
C449 source.n260 a_n3202_n3288# 0.012759f
C450 source.n261 a_n3202_n3288# 0.023743f
C451 source.n262 a_n3202_n3288# 0.023743f
C452 source.n263 a_n3202_n3288# 0.012759f
C453 source.n264 a_n3202_n3288# 0.013509f
C454 source.n265 a_n3202_n3288# 0.030157f
C455 source.n266 a_n3202_n3288# 0.030157f
C456 source.n267 a_n3202_n3288# 0.013509f
C457 source.n268 a_n3202_n3288# 0.012759f
C458 source.n269 a_n3202_n3288# 0.023743f
C459 source.n270 a_n3202_n3288# 0.023743f
C460 source.n271 a_n3202_n3288# 0.012759f
C461 source.n272 a_n3202_n3288# 0.013509f
C462 source.n273 a_n3202_n3288# 0.030157f
C463 source.n274 a_n3202_n3288# 0.061885f
C464 source.n275 a_n3202_n3288# 0.013509f
C465 source.n276 a_n3202_n3288# 0.012759f
C466 source.n277 a_n3202_n3288# 0.050989f
C467 source.n278 a_n3202_n3288# 0.034154f
C468 source.n279 a_n3202_n3288# 1.39485f
C469 source.n280 a_n3202_n3288# 0.031451f
C470 source.n281 a_n3202_n3288# 0.023743f
C471 source.n282 a_n3202_n3288# 0.012759f
C472 source.n283 a_n3202_n3288# 0.030157f
C473 source.n284 a_n3202_n3288# 0.013509f
C474 source.n285 a_n3202_n3288# 0.023743f
C475 source.n286 a_n3202_n3288# 0.012759f
C476 source.n287 a_n3202_n3288# 0.030157f
C477 source.n288 a_n3202_n3288# 0.013509f
C478 source.n289 a_n3202_n3288# 0.023743f
C479 source.n290 a_n3202_n3288# 0.013134f
C480 source.n291 a_n3202_n3288# 0.030157f
C481 source.n292 a_n3202_n3288# 0.013509f
C482 source.n293 a_n3202_n3288# 0.023743f
C483 source.n294 a_n3202_n3288# 0.012759f
C484 source.n295 a_n3202_n3288# 0.030157f
C485 source.n296 a_n3202_n3288# 0.013509f
C486 source.n297 a_n3202_n3288# 0.023743f
C487 source.n298 a_n3202_n3288# 0.012759f
C488 source.n299 a_n3202_n3288# 0.022618f
C489 source.n300 a_n3202_n3288# 0.021319f
C490 source.t13 a_n3202_n3288# 0.050933f
C491 source.n301 a_n3202_n3288# 0.171186f
C492 source.n302 a_n3202_n3288# 1.19781f
C493 source.n303 a_n3202_n3288# 0.012759f
C494 source.n304 a_n3202_n3288# 0.013509f
C495 source.n305 a_n3202_n3288# 0.030157f
C496 source.n306 a_n3202_n3288# 0.030157f
C497 source.n307 a_n3202_n3288# 0.013509f
C498 source.n308 a_n3202_n3288# 0.012759f
C499 source.n309 a_n3202_n3288# 0.023743f
C500 source.n310 a_n3202_n3288# 0.023743f
C501 source.n311 a_n3202_n3288# 0.012759f
C502 source.n312 a_n3202_n3288# 0.013509f
C503 source.n313 a_n3202_n3288# 0.030157f
C504 source.n314 a_n3202_n3288# 0.030157f
C505 source.n315 a_n3202_n3288# 0.013509f
C506 source.n316 a_n3202_n3288# 0.012759f
C507 source.n317 a_n3202_n3288# 0.023743f
C508 source.n318 a_n3202_n3288# 0.023743f
C509 source.n319 a_n3202_n3288# 0.012759f
C510 source.n320 a_n3202_n3288# 0.012759f
C511 source.n321 a_n3202_n3288# 0.013509f
C512 source.n322 a_n3202_n3288# 0.030157f
C513 source.n323 a_n3202_n3288# 0.030157f
C514 source.n324 a_n3202_n3288# 0.030157f
C515 source.n325 a_n3202_n3288# 0.013134f
C516 source.n326 a_n3202_n3288# 0.012759f
C517 source.n327 a_n3202_n3288# 0.023743f
C518 source.n328 a_n3202_n3288# 0.023743f
C519 source.n329 a_n3202_n3288# 0.012759f
C520 source.n330 a_n3202_n3288# 0.013509f
C521 source.n331 a_n3202_n3288# 0.030157f
C522 source.n332 a_n3202_n3288# 0.030157f
C523 source.n333 a_n3202_n3288# 0.013509f
C524 source.n334 a_n3202_n3288# 0.012759f
C525 source.n335 a_n3202_n3288# 0.023743f
C526 source.n336 a_n3202_n3288# 0.023743f
C527 source.n337 a_n3202_n3288# 0.012759f
C528 source.n338 a_n3202_n3288# 0.013509f
C529 source.n339 a_n3202_n3288# 0.030157f
C530 source.n340 a_n3202_n3288# 0.061885f
C531 source.n341 a_n3202_n3288# 0.013509f
C532 source.n342 a_n3202_n3288# 0.012759f
C533 source.n343 a_n3202_n3288# 0.050989f
C534 source.n344 a_n3202_n3288# 0.034154f
C535 source.n345 a_n3202_n3288# 1.39485f
C536 source.t7 a_n3202_n3288# 0.225152f
C537 source.t9 a_n3202_n3288# 0.225152f
C538 source.n346 a_n3202_n3288# 1.92775f
C539 source.n347 a_n3202_n3288# 0.391812f
C540 source.t1 a_n3202_n3288# 0.225152f
C541 source.t5 a_n3202_n3288# 0.225152f
C542 source.n348 a_n3202_n3288# 1.92775f
C543 source.n349 a_n3202_n3288# 0.391812f
C544 source.t0 a_n3202_n3288# 0.225152f
C545 source.t6 a_n3202_n3288# 0.225152f
C546 source.n350 a_n3202_n3288# 1.92775f
C547 source.n351 a_n3202_n3288# 0.391812f
C548 source.t18 a_n3202_n3288# 0.225152f
C549 source.t15 a_n3202_n3288# 0.225152f
C550 source.n352 a_n3202_n3288# 1.92775f
C551 source.n353 a_n3202_n3288# 0.391812f
C552 source.n354 a_n3202_n3288# 0.031451f
C553 source.n355 a_n3202_n3288# 0.023743f
C554 source.n356 a_n3202_n3288# 0.012759f
C555 source.n357 a_n3202_n3288# 0.030157f
C556 source.n358 a_n3202_n3288# 0.013509f
C557 source.n359 a_n3202_n3288# 0.023743f
C558 source.n360 a_n3202_n3288# 0.012759f
C559 source.n361 a_n3202_n3288# 0.030157f
C560 source.n362 a_n3202_n3288# 0.013509f
C561 source.n363 a_n3202_n3288# 0.023743f
C562 source.n364 a_n3202_n3288# 0.013134f
C563 source.n365 a_n3202_n3288# 0.030157f
C564 source.n366 a_n3202_n3288# 0.013509f
C565 source.n367 a_n3202_n3288# 0.023743f
C566 source.n368 a_n3202_n3288# 0.012759f
C567 source.n369 a_n3202_n3288# 0.030157f
C568 source.n370 a_n3202_n3288# 0.013509f
C569 source.n371 a_n3202_n3288# 0.023743f
C570 source.n372 a_n3202_n3288# 0.012759f
C571 source.n373 a_n3202_n3288# 0.022618f
C572 source.n374 a_n3202_n3288# 0.021319f
C573 source.t39 a_n3202_n3288# 0.050933f
C574 source.n375 a_n3202_n3288# 0.171186f
C575 source.n376 a_n3202_n3288# 1.19781f
C576 source.n377 a_n3202_n3288# 0.012759f
C577 source.n378 a_n3202_n3288# 0.013509f
C578 source.n379 a_n3202_n3288# 0.030157f
C579 source.n380 a_n3202_n3288# 0.030157f
C580 source.n381 a_n3202_n3288# 0.013509f
C581 source.n382 a_n3202_n3288# 0.012759f
C582 source.n383 a_n3202_n3288# 0.023743f
C583 source.n384 a_n3202_n3288# 0.023743f
C584 source.n385 a_n3202_n3288# 0.012759f
C585 source.n386 a_n3202_n3288# 0.013509f
C586 source.n387 a_n3202_n3288# 0.030157f
C587 source.n388 a_n3202_n3288# 0.030157f
C588 source.n389 a_n3202_n3288# 0.013509f
C589 source.n390 a_n3202_n3288# 0.012759f
C590 source.n391 a_n3202_n3288# 0.023743f
C591 source.n392 a_n3202_n3288# 0.023743f
C592 source.n393 a_n3202_n3288# 0.012759f
C593 source.n394 a_n3202_n3288# 0.012759f
C594 source.n395 a_n3202_n3288# 0.013509f
C595 source.n396 a_n3202_n3288# 0.030157f
C596 source.n397 a_n3202_n3288# 0.030157f
C597 source.n398 a_n3202_n3288# 0.030157f
C598 source.n399 a_n3202_n3288# 0.013134f
C599 source.n400 a_n3202_n3288# 0.012759f
C600 source.n401 a_n3202_n3288# 0.023743f
C601 source.n402 a_n3202_n3288# 0.023743f
C602 source.n403 a_n3202_n3288# 0.012759f
C603 source.n404 a_n3202_n3288# 0.013509f
C604 source.n405 a_n3202_n3288# 0.030157f
C605 source.n406 a_n3202_n3288# 0.030157f
C606 source.n407 a_n3202_n3288# 0.013509f
C607 source.n408 a_n3202_n3288# 0.012759f
C608 source.n409 a_n3202_n3288# 0.023743f
C609 source.n410 a_n3202_n3288# 0.023743f
C610 source.n411 a_n3202_n3288# 0.012759f
C611 source.n412 a_n3202_n3288# 0.013509f
C612 source.n413 a_n3202_n3288# 0.030157f
C613 source.n414 a_n3202_n3288# 0.061885f
C614 source.n415 a_n3202_n3288# 0.013509f
C615 source.n416 a_n3202_n3288# 0.012759f
C616 source.n417 a_n3202_n3288# 0.050989f
C617 source.n418 a_n3202_n3288# 0.034154f
C618 source.n419 a_n3202_n3288# 0.128558f
C619 source.n420 a_n3202_n3288# 0.031451f
C620 source.n421 a_n3202_n3288# 0.023743f
C621 source.n422 a_n3202_n3288# 0.012759f
C622 source.n423 a_n3202_n3288# 0.030157f
C623 source.n424 a_n3202_n3288# 0.013509f
C624 source.n425 a_n3202_n3288# 0.023743f
C625 source.n426 a_n3202_n3288# 0.012759f
C626 source.n427 a_n3202_n3288# 0.030157f
C627 source.n428 a_n3202_n3288# 0.013509f
C628 source.n429 a_n3202_n3288# 0.023743f
C629 source.n430 a_n3202_n3288# 0.013134f
C630 source.n431 a_n3202_n3288# 0.030157f
C631 source.n432 a_n3202_n3288# 0.013509f
C632 source.n433 a_n3202_n3288# 0.023743f
C633 source.n434 a_n3202_n3288# 0.012759f
C634 source.n435 a_n3202_n3288# 0.030157f
C635 source.n436 a_n3202_n3288# 0.013509f
C636 source.n437 a_n3202_n3288# 0.023743f
C637 source.n438 a_n3202_n3288# 0.012759f
C638 source.n439 a_n3202_n3288# 0.022618f
C639 source.n440 a_n3202_n3288# 0.021319f
C640 source.t28 a_n3202_n3288# 0.050933f
C641 source.n441 a_n3202_n3288# 0.171186f
C642 source.n442 a_n3202_n3288# 1.19781f
C643 source.n443 a_n3202_n3288# 0.012759f
C644 source.n444 a_n3202_n3288# 0.013509f
C645 source.n445 a_n3202_n3288# 0.030157f
C646 source.n446 a_n3202_n3288# 0.030157f
C647 source.n447 a_n3202_n3288# 0.013509f
C648 source.n448 a_n3202_n3288# 0.012759f
C649 source.n449 a_n3202_n3288# 0.023743f
C650 source.n450 a_n3202_n3288# 0.023743f
C651 source.n451 a_n3202_n3288# 0.012759f
C652 source.n452 a_n3202_n3288# 0.013509f
C653 source.n453 a_n3202_n3288# 0.030157f
C654 source.n454 a_n3202_n3288# 0.030157f
C655 source.n455 a_n3202_n3288# 0.013509f
C656 source.n456 a_n3202_n3288# 0.012759f
C657 source.n457 a_n3202_n3288# 0.023743f
C658 source.n458 a_n3202_n3288# 0.023743f
C659 source.n459 a_n3202_n3288# 0.012759f
C660 source.n460 a_n3202_n3288# 0.012759f
C661 source.n461 a_n3202_n3288# 0.013509f
C662 source.n462 a_n3202_n3288# 0.030157f
C663 source.n463 a_n3202_n3288# 0.030157f
C664 source.n464 a_n3202_n3288# 0.030157f
C665 source.n465 a_n3202_n3288# 0.013134f
C666 source.n466 a_n3202_n3288# 0.012759f
C667 source.n467 a_n3202_n3288# 0.023743f
C668 source.n468 a_n3202_n3288# 0.023743f
C669 source.n469 a_n3202_n3288# 0.012759f
C670 source.n470 a_n3202_n3288# 0.013509f
C671 source.n471 a_n3202_n3288# 0.030157f
C672 source.n472 a_n3202_n3288# 0.030157f
C673 source.n473 a_n3202_n3288# 0.013509f
C674 source.n474 a_n3202_n3288# 0.012759f
C675 source.n475 a_n3202_n3288# 0.023743f
C676 source.n476 a_n3202_n3288# 0.023743f
C677 source.n477 a_n3202_n3288# 0.012759f
C678 source.n478 a_n3202_n3288# 0.013509f
C679 source.n479 a_n3202_n3288# 0.030157f
C680 source.n480 a_n3202_n3288# 0.061885f
C681 source.n481 a_n3202_n3288# 0.013509f
C682 source.n482 a_n3202_n3288# 0.012759f
C683 source.n483 a_n3202_n3288# 0.050989f
C684 source.n484 a_n3202_n3288# 0.034154f
C685 source.n485 a_n3202_n3288# 0.128558f
C686 source.t23 a_n3202_n3288# 0.225152f
C687 source.t33 a_n3202_n3288# 0.225152f
C688 source.n486 a_n3202_n3288# 1.92775f
C689 source.n487 a_n3202_n3288# 0.391812f
C690 source.t29 a_n3202_n3288# 0.225152f
C691 source.t37 a_n3202_n3288# 0.225152f
C692 source.n488 a_n3202_n3288# 1.92775f
C693 source.n489 a_n3202_n3288# 0.391812f
C694 source.t25 a_n3202_n3288# 0.225152f
C695 source.t21 a_n3202_n3288# 0.225152f
C696 source.n490 a_n3202_n3288# 1.92775f
C697 source.n491 a_n3202_n3288# 0.391812f
C698 source.t38 a_n3202_n3288# 0.225152f
C699 source.t20 a_n3202_n3288# 0.225152f
C700 source.n492 a_n3202_n3288# 1.92775f
C701 source.n493 a_n3202_n3288# 0.391812f
C702 source.n494 a_n3202_n3288# 0.031451f
C703 source.n495 a_n3202_n3288# 0.023743f
C704 source.n496 a_n3202_n3288# 0.012759f
C705 source.n497 a_n3202_n3288# 0.030157f
C706 source.n498 a_n3202_n3288# 0.013509f
C707 source.n499 a_n3202_n3288# 0.023743f
C708 source.n500 a_n3202_n3288# 0.012759f
C709 source.n501 a_n3202_n3288# 0.030157f
C710 source.n502 a_n3202_n3288# 0.013509f
C711 source.n503 a_n3202_n3288# 0.023743f
C712 source.n504 a_n3202_n3288# 0.013134f
C713 source.n505 a_n3202_n3288# 0.030157f
C714 source.n506 a_n3202_n3288# 0.013509f
C715 source.n507 a_n3202_n3288# 0.023743f
C716 source.n508 a_n3202_n3288# 0.012759f
C717 source.n509 a_n3202_n3288# 0.030157f
C718 source.n510 a_n3202_n3288# 0.013509f
C719 source.n511 a_n3202_n3288# 0.023743f
C720 source.n512 a_n3202_n3288# 0.012759f
C721 source.n513 a_n3202_n3288# 0.022618f
C722 source.n514 a_n3202_n3288# 0.021319f
C723 source.t22 a_n3202_n3288# 0.050933f
C724 source.n515 a_n3202_n3288# 0.171186f
C725 source.n516 a_n3202_n3288# 1.19781f
C726 source.n517 a_n3202_n3288# 0.012759f
C727 source.n518 a_n3202_n3288# 0.013509f
C728 source.n519 a_n3202_n3288# 0.030157f
C729 source.n520 a_n3202_n3288# 0.030157f
C730 source.n521 a_n3202_n3288# 0.013509f
C731 source.n522 a_n3202_n3288# 0.012759f
C732 source.n523 a_n3202_n3288# 0.023743f
C733 source.n524 a_n3202_n3288# 0.023743f
C734 source.n525 a_n3202_n3288# 0.012759f
C735 source.n526 a_n3202_n3288# 0.013509f
C736 source.n527 a_n3202_n3288# 0.030157f
C737 source.n528 a_n3202_n3288# 0.030157f
C738 source.n529 a_n3202_n3288# 0.013509f
C739 source.n530 a_n3202_n3288# 0.012759f
C740 source.n531 a_n3202_n3288# 0.023743f
C741 source.n532 a_n3202_n3288# 0.023743f
C742 source.n533 a_n3202_n3288# 0.012759f
C743 source.n534 a_n3202_n3288# 0.012759f
C744 source.n535 a_n3202_n3288# 0.013509f
C745 source.n536 a_n3202_n3288# 0.030157f
C746 source.n537 a_n3202_n3288# 0.030157f
C747 source.n538 a_n3202_n3288# 0.030157f
C748 source.n539 a_n3202_n3288# 0.013134f
C749 source.n540 a_n3202_n3288# 0.012759f
C750 source.n541 a_n3202_n3288# 0.023743f
C751 source.n542 a_n3202_n3288# 0.023743f
C752 source.n543 a_n3202_n3288# 0.012759f
C753 source.n544 a_n3202_n3288# 0.013509f
C754 source.n545 a_n3202_n3288# 0.030157f
C755 source.n546 a_n3202_n3288# 0.030157f
C756 source.n547 a_n3202_n3288# 0.013509f
C757 source.n548 a_n3202_n3288# 0.012759f
C758 source.n549 a_n3202_n3288# 0.023743f
C759 source.n550 a_n3202_n3288# 0.023743f
C760 source.n551 a_n3202_n3288# 0.012759f
C761 source.n552 a_n3202_n3288# 0.013509f
C762 source.n553 a_n3202_n3288# 0.030157f
C763 source.n554 a_n3202_n3288# 0.061885f
C764 source.n555 a_n3202_n3288# 0.013509f
C765 source.n556 a_n3202_n3288# 0.012759f
C766 source.n557 a_n3202_n3288# 0.050989f
C767 source.n558 a_n3202_n3288# 0.034154f
C768 source.n559 a_n3202_n3288# 0.288577f
C769 source.n560 a_n3202_n3288# 1.50841f
C770 minus.n0 a_n3202_n3288# 0.037669f
C771 minus.n1 a_n3202_n3288# 0.008548f
C772 minus.t12 a_n3202_n3288# 1.03116f
C773 minus.n2 a_n3202_n3288# 0.062742f
C774 minus.t10 a_n3202_n3288# 1.03116f
C775 minus.n3 a_n3202_n3288# 0.407803f
C776 minus.n4 a_n3202_n3288# 0.037669f
C777 minus.t11 a_n3202_n3288# 1.03116f
C778 minus.n5 a_n3202_n3288# 0.418557f
C779 minus.n6 a_n3202_n3288# 0.173388f
C780 minus.t9 a_n3202_n3288# 1.05182f
C781 minus.n7 a_n3202_n3288# 0.392977f
C782 minus.t7 a_n3202_n3288# 1.03116f
C783 minus.n8 a_n3202_n3288# 0.410969f
C784 minus.n9 a_n3202_n3288# 0.008548f
C785 minus.t6 a_n3202_n3288# 1.03116f
C786 minus.n10 a_n3202_n3288# 0.418093f
C787 minus.n11 a_n3202_n3288# 0.062742f
C788 minus.n12 a_n3202_n3288# 0.062742f
C789 minus.n13 a_n3202_n3288# 0.050264f
C790 minus.n14 a_n3202_n3288# 0.008548f
C791 minus.t13 a_n3202_n3288# 1.03116f
C792 minus.n15 a_n3202_n3288# 0.407803f
C793 minus.n16 a_n3202_n3288# 0.008548f
C794 minus.n17 a_n3202_n3288# 0.037669f
C795 minus.n18 a_n3202_n3288# 0.037669f
C796 minus.n19 a_n3202_n3288# 0.050264f
C797 minus.n20 a_n3202_n3288# 0.008548f
C798 minus.t8 a_n3202_n3288# 1.03116f
C799 minus.n21 a_n3202_n3288# 0.418557f
C800 minus.t17 a_n3202_n3288# 1.03116f
C801 minus.n22 a_n3202_n3288# 0.418093f
C802 minus.n23 a_n3202_n3288# 0.062742f
C803 minus.n24 a_n3202_n3288# 0.050264f
C804 minus.n25 a_n3202_n3288# 0.037669f
C805 minus.n26 a_n3202_n3288# 0.407803f
C806 minus.n27 a_n3202_n3288# 0.008548f
C807 minus.t4 a_n3202_n3288# 1.03116f
C808 minus.n28 a_n3202_n3288# 0.407455f
C809 minus.n29 a_n3202_n3288# 1.64156f
C810 minus.n30 a_n3202_n3288# 0.037669f
C811 minus.n31 a_n3202_n3288# 0.008548f
C812 minus.n32 a_n3202_n3288# 0.062742f
C813 minus.t2 a_n3202_n3288# 1.03116f
C814 minus.n33 a_n3202_n3288# 0.407803f
C815 minus.n34 a_n3202_n3288# 0.037669f
C816 minus.t3 a_n3202_n3288# 1.03116f
C817 minus.n35 a_n3202_n3288# 0.418557f
C818 minus.n36 a_n3202_n3288# 0.173388f
C819 minus.t19 a_n3202_n3288# 1.05182f
C820 minus.n37 a_n3202_n3288# 0.392977f
C821 minus.t5 a_n3202_n3288# 1.03116f
C822 minus.n38 a_n3202_n3288# 0.410969f
C823 minus.n39 a_n3202_n3288# 0.008548f
C824 minus.t16 a_n3202_n3288# 1.03116f
C825 minus.n40 a_n3202_n3288# 0.418093f
C826 minus.n41 a_n3202_n3288# 0.062742f
C827 minus.n42 a_n3202_n3288# 0.062742f
C828 minus.n43 a_n3202_n3288# 0.050264f
C829 minus.n44 a_n3202_n3288# 0.008548f
C830 minus.t18 a_n3202_n3288# 1.03116f
C831 minus.n45 a_n3202_n3288# 0.407803f
C832 minus.n46 a_n3202_n3288# 0.008548f
C833 minus.n47 a_n3202_n3288# 0.037669f
C834 minus.n48 a_n3202_n3288# 0.037669f
C835 minus.n49 a_n3202_n3288# 0.050264f
C836 minus.n50 a_n3202_n3288# 0.008548f
C837 minus.t14 a_n3202_n3288# 1.03116f
C838 minus.n51 a_n3202_n3288# 0.418557f
C839 minus.t0 a_n3202_n3288# 1.03116f
C840 minus.n52 a_n3202_n3288# 0.418093f
C841 minus.n53 a_n3202_n3288# 0.062742f
C842 minus.n54 a_n3202_n3288# 0.050264f
C843 minus.n55 a_n3202_n3288# 0.037669f
C844 minus.t15 a_n3202_n3288# 1.03116f
C845 minus.n56 a_n3202_n3288# 0.407803f
C846 minus.n57 a_n3202_n3288# 0.008548f
C847 minus.t1 a_n3202_n3288# 1.03116f
C848 minus.n58 a_n3202_n3288# 0.407455f
C849 minus.n59 a_n3202_n3288# 0.264293f
C850 minus.n60 a_n3202_n3288# 1.95906f
.ends

