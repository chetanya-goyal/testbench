* NGSPICE file created from diffpair376.ext - technology: sky130A

.subckt diffpair376 minus drain_right drain_left source plus
X0 drain_left.t13 plus.t0 source.t20 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X1 source.t24 plus.t1 drain_left.t12 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X2 drain_right.t13 minus.t0 source.t4 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X3 drain_right.t12 minus.t1 source.t7 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X4 drain_right.t11 minus.t2 source.t10 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X5 source.t25 plus.t2 drain_left.t11 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X6 source.t3 minus.t3 drain_right.t10 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X7 drain_right.t9 minus.t4 source.t8 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X8 drain_right.t8 minus.t5 source.t9 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X9 drain_left.t10 plus.t3 source.t17 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X10 drain_left.t9 plus.t4 source.t15 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X11 drain_left.t8 plus.t5 source.t18 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X12 source.t0 minus.t6 drain_right.t7 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X13 drain_right.t6 minus.t7 source.t1 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X14 a_n2204_n2688# a_n2204_n2688# a_n2204_n2688# a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.6
X15 source.t26 plus.t6 drain_left.t7 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X16 source.t2 minus.t8 drain_right.t5 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X17 a_n2204_n2688# a_n2204_n2688# a_n2204_n2688# a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X18 drain_left.t6 plus.t7 source.t19 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X19 drain_right.t4 minus.t9 source.t11 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X20 a_n2204_n2688# a_n2204_n2688# a_n2204_n2688# a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X21 source.t16 plus.t8 drain_left.t5 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X22 drain_left.t4 plus.t9 source.t21 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X23 a_n2204_n2688# a_n2204_n2688# a_n2204_n2688# a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X24 source.t27 minus.t10 drain_right.t3 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X25 drain_left.t3 plus.t10 source.t14 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X26 source.t13 plus.t11 drain_left.t2 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X27 source.t6 minus.t11 drain_right.t2 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X28 drain_left.t1 plus.t12 source.t22 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X29 drain_right.t1 minus.t12 source.t5 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X30 source.t12 minus.t13 drain_right.t0 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X31 source.t23 plus.t13 drain_left.t0 a_n2204_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
R0 plus.n5 plus.t9 450.818
R1 plus.n23 plus.t10 450.818
R2 plus.n16 plus.t0 426.973
R3 plus.n14 plus.t1 426.973
R4 plus.n2 plus.t3 426.973
R5 plus.n9 plus.t6 426.973
R6 plus.n8 plus.t7 426.973
R7 plus.n4 plus.t8 426.973
R8 plus.n34 plus.t5 426.973
R9 plus.n32 plus.t13 426.973
R10 plus.n20 plus.t12 426.973
R11 plus.n27 plus.t11 426.973
R12 plus.n26 plus.t4 426.973
R13 plus.n22 plus.t2 426.973
R14 plus.n7 plus.n6 161.3
R15 plus.n8 plus.n3 161.3
R16 plus.n11 plus.n2 161.3
R17 plus.n13 plus.n12 161.3
R18 plus.n14 plus.n1 161.3
R19 plus.n15 plus.n0 161.3
R20 plus.n17 plus.n16 161.3
R21 plus.n25 plus.n24 161.3
R22 plus.n26 plus.n21 161.3
R23 plus.n29 plus.n20 161.3
R24 plus.n31 plus.n30 161.3
R25 plus.n32 plus.n19 161.3
R26 plus.n33 plus.n18 161.3
R27 plus.n35 plus.n34 161.3
R28 plus.n10 plus.n9 80.6037
R29 plus.n28 plus.n27 80.6037
R30 plus.n9 plus.n2 48.2005
R31 plus.n9 plus.n8 48.2005
R32 plus.n27 plus.n20 48.2005
R33 plus.n27 plus.n26 48.2005
R34 plus.n14 plus.n13 45.2793
R35 plus.n7 plus.n4 45.2793
R36 plus.n32 plus.n31 45.2793
R37 plus.n25 plus.n22 45.2793
R38 plus.n24 plus.n23 44.9119
R39 plus.n6 plus.n5 44.9119
R40 plus.n16 plus.n15 35.055
R41 plus.n34 plus.n33 35.055
R42 plus plus.n35 30.2888
R43 plus.n23 plus.n22 17.739
R44 plus.n5 plus.n4 17.739
R45 plus.n15 plus.n14 13.146
R46 plus.n33 plus.n32 13.146
R47 plus plus.n17 11.0819
R48 plus.n13 plus.n2 2.92171
R49 plus.n8 plus.n7 2.92171
R50 plus.n31 plus.n20 2.92171
R51 plus.n26 plus.n25 2.92171
R52 plus.n10 plus.n3 0.285035
R53 plus.n11 plus.n10 0.285035
R54 plus.n29 plus.n28 0.285035
R55 plus.n28 plus.n21 0.285035
R56 plus.n6 plus.n3 0.189894
R57 plus.n12 plus.n11 0.189894
R58 plus.n12 plus.n1 0.189894
R59 plus.n1 plus.n0 0.189894
R60 plus.n17 plus.n0 0.189894
R61 plus.n35 plus.n18 0.189894
R62 plus.n19 plus.n18 0.189894
R63 plus.n30 plus.n19 0.189894
R64 plus.n30 plus.n29 0.189894
R65 plus.n24 plus.n21 0.189894
R66 source.n7 source.t11 51.0588
R67 source.n27 source.t8 51.0586
R68 source.n20 source.t14 51.0586
R69 source.n0 source.t20 51.0586
R70 source.n2 source.n1 48.8588
R71 source.n4 source.n3 48.8588
R72 source.n6 source.n5 48.8588
R73 source.n9 source.n8 48.8588
R74 source.n11 source.n10 48.8588
R75 source.n13 source.n12 48.8588
R76 source.n26 source.n25 48.8586
R77 source.n24 source.n23 48.8586
R78 source.n22 source.n21 48.8586
R79 source.n19 source.n18 48.8586
R80 source.n17 source.n16 48.8586
R81 source.n15 source.n14 48.8586
R82 source.n15 source.n13 20.6184
R83 source.n28 source.n0 14.1529
R84 source.n28 source.n27 5.66429
R85 source.n25 source.t5 2.2005
R86 source.n25 source.t6 2.2005
R87 source.n23 source.t4 2.2005
R88 source.n23 source.t27 2.2005
R89 source.n21 source.t9 2.2005
R90 source.n21 source.t12 2.2005
R91 source.n18 source.t15 2.2005
R92 source.n18 source.t25 2.2005
R93 source.n16 source.t22 2.2005
R94 source.n16 source.t13 2.2005
R95 source.n14 source.t18 2.2005
R96 source.n14 source.t23 2.2005
R97 source.n1 source.t17 2.2005
R98 source.n1 source.t24 2.2005
R99 source.n3 source.t19 2.2005
R100 source.n3 source.t26 2.2005
R101 source.n5 source.t21 2.2005
R102 source.n5 source.t16 2.2005
R103 source.n8 source.t1 2.2005
R104 source.n8 source.t2 2.2005
R105 source.n10 source.t7 2.2005
R106 source.n10 source.t0 2.2005
R107 source.n12 source.t10 2.2005
R108 source.n12 source.t3 2.2005
R109 source.n7 source.n6 0.87119
R110 source.n22 source.n20 0.87119
R111 source.n13 source.n11 0.802224
R112 source.n11 source.n9 0.802224
R113 source.n9 source.n7 0.802224
R114 source.n6 source.n4 0.802224
R115 source.n4 source.n2 0.802224
R116 source.n2 source.n0 0.802224
R117 source.n17 source.n15 0.802224
R118 source.n19 source.n17 0.802224
R119 source.n20 source.n19 0.802224
R120 source.n24 source.n22 0.802224
R121 source.n26 source.n24 0.802224
R122 source.n27 source.n26 0.802224
R123 source source.n28 0.188
R124 drain_left.n7 drain_left.t4 68.5393
R125 drain_left.n1 drain_left.t8 68.5391
R126 drain_left.n4 drain_left.n2 66.3391
R127 drain_left.n9 drain_left.n8 65.5376
R128 drain_left.n7 drain_left.n6 65.5376
R129 drain_left.n11 drain_left.n10 65.5374
R130 drain_left.n4 drain_left.n3 65.5373
R131 drain_left.n1 drain_left.n0 65.5373
R132 drain_left drain_left.n5 29.7043
R133 drain_left drain_left.n11 6.45494
R134 drain_left.n2 drain_left.t11 2.2005
R135 drain_left.n2 drain_left.t3 2.2005
R136 drain_left.n3 drain_left.t2 2.2005
R137 drain_left.n3 drain_left.t9 2.2005
R138 drain_left.n0 drain_left.t0 2.2005
R139 drain_left.n0 drain_left.t1 2.2005
R140 drain_left.n10 drain_left.t12 2.2005
R141 drain_left.n10 drain_left.t13 2.2005
R142 drain_left.n8 drain_left.t7 2.2005
R143 drain_left.n8 drain_left.t10 2.2005
R144 drain_left.n6 drain_left.t5 2.2005
R145 drain_left.n6 drain_left.t6 2.2005
R146 drain_left.n9 drain_left.n7 0.802224
R147 drain_left.n11 drain_left.n9 0.802224
R148 drain_left.n5 drain_left.n1 0.546447
R149 drain_left.n5 drain_left.n4 0.145585
R150 minus.n5 minus.t9 450.818
R151 minus.n23 minus.t5 450.818
R152 minus.n4 minus.t8 426.973
R153 minus.n8 minus.t7 426.973
R154 minus.n9 minus.t6 426.973
R155 minus.n10 minus.t1 426.973
R156 minus.n14 minus.t3 426.973
R157 minus.n16 minus.t2 426.973
R158 minus.n22 minus.t13 426.973
R159 minus.n26 minus.t0 426.973
R160 minus.n27 minus.t10 426.973
R161 minus.n28 minus.t12 426.973
R162 minus.n32 minus.t11 426.973
R163 minus.n34 minus.t4 426.973
R164 minus.n17 minus.n16 161.3
R165 minus.n15 minus.n0 161.3
R166 minus.n14 minus.n13 161.3
R167 minus.n12 minus.n1 161.3
R168 minus.n11 minus.n10 161.3
R169 minus.n8 minus.n7 161.3
R170 minus.n6 minus.n3 161.3
R171 minus.n35 minus.n34 161.3
R172 minus.n33 minus.n18 161.3
R173 minus.n32 minus.n31 161.3
R174 minus.n30 minus.n19 161.3
R175 minus.n29 minus.n28 161.3
R176 minus.n26 minus.n25 161.3
R177 minus.n24 minus.n21 161.3
R178 minus.n9 minus.n2 80.6037
R179 minus.n27 minus.n20 80.6037
R180 minus.n9 minus.n8 48.2005
R181 minus.n10 minus.n9 48.2005
R182 minus.n27 minus.n26 48.2005
R183 minus.n28 minus.n27 48.2005
R184 minus.n4 minus.n3 45.2793
R185 minus.n14 minus.n1 45.2793
R186 minus.n22 minus.n21 45.2793
R187 minus.n32 minus.n19 45.2793
R188 minus.n6 minus.n5 44.9119
R189 minus.n24 minus.n23 44.9119
R190 minus.n36 minus.n17 35.2713
R191 minus.n16 minus.n15 35.055
R192 minus.n34 minus.n33 35.055
R193 minus.n5 minus.n4 17.739
R194 minus.n23 minus.n22 17.739
R195 minus.n15 minus.n14 13.146
R196 minus.n33 minus.n32 13.146
R197 minus.n36 minus.n35 6.57436
R198 minus.n8 minus.n3 2.92171
R199 minus.n10 minus.n1 2.92171
R200 minus.n26 minus.n21 2.92171
R201 minus.n28 minus.n19 2.92171
R202 minus.n11 minus.n2 0.285035
R203 minus.n7 minus.n2 0.285035
R204 minus.n25 minus.n20 0.285035
R205 minus.n29 minus.n20 0.285035
R206 minus.n17 minus.n0 0.189894
R207 minus.n13 minus.n0 0.189894
R208 minus.n13 minus.n12 0.189894
R209 minus.n12 minus.n11 0.189894
R210 minus.n7 minus.n6 0.189894
R211 minus.n25 minus.n24 0.189894
R212 minus.n30 minus.n29 0.189894
R213 minus.n31 minus.n30 0.189894
R214 minus.n31 minus.n18 0.189894
R215 minus.n35 minus.n18 0.189894
R216 minus minus.n36 0.188
R217 drain_right.n1 drain_right.t8 68.5391
R218 drain_right.n11 drain_right.t11 67.7376
R219 drain_right.n8 drain_right.n6 66.3391
R220 drain_right.n4 drain_right.n2 66.3391
R221 drain_right.n8 drain_right.n7 65.5376
R222 drain_right.n10 drain_right.n9 65.5376
R223 drain_right.n4 drain_right.n3 65.5373
R224 drain_right.n1 drain_right.n0 65.5373
R225 drain_right drain_right.n5 29.151
R226 drain_right drain_right.n11 6.05408
R227 drain_right.n2 drain_right.t2 2.2005
R228 drain_right.n2 drain_right.t9 2.2005
R229 drain_right.n3 drain_right.t3 2.2005
R230 drain_right.n3 drain_right.t1 2.2005
R231 drain_right.n0 drain_right.t0 2.2005
R232 drain_right.n0 drain_right.t13 2.2005
R233 drain_right.n6 drain_right.t5 2.2005
R234 drain_right.n6 drain_right.t4 2.2005
R235 drain_right.n7 drain_right.t7 2.2005
R236 drain_right.n7 drain_right.t6 2.2005
R237 drain_right.n9 drain_right.t10 2.2005
R238 drain_right.n9 drain_right.t12 2.2005
R239 drain_right.n11 drain_right.n10 0.802224
R240 drain_right.n10 drain_right.n8 0.802224
R241 drain_right.n5 drain_right.n1 0.546447
R242 drain_right.n5 drain_right.n4 0.145585
C0 source minus 6.36834f
C1 drain_left minus 0.172803f
C2 source drain_left 15.809299f
C3 drain_right plus 0.374006f
C4 plus minus 5.34269f
C5 source plus 6.38278f
C6 drain_left plus 6.5649f
C7 drain_right minus 6.35021f
C8 source drain_right 15.8041f
C9 drain_left drain_right 1.14729f
C10 drain_right a_n2204_n2688# 6.60876f
C11 drain_left a_n2204_n2688# 6.94194f
C12 source a_n2204_n2688# 5.497022f
C13 minus a_n2204_n2688# 8.516848f
C14 plus a_n2204_n2688# 10.13763f
C15 drain_right.t8 a_n2204_n2688# 2.0428f
C16 drain_right.t0 a_n2204_n2688# 0.183115f
C17 drain_right.t13 a_n2204_n2688# 0.183115f
C18 drain_right.n0 a_n2204_n2688# 1.60164f
C19 drain_right.n1 a_n2204_n2688# 0.660508f
C20 drain_right.t2 a_n2204_n2688# 0.183115f
C21 drain_right.t9 a_n2204_n2688# 0.183115f
C22 drain_right.n2 a_n2204_n2688# 1.60587f
C23 drain_right.t3 a_n2204_n2688# 0.183115f
C24 drain_right.t1 a_n2204_n2688# 0.183115f
C25 drain_right.n3 a_n2204_n2688# 1.60164f
C26 drain_right.n4 a_n2204_n2688# 0.634309f
C27 drain_right.n5 a_n2204_n2688# 1.14601f
C28 drain_right.t5 a_n2204_n2688# 0.183115f
C29 drain_right.t4 a_n2204_n2688# 0.183115f
C30 drain_right.n6 a_n2204_n2688# 1.60587f
C31 drain_right.t7 a_n2204_n2688# 0.183115f
C32 drain_right.t6 a_n2204_n2688# 0.183115f
C33 drain_right.n7 a_n2204_n2688# 1.60165f
C34 drain_right.n8 a_n2204_n2688# 0.684672f
C35 drain_right.t10 a_n2204_n2688# 0.183115f
C36 drain_right.t12 a_n2204_n2688# 0.183115f
C37 drain_right.n9 a_n2204_n2688# 1.60165f
C38 drain_right.n10 a_n2204_n2688# 0.33926f
C39 drain_right.t11 a_n2204_n2688# 2.03876f
C40 drain_right.n11 a_n2204_n2688# 0.57662f
C41 minus.n0 a_n2204_n2688# 0.043533f
C42 minus.n1 a_n2204_n2688# 0.009879f
C43 minus.t3 a_n2204_n2688# 0.674176f
C44 minus.n2 a_n2204_n2688# 0.057954f
C45 minus.n3 a_n2204_n2688# 0.009879f
C46 minus.t7 a_n2204_n2688# 0.674176f
C47 minus.t9 a_n2204_n2688# 0.689229f
C48 minus.t8 a_n2204_n2688# 0.674176f
C49 minus.n4 a_n2204_n2688# 0.292627f
C50 minus.n5 a_n2204_n2688# 0.273238f
C51 minus.n6 a_n2204_n2688# 0.178099f
C52 minus.n7 a_n2204_n2688# 0.05809f
C53 minus.n8 a_n2204_n2688# 0.285893f
C54 minus.t6 a_n2204_n2688# 0.674176f
C55 minus.n9 a_n2204_n2688# 0.295235f
C56 minus.t1 a_n2204_n2688# 0.674176f
C57 minus.n10 a_n2204_n2688# 0.285893f
C58 minus.n11 a_n2204_n2688# 0.05809f
C59 minus.n12 a_n2204_n2688# 0.043533f
C60 minus.n13 a_n2204_n2688# 0.043533f
C61 minus.n14 a_n2204_n2688# 0.287235f
C62 minus.n15 a_n2204_n2688# 0.009879f
C63 minus.t2 a_n2204_n2688# 0.674176f
C64 minus.n16 a_n2204_n2688# 0.28294f
C65 minus.n17 a_n2204_n2688# 1.47987f
C66 minus.n18 a_n2204_n2688# 0.043533f
C67 minus.n19 a_n2204_n2688# 0.009879f
C68 minus.n20 a_n2204_n2688# 0.057954f
C69 minus.n21 a_n2204_n2688# 0.009879f
C70 minus.t5 a_n2204_n2688# 0.689229f
C71 minus.t13 a_n2204_n2688# 0.674176f
C72 minus.n22 a_n2204_n2688# 0.292627f
C73 minus.n23 a_n2204_n2688# 0.273238f
C74 minus.n24 a_n2204_n2688# 0.178099f
C75 minus.n25 a_n2204_n2688# 0.05809f
C76 minus.t0 a_n2204_n2688# 0.674176f
C77 minus.n26 a_n2204_n2688# 0.285893f
C78 minus.t10 a_n2204_n2688# 0.674176f
C79 minus.n27 a_n2204_n2688# 0.295235f
C80 minus.t12 a_n2204_n2688# 0.674176f
C81 minus.n28 a_n2204_n2688# 0.285893f
C82 minus.n29 a_n2204_n2688# 0.05809f
C83 minus.n30 a_n2204_n2688# 0.043533f
C84 minus.n31 a_n2204_n2688# 0.043533f
C85 minus.t11 a_n2204_n2688# 0.674176f
C86 minus.n32 a_n2204_n2688# 0.287235f
C87 minus.n33 a_n2204_n2688# 0.009879f
C88 minus.t4 a_n2204_n2688# 0.674176f
C89 minus.n34 a_n2204_n2688# 0.28294f
C90 minus.n35 a_n2204_n2688# 0.292209f
C91 minus.n36 a_n2204_n2688# 1.79971f
C92 drain_left.t8 a_n2204_n2688# 2.05189f
C93 drain_left.t0 a_n2204_n2688# 0.18393f
C94 drain_left.t1 a_n2204_n2688# 0.18393f
C95 drain_left.n0 a_n2204_n2688# 1.60877f
C96 drain_left.n1 a_n2204_n2688# 0.663449f
C97 drain_left.t11 a_n2204_n2688# 0.18393f
C98 drain_left.t3 a_n2204_n2688# 0.18393f
C99 drain_left.n2 a_n2204_n2688# 1.61302f
C100 drain_left.t2 a_n2204_n2688# 0.18393f
C101 drain_left.t9 a_n2204_n2688# 0.18393f
C102 drain_left.n3 a_n2204_n2688# 1.60877f
C103 drain_left.n4 a_n2204_n2688# 0.637133f
C104 drain_left.n5 a_n2204_n2688# 1.20402f
C105 drain_left.t4 a_n2204_n2688# 2.05189f
C106 drain_left.t5 a_n2204_n2688# 0.18393f
C107 drain_left.t6 a_n2204_n2688# 0.18393f
C108 drain_left.n6 a_n2204_n2688# 1.60878f
C109 drain_left.n7 a_n2204_n2688# 0.683659f
C110 drain_left.t7 a_n2204_n2688# 0.18393f
C111 drain_left.t10 a_n2204_n2688# 0.18393f
C112 drain_left.n8 a_n2204_n2688# 1.60878f
C113 drain_left.n9 a_n2204_n2688# 0.34077f
C114 drain_left.t12 a_n2204_n2688# 0.18393f
C115 drain_left.t13 a_n2204_n2688# 0.18393f
C116 drain_left.n10 a_n2204_n2688# 1.60877f
C117 drain_left.n11 a_n2204_n2688# 0.566289f
C118 source.t20 a_n2204_n2688# 2.09145f
C119 source.n0 a_n2204_n2688# 1.24108f
C120 source.t17 a_n2204_n2688# 0.196132f
C121 source.t24 a_n2204_n2688# 0.196132f
C122 source.n1 a_n2204_n2688# 1.64189f
C123 source.n2 a_n2204_n2688# 0.399509f
C124 source.t19 a_n2204_n2688# 0.196132f
C125 source.t26 a_n2204_n2688# 0.196132f
C126 source.n3 a_n2204_n2688# 1.64189f
C127 source.n4 a_n2204_n2688# 0.399509f
C128 source.t21 a_n2204_n2688# 0.196132f
C129 source.t16 a_n2204_n2688# 0.196132f
C130 source.n5 a_n2204_n2688# 1.64189f
C131 source.n6 a_n2204_n2688# 0.405637f
C132 source.t11 a_n2204_n2688# 2.09145f
C133 source.n7 a_n2204_n2688# 0.49098f
C134 source.t1 a_n2204_n2688# 0.196132f
C135 source.t2 a_n2204_n2688# 0.196132f
C136 source.n8 a_n2204_n2688# 1.64189f
C137 source.n9 a_n2204_n2688# 0.399509f
C138 source.t7 a_n2204_n2688# 0.196132f
C139 source.t0 a_n2204_n2688# 0.196132f
C140 source.n10 a_n2204_n2688# 1.64189f
C141 source.n11 a_n2204_n2688# 0.399509f
C142 source.t10 a_n2204_n2688# 0.196132f
C143 source.t3 a_n2204_n2688# 0.196132f
C144 source.n12 a_n2204_n2688# 1.64189f
C145 source.n13 a_n2204_n2688# 1.63519f
C146 source.t18 a_n2204_n2688# 0.196132f
C147 source.t23 a_n2204_n2688# 0.196132f
C148 source.n14 a_n2204_n2688# 1.64189f
C149 source.n15 a_n2204_n2688# 1.6352f
C150 source.t22 a_n2204_n2688# 0.196132f
C151 source.t13 a_n2204_n2688# 0.196132f
C152 source.n16 a_n2204_n2688# 1.64189f
C153 source.n17 a_n2204_n2688# 0.399514f
C154 source.t15 a_n2204_n2688# 0.196132f
C155 source.t25 a_n2204_n2688# 0.196132f
C156 source.n18 a_n2204_n2688# 1.64189f
C157 source.n19 a_n2204_n2688# 0.399514f
C158 source.t14 a_n2204_n2688# 2.09145f
C159 source.n20 a_n2204_n2688# 0.490985f
C160 source.t9 a_n2204_n2688# 0.196132f
C161 source.t12 a_n2204_n2688# 0.196132f
C162 source.n21 a_n2204_n2688# 1.64189f
C163 source.n22 a_n2204_n2688# 0.405642f
C164 source.t4 a_n2204_n2688# 0.196132f
C165 source.t27 a_n2204_n2688# 0.196132f
C166 source.n23 a_n2204_n2688# 1.64189f
C167 source.n24 a_n2204_n2688# 0.399514f
C168 source.t5 a_n2204_n2688# 0.196132f
C169 source.t6 a_n2204_n2688# 0.196132f
C170 source.n25 a_n2204_n2688# 1.64189f
C171 source.n26 a_n2204_n2688# 0.399514f
C172 source.t8 a_n2204_n2688# 2.09145f
C173 source.n27 a_n2204_n2688# 0.62925f
C174 source.n28 a_n2204_n2688# 1.44789f
C175 plus.n0 a_n2204_n2688# 0.044229f
C176 plus.t0 a_n2204_n2688# 0.684957f
C177 plus.t1 a_n2204_n2688# 0.684957f
C178 plus.n1 a_n2204_n2688# 0.044229f
C179 plus.t3 a_n2204_n2688# 0.684957f
C180 plus.n2 a_n2204_n2688# 0.290465f
C181 plus.n3 a_n2204_n2688# 0.059019f
C182 plus.t6 a_n2204_n2688# 0.684957f
C183 plus.t7 a_n2204_n2688# 0.684957f
C184 plus.t8 a_n2204_n2688# 0.684957f
C185 plus.n4 a_n2204_n2688# 0.297307f
C186 plus.t9 a_n2204_n2688# 0.700251f
C187 plus.n5 a_n2204_n2688# 0.277608f
C188 plus.n6 a_n2204_n2688# 0.180947f
C189 plus.n7 a_n2204_n2688# 0.010037f
C190 plus.n8 a_n2204_n2688# 0.290465f
C191 plus.n9 a_n2204_n2688# 0.299956f
C192 plus.n10 a_n2204_n2688# 0.058881f
C193 plus.n11 a_n2204_n2688# 0.059019f
C194 plus.n12 a_n2204_n2688# 0.044229f
C195 plus.n13 a_n2204_n2688# 0.010037f
C196 plus.n14 a_n2204_n2688# 0.291828f
C197 plus.n15 a_n2204_n2688# 0.010037f
C198 plus.n16 a_n2204_n2688# 0.287465f
C199 plus.n17 a_n2204_n2688# 0.442426f
C200 plus.n18 a_n2204_n2688# 0.044229f
C201 plus.t5 a_n2204_n2688# 0.684957f
C202 plus.n19 a_n2204_n2688# 0.044229f
C203 plus.t13 a_n2204_n2688# 0.684957f
C204 plus.t12 a_n2204_n2688# 0.684957f
C205 plus.n20 a_n2204_n2688# 0.290465f
C206 plus.n21 a_n2204_n2688# 0.059019f
C207 plus.t11 a_n2204_n2688# 0.684957f
C208 plus.t4 a_n2204_n2688# 0.684957f
C209 plus.t2 a_n2204_n2688# 0.684957f
C210 plus.n22 a_n2204_n2688# 0.297307f
C211 plus.t10 a_n2204_n2688# 0.700251f
C212 plus.n23 a_n2204_n2688# 0.277608f
C213 plus.n24 a_n2204_n2688# 0.180947f
C214 plus.n25 a_n2204_n2688# 0.010037f
C215 plus.n26 a_n2204_n2688# 0.290465f
C216 plus.n27 a_n2204_n2688# 0.299956f
C217 plus.n28 a_n2204_n2688# 0.058881f
C218 plus.n29 a_n2204_n2688# 0.059019f
C219 plus.n30 a_n2204_n2688# 0.044229f
C220 plus.n31 a_n2204_n2688# 0.010037f
C221 plus.n32 a_n2204_n2688# 0.291828f
C222 plus.n33 a_n2204_n2688# 0.010037f
C223 plus.n34 a_n2204_n2688# 0.287465f
C224 plus.n35 a_n2204_n2688# 1.31468f
.ends

