* NGSPICE file created from diffpair483.ext - technology: sky130A

.subckt diffpair483 minus drain_right drain_left source plus
X0 a_n1366_n3888# a_n1366_n3888# a_n1366_n3888# a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=57 ps=247.6 w=15 l=0.15
X1 drain_right.t7 minus.t0 source.t4 a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X2 source.t11 minus.t1 drain_right.t6 a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X3 drain_left.t7 plus.t0 source.t1 a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X4 a_n1366_n3888# a_n1366_n3888# a_n1366_n3888# a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X5 source.t8 minus.t2 drain_right.t5 a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X6 drain_right.t4 minus.t3 source.t7 a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X7 a_n1366_n3888# a_n1366_n3888# a_n1366_n3888# a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X8 source.t12 plus.t1 drain_left.t6 a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X9 source.t9 minus.t4 drain_right.t3 a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X10 a_n1366_n3888# a_n1366_n3888# a_n1366_n3888# a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X11 source.t13 plus.t2 drain_left.t5 a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X12 drain_right.t2 minus.t5 source.t10 a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X13 drain_left.t4 plus.t3 source.t14 a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X14 drain_left.t3 plus.t4 source.t15 a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X15 drain_right.t1 minus.t6 source.t5 a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X16 source.t0 plus.t5 drain_left.t2 a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X17 drain_left.t1 plus.t6 source.t3 a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X18 source.t2 plus.t7 drain_left.t0 a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X19 source.t6 minus.t7 drain_right.t0 a_n1366_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
R0 minus.n5 minus.t4 2688.25
R1 minus.n1 minus.t3 2688.25
R2 minus.n12 minus.t0 2688.25
R3 minus.n8 minus.t1 2688.25
R4 minus.n4 minus.t5 2618.87
R5 minus.n2 minus.t2 2618.87
R6 minus.n11 minus.t7 2618.87
R7 minus.n9 minus.t6 2618.87
R8 minus.n1 minus.n0 161.489
R9 minus.n8 minus.n7 161.489
R10 minus.n6 minus.n5 161.3
R11 minus.n3 minus.n0 161.3
R12 minus.n13 minus.n12 161.3
R13 minus.n10 minus.n7 161.3
R14 minus.n4 minus.n3 47.4702
R15 minus.n3 minus.n2 47.4702
R16 minus.n10 minus.n9 47.4702
R17 minus.n11 minus.n10 47.4702
R18 minus.n14 minus.n6 36.6482
R19 minus.n5 minus.n4 25.5611
R20 minus.n2 minus.n1 25.5611
R21 minus.n9 minus.n8 25.5611
R22 minus.n12 minus.n11 25.5611
R23 minus.n14 minus.n13 6.58005
R24 minus.n6 minus.n0 0.189894
R25 minus.n13 minus.n7 0.189894
R26 minus minus.n14 0.188
R27 source.n3 source.t13 46.201
R28 source.n4 source.t7 46.201
R29 source.n7 source.t9 46.201
R30 source.n15 source.t4 46.2008
R31 source.n12 source.t11 46.2008
R32 source.n11 source.t14 46.2008
R33 source.n8 source.t12 46.2008
R34 source.n0 source.t15 46.2008
R35 source.n2 source.n1 44.201
R36 source.n6 source.n5 44.201
R37 source.n14 source.n13 44.2008
R38 source.n10 source.n9 44.2008
R39 source.n8 source.n7 24.1208
R40 source.n16 source.n0 18.5777
R41 source.n16 source.n15 5.5436
R42 source.n13 source.t5 2.0005
R43 source.n13 source.t6 2.0005
R44 source.n9 source.t1 2.0005
R45 source.n9 source.t2 2.0005
R46 source.n1 source.t3 2.0005
R47 source.n1 source.t0 2.0005
R48 source.n5 source.t10 2.0005
R49 source.n5 source.t8 2.0005
R50 source.n7 source.n6 0.560845
R51 source.n6 source.n4 0.560845
R52 source.n3 source.n2 0.560845
R53 source.n2 source.n0 0.560845
R54 source.n10 source.n8 0.560845
R55 source.n11 source.n10 0.560845
R56 source.n14 source.n12 0.560845
R57 source.n15 source.n14 0.560845
R58 source.n4 source.n3 0.470328
R59 source.n12 source.n11 0.470328
R60 source source.n16 0.188
R61 drain_right.n5 drain_right.n3 61.44
R62 drain_right.n2 drain_right.n1 61.1044
R63 drain_right.n2 drain_right.n0 61.1044
R64 drain_right.n5 drain_right.n4 60.8798
R65 drain_right drain_right.n2 31.0478
R66 drain_right drain_right.n5 6.21356
R67 drain_right.n1 drain_right.t0 2.0005
R68 drain_right.n1 drain_right.t7 2.0005
R69 drain_right.n0 drain_right.t6 2.0005
R70 drain_right.n0 drain_right.t1 2.0005
R71 drain_right.n3 drain_right.t5 2.0005
R72 drain_right.n3 drain_right.t4 2.0005
R73 drain_right.n4 drain_right.t3 2.0005
R74 drain_right.n4 drain_right.t2 2.0005
R75 plus.n1 plus.t2 2688.25
R76 plus.n5 plus.t4 2688.25
R77 plus.n8 plus.t3 2688.25
R78 plus.n12 plus.t1 2688.25
R79 plus.n2 plus.t6 2618.87
R80 plus.n4 plus.t5 2618.87
R81 plus.n9 plus.t7 2618.87
R82 plus.n11 plus.t0 2618.87
R83 plus.n1 plus.n0 161.489
R84 plus.n8 plus.n7 161.489
R85 plus.n3 plus.n0 161.3
R86 plus.n6 plus.n5 161.3
R87 plus.n10 plus.n7 161.3
R88 plus.n13 plus.n12 161.3
R89 plus.n3 plus.n2 47.4702
R90 plus.n4 plus.n3 47.4702
R91 plus.n11 plus.n10 47.4702
R92 plus.n10 plus.n9 47.4702
R93 plus plus.n13 29.393
R94 plus.n2 plus.n1 25.5611
R95 plus.n5 plus.n4 25.5611
R96 plus.n12 plus.n11 25.5611
R97 plus.n9 plus.n8 25.5611
R98 plus plus.n6 13.3603
R99 plus.n6 plus.n0 0.189894
R100 plus.n13 plus.n7 0.189894
R101 drain_left.n5 drain_left.n3 61.4402
R102 drain_left.n2 drain_left.n1 61.1044
R103 drain_left.n2 drain_left.n0 61.1044
R104 drain_left.n5 drain_left.n4 60.8796
R105 drain_left drain_left.n2 31.601
R106 drain_left drain_left.n5 6.21356
R107 drain_left.n1 drain_left.t0 2.0005
R108 drain_left.n1 drain_left.t4 2.0005
R109 drain_left.n0 drain_left.t6 2.0005
R110 drain_left.n0 drain_left.t7 2.0005
R111 drain_left.n4 drain_left.t2 2.0005
R112 drain_left.n4 drain_left.t3 2.0005
R113 drain_left.n3 drain_left.t5 2.0005
R114 drain_left.n3 drain_left.t1 2.0005
C0 source plus 1.94565f
C1 source minus 1.93161f
C2 minus plus 5.39063f
C3 drain_right drain_left 0.640281f
C4 drain_right source 20.662802f
C5 drain_right plus 0.282599f
C6 drain_right minus 2.63358f
C7 source drain_left 20.6635f
C8 drain_left plus 2.76298f
C9 drain_left minus 0.170499f
C10 drain_right a_n1366_n3888# 5.91171f
C11 drain_left a_n1366_n3888# 6.11775f
C12 source a_n1366_n3888# 10.194994f
C13 minus a_n1366_n3888# 5.187947f
C14 plus a_n1366_n3888# 7.1559f
C15 drain_left.t6 a_n1366_n3888# 0.506978f
C16 drain_left.t7 a_n1366_n3888# 0.506978f
C17 drain_left.n0 a_n1366_n3888# 3.37036f
C18 drain_left.t0 a_n1366_n3888# 0.506978f
C19 drain_left.t4 a_n1366_n3888# 0.506978f
C20 drain_left.n1 a_n1366_n3888# 3.37036f
C21 drain_left.n2 a_n1366_n3888# 2.07552f
C22 drain_left.t5 a_n1366_n3888# 0.506978f
C23 drain_left.t1 a_n1366_n3888# 0.506978f
C24 drain_left.n3 a_n1366_n3888# 3.37233f
C25 drain_left.t2 a_n1366_n3888# 0.506978f
C26 drain_left.t3 a_n1366_n3888# 0.506978f
C27 drain_left.n4 a_n1366_n3888# 3.36918f
C28 drain_left.n5 a_n1366_n3888# 0.910262f
C29 plus.n0 a_n1366_n3888# 0.118203f
C30 plus.t5 a_n1366_n3888# 0.31681f
C31 plus.t6 a_n1366_n3888# 0.31681f
C32 plus.t2 a_n1366_n3888# 0.320248f
C33 plus.n1 a_n1366_n3888# 0.151042f
C34 plus.n2 a_n1366_n3888# 0.129382f
C35 plus.n3 a_n1366_n3888# 0.021173f
C36 plus.n4 a_n1366_n3888# 0.129382f
C37 plus.t4 a_n1366_n3888# 0.320248f
C38 plus.n5 a_n1366_n3888# 0.150962f
C39 plus.n6 a_n1366_n3888# 0.640102f
C40 plus.n7 a_n1366_n3888# 0.118203f
C41 plus.t1 a_n1366_n3888# 0.320248f
C42 plus.t0 a_n1366_n3888# 0.31681f
C43 plus.t7 a_n1366_n3888# 0.31681f
C44 plus.t3 a_n1366_n3888# 0.320248f
C45 plus.n8 a_n1366_n3888# 0.151042f
C46 plus.n9 a_n1366_n3888# 0.129382f
C47 plus.n10 a_n1366_n3888# 0.021173f
C48 plus.n11 a_n1366_n3888# 0.129382f
C49 plus.n12 a_n1366_n3888# 0.150962f
C50 plus.n13 a_n1366_n3888# 1.47654f
C51 drain_right.t6 a_n1366_n3888# 0.505037f
C52 drain_right.t1 a_n1366_n3888# 0.505037f
C53 drain_right.n0 a_n1366_n3888# 3.35745f
C54 drain_right.t0 a_n1366_n3888# 0.505037f
C55 drain_right.t7 a_n1366_n3888# 0.505037f
C56 drain_right.n1 a_n1366_n3888# 3.35745f
C57 drain_right.n2 a_n1366_n3888# 2.00854f
C58 drain_right.t5 a_n1366_n3888# 0.505037f
C59 drain_right.t4 a_n1366_n3888# 0.505037f
C60 drain_right.n3 a_n1366_n3888# 3.35941f
C61 drain_right.t3 a_n1366_n3888# 0.505037f
C62 drain_right.t2 a_n1366_n3888# 0.505037f
C63 drain_right.n4 a_n1366_n3888# 3.35629f
C64 drain_right.n5 a_n1366_n3888# 0.906776f
C65 source.t15 a_n1366_n3888# 2.68396f
C66 source.n0 a_n1366_n3888# 1.19483f
C67 source.t3 a_n1366_n3888# 0.337075f
C68 source.t0 a_n1366_n3888# 0.337075f
C69 source.n1 a_n1366_n3888# 2.18342f
C70 source.n2 a_n1366_n3888# 0.252645f
C71 source.t13 a_n1366_n3888# 2.68396f
C72 source.n3 a_n1366_n3888# 0.353363f
C73 source.t7 a_n1366_n3888# 2.68396f
C74 source.n4 a_n1366_n3888# 0.353363f
C75 source.t10 a_n1366_n3888# 0.337075f
C76 source.t8 a_n1366_n3888# 0.337075f
C77 source.n5 a_n1366_n3888# 2.18342f
C78 source.n6 a_n1366_n3888# 0.252645f
C79 source.t9 a_n1366_n3888# 2.68396f
C80 source.n7 a_n1366_n3888# 1.50727f
C81 source.t12 a_n1366_n3888# 2.68396f
C82 source.n8 a_n1366_n3888# 1.50728f
C83 source.t1 a_n1366_n3888# 0.337075f
C84 source.t2 a_n1366_n3888# 0.337075f
C85 source.n9 a_n1366_n3888# 2.18341f
C86 source.n10 a_n1366_n3888# 0.252647f
C87 source.t14 a_n1366_n3888# 2.68396f
C88 source.n11 a_n1366_n3888# 0.353366f
C89 source.t11 a_n1366_n3888# 2.68396f
C90 source.n12 a_n1366_n3888# 0.353366f
C91 source.t5 a_n1366_n3888# 0.337075f
C92 source.t6 a_n1366_n3888# 0.337075f
C93 source.n13 a_n1366_n3888# 2.18341f
C94 source.n14 a_n1366_n3888# 0.252647f
C95 source.t4 a_n1366_n3888# 2.68396f
C96 source.n15 a_n1366_n3888# 0.460146f
C97 source.n16 a_n1366_n3888# 1.37292f
C98 minus.n0 a_n1366_n3888# 0.113918f
C99 minus.t4 a_n1366_n3888# 0.308638f
C100 minus.t5 a_n1366_n3888# 0.305325f
C101 minus.t2 a_n1366_n3888# 0.305325f
C102 minus.t3 a_n1366_n3888# 0.308638f
C103 minus.n1 a_n1366_n3888# 0.145567f
C104 minus.n2 a_n1366_n3888# 0.124691f
C105 minus.n3 a_n1366_n3888# 0.020405f
C106 minus.n4 a_n1366_n3888# 0.124691f
C107 minus.n5 a_n1366_n3888# 0.145489f
C108 minus.n6 a_n1366_n3888# 1.73627f
C109 minus.n7 a_n1366_n3888# 0.113918f
C110 minus.t7 a_n1366_n3888# 0.305325f
C111 minus.t6 a_n1366_n3888# 0.305325f
C112 minus.t1 a_n1366_n3888# 0.308638f
C113 minus.n8 a_n1366_n3888# 0.145567f
C114 minus.n9 a_n1366_n3888# 0.124691f
C115 minus.n10 a_n1366_n3888# 0.020405f
C116 minus.n11 a_n1366_n3888# 0.124691f
C117 minus.t0 a_n1366_n3888# 0.308638f
C118 minus.n12 a_n1366_n3888# 0.145489f
C119 minus.n13 a_n1366_n3888# 0.323508f
C120 minus.n14 a_n1366_n3888# 2.10326f
.ends

