* NGSPICE file created from diffpair556.ext - technology: sky130A

.subckt diffpair556 minus drain_right drain_left source plus
X0 drain_left.t13 plus.t0 source.t26 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X1 drain_right.t13 minus.t0 source.t6 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X2 drain_right.t12 minus.t1 source.t1 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X3 source.t23 plus.t1 drain_left.t12 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X4 a_n2524_n3888# a_n2524_n3888# a_n2524_n3888# a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.8
X5 a_n2524_n3888# a_n2524_n3888# a_n2524_n3888# a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X6 a_n2524_n3888# a_n2524_n3888# a_n2524_n3888# a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X7 a_n2524_n3888# a_n2524_n3888# a_n2524_n3888# a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.8
X8 source.t9 minus.t2 drain_right.t11 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X9 drain_right.t10 minus.t3 source.t11 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X10 source.t10 minus.t4 drain_right.t9 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X11 source.t14 plus.t2 drain_left.t11 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X12 source.t2 minus.t5 drain_right.t8 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X13 drain_right.t7 minus.t6 source.t7 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X14 source.t25 plus.t3 drain_left.t10 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X15 drain_right.t6 minus.t7 source.t8 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X16 source.t0 minus.t8 drain_right.t5 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X17 source.t3 minus.t9 drain_right.t4 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X18 drain_left.t9 plus.t4 source.t19 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X19 source.t27 minus.t10 drain_right.t3 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X20 drain_right.t2 minus.t11 source.t5 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X21 drain_left.t8 plus.t5 source.t20 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X22 source.t21 plus.t6 drain_left.t7 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X23 source.t22 plus.t7 drain_left.t6 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X24 drain_left.t5 plus.t8 source.t18 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X25 drain_left.t4 plus.t9 source.t16 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X26 drain_left.t3 plus.t10 source.t15 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X27 source.t24 plus.t11 drain_left.t2 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X28 drain_left.t1 plus.t12 source.t13 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
X29 drain_right.t1 minus.t12 source.t4 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.8
X30 drain_left.t0 plus.t13 source.t17 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.8
X31 drain_right.t0 minus.t13 source.t12 a_n2524_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.8
R0 plus.n5 plus.t13 524.826
R1 plus.n23 plus.t0 524.826
R2 plus.n16 plus.t5 500.979
R3 plus.n14 plus.t6 500.979
R4 plus.n2 plus.t10 500.979
R5 plus.n9 plus.t7 500.979
R6 plus.n8 plus.t8 500.979
R7 plus.n4 plus.t11 500.979
R8 plus.n34 plus.t4 500.979
R9 plus.n32 plus.t1 500.979
R10 plus.n20 plus.t9 500.979
R11 plus.n27 plus.t2 500.979
R12 plus.n26 plus.t12 500.979
R13 plus.n22 plus.t3 500.979
R14 plus.n7 plus.n6 161.3
R15 plus.n13 plus.n12 161.3
R16 plus.n14 plus.n1 161.3
R17 plus.n15 plus.n0 161.3
R18 plus.n17 plus.n16 161.3
R19 plus.n25 plus.n24 161.3
R20 plus.n31 plus.n30 161.3
R21 plus.n32 plus.n19 161.3
R22 plus.n33 plus.n18 161.3
R23 plus.n35 plus.n34 161.3
R24 plus.n8 plus.n3 80.6037
R25 plus.n10 plus.n9 80.6037
R26 plus.n11 plus.n2 80.6037
R27 plus.n26 plus.n21 80.6037
R28 plus.n28 plus.n27 80.6037
R29 plus.n29 plus.n20 80.6037
R30 plus.n9 plus.n2 48.2005
R31 plus.n9 plus.n8 48.2005
R32 plus.n27 plus.n20 48.2005
R33 plus.n27 plus.n26 48.2005
R34 plus.n24 plus.n23 44.9119
R35 plus.n6 plus.n5 44.9119
R36 plus.n16 plus.n15 35.055
R37 plus.n34 plus.n33 35.055
R38 plus plus.n35 33.9252
R39 plus.n13 plus.n2 32.1338
R40 plus.n8 plus.n7 32.1338
R41 plus.n31 plus.n20 32.1338
R42 plus.n26 plus.n25 32.1338
R43 plus.n23 plus.n22 17.739
R44 plus.n5 plus.n4 17.739
R45 plus.n14 plus.n13 16.0672
R46 plus.n7 plus.n4 16.0672
R47 plus.n32 plus.n31 16.0672
R48 plus.n25 plus.n22 16.0672
R49 plus plus.n17 13.5062
R50 plus.n15 plus.n14 13.146
R51 plus.n33 plus.n32 13.146
R52 plus.n10 plus.n3 0.380177
R53 plus.n11 plus.n10 0.380177
R54 plus.n29 plus.n28 0.380177
R55 plus.n28 plus.n21 0.380177
R56 plus.n6 plus.n3 0.285035
R57 plus.n12 plus.n11 0.285035
R58 plus.n30 plus.n29 0.285035
R59 plus.n24 plus.n21 0.285035
R60 plus.n12 plus.n1 0.189894
R61 plus.n1 plus.n0 0.189894
R62 plus.n17 plus.n0 0.189894
R63 plus.n35 plus.n18 0.189894
R64 plus.n19 plus.n18 0.189894
R65 plus.n30 plus.n19 0.189894
R66 source.n7 source.t8 45.521
R67 source.n27 source.t4 45.5208
R68 source.n20 source.t26 45.5208
R69 source.n0 source.t20 45.5208
R70 source.n2 source.n1 44.201
R71 source.n4 source.n3 44.201
R72 source.n6 source.n5 44.201
R73 source.n9 source.n8 44.201
R74 source.n11 source.n10 44.201
R75 source.n13 source.n12 44.201
R76 source.n26 source.n25 44.2008
R77 source.n24 source.n23 44.2008
R78 source.n22 source.n21 44.2008
R79 source.n19 source.n18 44.2008
R80 source.n17 source.n16 44.2008
R81 source.n15 source.n14 44.2008
R82 source.n15 source.n13 25.5087
R83 source.n28 source.n0 18.7846
R84 source.n28 source.n27 5.7505
R85 source.n25 source.t6 1.3205
R86 source.n25 source.t9 1.3205
R87 source.n23 source.t12 1.3205
R88 source.n23 source.t10 1.3205
R89 source.n21 source.t1 1.3205
R90 source.n21 source.t3 1.3205
R91 source.n18 source.t13 1.3205
R92 source.n18 source.t25 1.3205
R93 source.n16 source.t16 1.3205
R94 source.n16 source.t14 1.3205
R95 source.n14 source.t19 1.3205
R96 source.n14 source.t23 1.3205
R97 source.n1 source.t15 1.3205
R98 source.n1 source.t21 1.3205
R99 source.n3 source.t18 1.3205
R100 source.n3 source.t22 1.3205
R101 source.n5 source.t17 1.3205
R102 source.n5 source.t24 1.3205
R103 source.n8 source.t11 1.3205
R104 source.n8 source.t2 1.3205
R105 source.n10 source.t5 1.3205
R106 source.n10 source.t27 1.3205
R107 source.n12 source.t7 1.3205
R108 source.n12 source.t0 1.3205
R109 source.n13 source.n11 0.974638
R110 source.n11 source.n9 0.974638
R111 source.n9 source.n7 0.974638
R112 source.n6 source.n4 0.974638
R113 source.n4 source.n2 0.974638
R114 source.n2 source.n0 0.974638
R115 source.n17 source.n15 0.974638
R116 source.n19 source.n17 0.974638
R117 source.n20 source.n19 0.974638
R118 source.n24 source.n22 0.974638
R119 source.n26 source.n24 0.974638
R120 source.n27 source.n26 0.974638
R121 source.n7 source.n6 0.957397
R122 source.n22 source.n20 0.957397
R123 source source.n28 0.188
R124 drain_left.n7 drain_left.t0 63.1739
R125 drain_left.n1 drain_left.t9 63.1737
R126 drain_left.n4 drain_left.n2 61.8537
R127 drain_left.n9 drain_left.n8 60.8798
R128 drain_left.n7 drain_left.n6 60.8798
R129 drain_left.n11 drain_left.n10 60.8796
R130 drain_left.n4 drain_left.n3 60.8796
R131 drain_left.n1 drain_left.n0 60.8796
R132 drain_left drain_left.n5 35.2411
R133 drain_left drain_left.n11 6.62735
R134 drain_left.n2 drain_left.t10 1.3205
R135 drain_left.n2 drain_left.t13 1.3205
R136 drain_left.n3 drain_left.t11 1.3205
R137 drain_left.n3 drain_left.t1 1.3205
R138 drain_left.n0 drain_left.t12 1.3205
R139 drain_left.n0 drain_left.t4 1.3205
R140 drain_left.n10 drain_left.t7 1.3205
R141 drain_left.n10 drain_left.t8 1.3205
R142 drain_left.n8 drain_left.t6 1.3205
R143 drain_left.n8 drain_left.t3 1.3205
R144 drain_left.n6 drain_left.t2 1.3205
R145 drain_left.n6 drain_left.t5 1.3205
R146 drain_left.n9 drain_left.n7 0.974638
R147 drain_left.n11 drain_left.n9 0.974638
R148 drain_left.n5 drain_left.n1 0.675757
R149 drain_left.n5 drain_left.n4 0.188688
R150 minus.n5 minus.t7 524.826
R151 minus.n23 minus.t1 524.826
R152 minus.n4 minus.t5 500.979
R153 minus.n8 minus.t3 500.979
R154 minus.n9 minus.t10 500.979
R155 minus.n10 minus.t11 500.979
R156 minus.n14 minus.t8 500.979
R157 minus.n16 minus.t6 500.979
R158 minus.n22 minus.t9 500.979
R159 minus.n26 minus.t13 500.979
R160 minus.n27 minus.t4 500.979
R161 minus.n28 minus.t0 500.979
R162 minus.n32 minus.t2 500.979
R163 minus.n34 minus.t12 500.979
R164 minus.n17 minus.n16 161.3
R165 minus.n15 minus.n0 161.3
R166 minus.n14 minus.n13 161.3
R167 minus.n12 minus.n1 161.3
R168 minus.n6 minus.n3 161.3
R169 minus.n35 minus.n34 161.3
R170 minus.n33 minus.n18 161.3
R171 minus.n32 minus.n31 161.3
R172 minus.n30 minus.n19 161.3
R173 minus.n24 minus.n21 161.3
R174 minus.n11 minus.n10 80.6037
R175 minus.n9 minus.n2 80.6037
R176 minus.n8 minus.n7 80.6037
R177 minus.n29 minus.n28 80.6037
R178 minus.n27 minus.n20 80.6037
R179 minus.n26 minus.n25 80.6037
R180 minus.n9 minus.n8 48.2005
R181 minus.n10 minus.n9 48.2005
R182 minus.n27 minus.n26 48.2005
R183 minus.n28 minus.n27 48.2005
R184 minus.n6 minus.n5 44.9119
R185 minus.n24 minus.n23 44.9119
R186 minus.n36 minus.n17 41.1804
R187 minus.n16 minus.n15 35.055
R188 minus.n34 minus.n33 35.055
R189 minus.n8 minus.n3 32.1338
R190 minus.n10 minus.n1 32.1338
R191 minus.n26 minus.n21 32.1338
R192 minus.n28 minus.n19 32.1338
R193 minus.n5 minus.n4 17.739
R194 minus.n23 minus.n22 17.739
R195 minus.n4 minus.n3 16.0672
R196 minus.n14 minus.n1 16.0672
R197 minus.n22 minus.n21 16.0672
R198 minus.n32 minus.n19 16.0672
R199 minus.n15 minus.n14 13.146
R200 minus.n33 minus.n32 13.146
R201 minus.n36 minus.n35 6.72588
R202 minus.n11 minus.n2 0.380177
R203 minus.n7 minus.n2 0.380177
R204 minus.n25 minus.n20 0.380177
R205 minus.n29 minus.n20 0.380177
R206 minus.n12 minus.n11 0.285035
R207 minus.n7 minus.n6 0.285035
R208 minus.n25 minus.n24 0.285035
R209 minus.n30 minus.n29 0.285035
R210 minus.n17 minus.n0 0.189894
R211 minus.n13 minus.n0 0.189894
R212 minus.n13 minus.n12 0.189894
R213 minus.n31 minus.n30 0.189894
R214 minus.n31 minus.n18 0.189894
R215 minus.n35 minus.n18 0.189894
R216 minus minus.n36 0.188
R217 drain_right.n1 drain_right.t12 63.1737
R218 drain_right.n11 drain_right.t7 62.1998
R219 drain_right.n8 drain_right.n6 61.8538
R220 drain_right.n4 drain_right.n2 61.8537
R221 drain_right.n8 drain_right.n7 60.8798
R222 drain_right.n10 drain_right.n9 60.8798
R223 drain_right.n4 drain_right.n3 60.8796
R224 drain_right.n1 drain_right.n0 60.8796
R225 drain_right drain_right.n5 34.6879
R226 drain_right drain_right.n11 6.14028
R227 drain_right.n2 drain_right.t11 1.3205
R228 drain_right.n2 drain_right.t1 1.3205
R229 drain_right.n3 drain_right.t9 1.3205
R230 drain_right.n3 drain_right.t13 1.3205
R231 drain_right.n0 drain_right.t4 1.3205
R232 drain_right.n0 drain_right.t0 1.3205
R233 drain_right.n6 drain_right.t8 1.3205
R234 drain_right.n6 drain_right.t6 1.3205
R235 drain_right.n7 drain_right.t3 1.3205
R236 drain_right.n7 drain_right.t10 1.3205
R237 drain_right.n9 drain_right.t5 1.3205
R238 drain_right.n9 drain_right.t2 1.3205
R239 drain_right.n11 drain_right.n10 0.974638
R240 drain_right.n10 drain_right.n8 0.974638
R241 drain_right.n5 drain_right.n1 0.675757
R242 drain_right.n5 drain_right.n4 0.188688
C0 drain_right minus 12.016701f
C1 source drain_right 21.0801f
C2 drain_left drain_right 1.31793f
C3 source minus 11.929299f
C4 drain_left minus 0.173289f
C5 source drain_left 21.087198f
C6 drain_right plus 0.408742f
C7 plus minus 6.8422f
C8 source plus 11.943901f
C9 drain_left plus 12.2637f
C10 drain_right a_n2524_n3888# 8.51489f
C11 drain_left a_n2524_n3888# 8.8912f
C12 source a_n2524_n3888# 7.908649f
C13 minus a_n2524_n3888# 10.236322f
C14 plus a_n2524_n3888# 12.0517f
C15 drain_right.t12 a_n2524_n3888# 3.33745f
C16 drain_right.t4 a_n2524_n3888# 0.288797f
C17 drain_right.t0 a_n2524_n3888# 0.288797f
C18 drain_right.n0 a_n2524_n3888# 2.61038f
C19 drain_right.n1 a_n2524_n3888# 0.676282f
C20 drain_right.t11 a_n2524_n3888# 0.288797f
C21 drain_right.t1 a_n2524_n3888# 0.288797f
C22 drain_right.n2 a_n2524_n3888# 2.61609f
C23 drain_right.t9 a_n2524_n3888# 0.288797f
C24 drain_right.t13 a_n2524_n3888# 0.288797f
C25 drain_right.n3 a_n2524_n3888# 2.61038f
C26 drain_right.n4 a_n2524_n3888# 0.65042f
C27 drain_right.n5 a_n2524_n3888# 1.51543f
C28 drain_right.t8 a_n2524_n3888# 0.288797f
C29 drain_right.t6 a_n2524_n3888# 0.288797f
C30 drain_right.n6 a_n2524_n3888# 2.61608f
C31 drain_right.t3 a_n2524_n3888# 0.288797f
C32 drain_right.t10 a_n2524_n3888# 0.288797f
C33 drain_right.n7 a_n2524_n3888# 2.61039f
C34 drain_right.n8 a_n2524_n3888# 0.709125f
C35 drain_right.t5 a_n2524_n3888# 0.288797f
C36 drain_right.t2 a_n2524_n3888# 0.288797f
C37 drain_right.n9 a_n2524_n3888# 2.61039f
C38 drain_right.n10 a_n2524_n3888# 0.352504f
C39 drain_right.t7 a_n2524_n3888# 3.33203f
C40 drain_right.n11 a_n2524_n3888# 0.580847f
C41 minus.n0 a_n2524_n3888# 0.038714f
C42 minus.n1 a_n2524_n3888# 0.008785f
C43 minus.t8 a_n2524_n3888# 1.32017f
C44 minus.n2 a_n2524_n3888# 0.077428f
C45 minus.n3 a_n2524_n3888# 0.008785f
C46 minus.t3 a_n2524_n3888# 1.32017f
C47 minus.t7 a_n2524_n3888# 1.34327f
C48 minus.t5 a_n2524_n3888# 1.32017f
C49 minus.n4 a_n2524_n3888# 0.510712f
C50 minus.n5 a_n2524_n3888# 0.488608f
C51 minus.n6 a_n2524_n3888# 0.1808f
C52 minus.n7 a_n2524_n3888# 0.064483f
C53 minus.n8 a_n2524_n3888# 0.515179f
C54 minus.t10 a_n2524_n3888# 1.32017f
C55 minus.n9 a_n2524_n3888# 0.517805f
C56 minus.t11 a_n2524_n3888# 1.32017f
C57 minus.n10 a_n2524_n3888# 0.515179f
C58 minus.n11 a_n2524_n3888# 0.064483f
C59 minus.n12 a_n2524_n3888# 0.051659f
C60 minus.n13 a_n2524_n3888# 0.038714f
C61 minus.n14 a_n2524_n3888# 0.505917f
C62 minus.n15 a_n2524_n3888# 0.008785f
C63 minus.t6 a_n2524_n3888# 1.32017f
C64 minus.n16 a_n2524_n3888# 0.506872f
C65 minus.n17 a_n2524_n3888# 1.67122f
C66 minus.n18 a_n2524_n3888# 0.038714f
C67 minus.n19 a_n2524_n3888# 0.008785f
C68 minus.n20 a_n2524_n3888# 0.077428f
C69 minus.n21 a_n2524_n3888# 0.008785f
C70 minus.t1 a_n2524_n3888# 1.34327f
C71 minus.t9 a_n2524_n3888# 1.32017f
C72 minus.n22 a_n2524_n3888# 0.510712f
C73 minus.n23 a_n2524_n3888# 0.488608f
C74 minus.n24 a_n2524_n3888# 0.1808f
C75 minus.n25 a_n2524_n3888# 0.064483f
C76 minus.t13 a_n2524_n3888# 1.32017f
C77 minus.n26 a_n2524_n3888# 0.515179f
C78 minus.t4 a_n2524_n3888# 1.32017f
C79 minus.n27 a_n2524_n3888# 0.517805f
C80 minus.t0 a_n2524_n3888# 1.32017f
C81 minus.n28 a_n2524_n3888# 0.515179f
C82 minus.n29 a_n2524_n3888# 0.064483f
C83 minus.n30 a_n2524_n3888# 0.051659f
C84 minus.n31 a_n2524_n3888# 0.038714f
C85 minus.t2 a_n2524_n3888# 1.32017f
C86 minus.n32 a_n2524_n3888# 0.505917f
C87 minus.n33 a_n2524_n3888# 0.008785f
C88 minus.t12 a_n2524_n3888# 1.32017f
C89 minus.n34 a_n2524_n3888# 0.506872f
C90 minus.n35 a_n2524_n3888# 0.273491f
C91 minus.n36 a_n2524_n3888# 1.99548f
C92 drain_left.t9 a_n2524_n3888# 3.35803f
C93 drain_left.t12 a_n2524_n3888# 0.290577f
C94 drain_left.t4 a_n2524_n3888# 0.290577f
C95 drain_left.n0 a_n2524_n3888# 2.62648f
C96 drain_left.n1 a_n2524_n3888# 0.680453f
C97 drain_left.t10 a_n2524_n3888# 0.290577f
C98 drain_left.t13 a_n2524_n3888# 0.290577f
C99 drain_left.n2 a_n2524_n3888# 2.63222f
C100 drain_left.t11 a_n2524_n3888# 0.290577f
C101 drain_left.t1 a_n2524_n3888# 0.290577f
C102 drain_left.n3 a_n2524_n3888# 2.62648f
C103 drain_left.n4 a_n2524_n3888# 0.654431f
C104 drain_left.n5 a_n2524_n3888# 1.57526f
C105 drain_left.t0 a_n2524_n3888# 3.35803f
C106 drain_left.t2 a_n2524_n3888# 0.290577f
C107 drain_left.t5 a_n2524_n3888# 0.290577f
C108 drain_left.n6 a_n2524_n3888# 2.62648f
C109 drain_left.n7 a_n2524_n3888# 0.703215f
C110 drain_left.t6 a_n2524_n3888# 0.290577f
C111 drain_left.t3 a_n2524_n3888# 0.290577f
C112 drain_left.n8 a_n2524_n3888# 2.62648f
C113 drain_left.n9 a_n2524_n3888# 0.354678f
C114 drain_left.t7 a_n2524_n3888# 0.290577f
C115 drain_left.t8 a_n2524_n3888# 0.290577f
C116 drain_left.n10 a_n2524_n3888# 2.62647f
C117 drain_left.n11 a_n2524_n3888# 0.574504f
C118 source.t20 a_n2524_n3888# 3.38371f
C119 source.n0 a_n2524_n3888# 1.62429f
C120 source.t15 a_n2524_n3888# 0.301939f
C121 source.t21 a_n2524_n3888# 0.301939f
C122 source.n1 a_n2524_n3888# 2.65228f
C123 source.n2 a_n2524_n3888# 0.410821f
C124 source.t18 a_n2524_n3888# 0.301939f
C125 source.t22 a_n2524_n3888# 0.301939f
C126 source.n3 a_n2524_n3888# 2.65228f
C127 source.n4 a_n2524_n3888# 0.410821f
C128 source.t17 a_n2524_n3888# 0.301939f
C129 source.t24 a_n2524_n3888# 0.301939f
C130 source.n5 a_n2524_n3888# 2.65228f
C131 source.n6 a_n2524_n3888# 0.409405f
C132 source.t8 a_n2524_n3888# 3.38372f
C133 source.n7 a_n2524_n3888# 0.501439f
C134 source.t11 a_n2524_n3888# 0.301939f
C135 source.t2 a_n2524_n3888# 0.301939f
C136 source.n8 a_n2524_n3888# 2.65228f
C137 source.n9 a_n2524_n3888# 0.410821f
C138 source.t5 a_n2524_n3888# 0.301939f
C139 source.t27 a_n2524_n3888# 0.301939f
C140 source.n10 a_n2524_n3888# 2.65228f
C141 source.n11 a_n2524_n3888# 0.410821f
C142 source.t7 a_n2524_n3888# 0.301939f
C143 source.t0 a_n2524_n3888# 0.301939f
C144 source.n12 a_n2524_n3888# 2.65228f
C145 source.n13 a_n2524_n3888# 2.04945f
C146 source.t19 a_n2524_n3888# 0.301939f
C147 source.t23 a_n2524_n3888# 0.301939f
C148 source.n14 a_n2524_n3888# 2.65228f
C149 source.n15 a_n2524_n3888# 2.04946f
C150 source.t16 a_n2524_n3888# 0.301939f
C151 source.t14 a_n2524_n3888# 0.301939f
C152 source.n16 a_n2524_n3888# 2.65228f
C153 source.n17 a_n2524_n3888# 0.410824f
C154 source.t13 a_n2524_n3888# 0.301939f
C155 source.t25 a_n2524_n3888# 0.301939f
C156 source.n18 a_n2524_n3888# 2.65228f
C157 source.n19 a_n2524_n3888# 0.410824f
C158 source.t26 a_n2524_n3888# 3.38371f
C159 source.n20 a_n2524_n3888# 0.501443f
C160 source.t1 a_n2524_n3888# 0.301939f
C161 source.t3 a_n2524_n3888# 0.301939f
C162 source.n21 a_n2524_n3888# 2.65228f
C163 source.n22 a_n2524_n3888# 0.409409f
C164 source.t12 a_n2524_n3888# 0.301939f
C165 source.t10 a_n2524_n3888# 0.301939f
C166 source.n23 a_n2524_n3888# 2.65228f
C167 source.n24 a_n2524_n3888# 0.410824f
C168 source.t6 a_n2524_n3888# 0.301939f
C169 source.t9 a_n2524_n3888# 0.301939f
C170 source.n25 a_n2524_n3888# 2.65228f
C171 source.n26 a_n2524_n3888# 0.410824f
C172 source.t4 a_n2524_n3888# 3.38371f
C173 source.n27 a_n2524_n3888# 0.633139f
C174 source.n28 a_n2524_n3888# 1.88376f
C175 plus.n0 a_n2524_n3888# 0.039192f
C176 plus.t5 a_n2524_n3888# 1.33648f
C177 plus.t6 a_n2524_n3888# 1.33648f
C178 plus.n1 a_n2524_n3888# 0.039192f
C179 plus.t10 a_n2524_n3888# 1.33648f
C180 plus.n2 a_n2524_n3888# 0.521544f
C181 plus.n3 a_n2524_n3888# 0.06528f
C182 plus.t7 a_n2524_n3888# 1.33648f
C183 plus.t8 a_n2524_n3888# 1.33648f
C184 plus.t11 a_n2524_n3888# 1.33648f
C185 plus.n4 a_n2524_n3888# 0.517022f
C186 plus.t13 a_n2524_n3888# 1.35986f
C187 plus.n5 a_n2524_n3888# 0.494645f
C188 plus.n6 a_n2524_n3888# 0.183034f
C189 plus.n7 a_n2524_n3888# 0.008894f
C190 plus.n8 a_n2524_n3888# 0.521544f
C191 plus.n9 a_n2524_n3888# 0.524202f
C192 plus.n10 a_n2524_n3888# 0.078385f
C193 plus.n11 a_n2524_n3888# 0.06528f
C194 plus.n12 a_n2524_n3888# 0.052297f
C195 plus.n13 a_n2524_n3888# 0.008894f
C196 plus.n14 a_n2524_n3888# 0.512167f
C197 plus.n15 a_n2524_n3888# 0.008894f
C198 plus.n16 a_n2524_n3888# 0.513133f
C199 plus.n17 a_n2524_n3888# 0.516016f
C200 plus.n18 a_n2524_n3888# 0.039192f
C201 plus.t4 a_n2524_n3888# 1.33648f
C202 plus.n19 a_n2524_n3888# 0.039192f
C203 plus.t1 a_n2524_n3888# 1.33648f
C204 plus.t9 a_n2524_n3888# 1.33648f
C205 plus.n20 a_n2524_n3888# 0.521544f
C206 plus.n21 a_n2524_n3888# 0.06528f
C207 plus.t2 a_n2524_n3888# 1.33648f
C208 plus.t12 a_n2524_n3888# 1.33648f
C209 plus.t3 a_n2524_n3888# 1.33648f
C210 plus.n22 a_n2524_n3888# 0.517022f
C211 plus.t0 a_n2524_n3888# 1.35986f
C212 plus.n23 a_n2524_n3888# 0.494645f
C213 plus.n24 a_n2524_n3888# 0.183034f
C214 plus.n25 a_n2524_n3888# 0.008894f
C215 plus.n26 a_n2524_n3888# 0.521544f
C216 plus.n27 a_n2524_n3888# 0.524202f
C217 plus.n28 a_n2524_n3888# 0.078385f
C218 plus.n29 a_n2524_n3888# 0.06528f
C219 plus.n30 a_n2524_n3888# 0.052297f
C220 plus.n31 a_n2524_n3888# 0.008894f
C221 plus.n32 a_n2524_n3888# 0.512167f
C222 plus.n33 a_n2524_n3888# 0.008894f
C223 plus.n34 a_n2524_n3888# 0.513133f
C224 plus.n35 a_n2524_n3888# 1.40633f
.ends

