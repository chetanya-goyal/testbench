* NGSPICE file created from diffpair548.ext - technology: sky130A

.subckt diffpair548 minus drain_right drain_left source plus
X0 source.t37 plus.t0 drain_left.t7 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X1 source.t36 plus.t1 drain_left.t6 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X2 source.t3 minus.t0 drain_right.t19 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X3 drain_left.t13 plus.t2 source.t35 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X4 source.t34 plus.t3 drain_left.t12 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X5 source.t33 plus.t4 drain_left.t15 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X6 source.t7 minus.t1 drain_right.t18 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X7 drain_right.t17 minus.t2 source.t8 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X8 a_n2982_n3888# a_n2982_n3888# a_n2982_n3888# a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.7
X9 drain_left.t14 plus.t5 source.t32 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X10 source.t31 plus.t6 drain_left.t3 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X11 source.t30 plus.t7 drain_left.t2 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X12 source.t2 minus.t3 drain_right.t16 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X13 source.t29 plus.t8 drain_left.t1 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X14 drain_left.t0 plus.t9 source.t28 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X15 drain_right.t15 minus.t4 source.t0 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X16 source.t14 minus.t5 drain_right.t14 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X17 drain_right.t13 minus.t6 source.t6 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X18 a_n2982_n3888# a_n2982_n3888# a_n2982_n3888# a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.7
X19 drain_right.t12 minus.t7 source.t10 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X20 drain_right.t11 minus.t8 source.t5 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X21 drain_right.t10 minus.t9 source.t15 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X22 drain_left.t17 plus.t10 source.t27 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X23 drain_right.t9 minus.t10 source.t17 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X24 drain_left.t16 plus.t11 source.t26 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X25 drain_left.t5 plus.t12 source.t25 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X26 drain_right.t8 minus.t11 source.t4 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.7
X27 source.t24 plus.t13 drain_left.t4 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X28 drain_left.t9 plus.t14 source.t23 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X29 drain_left.t8 plus.t15 source.t22 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X30 a_n2982_n3888# a_n2982_n3888# a_n2982_n3888# a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.7
X31 source.t9 minus.t12 drain_right.t7 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X32 drain_right.t6 minus.t13 source.t39 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X33 a_n2982_n3888# a_n2982_n3888# a_n2982_n3888# a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.7
X34 source.t12 minus.t14 drain_right.t5 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X35 drain_left.t19 plus.t16 source.t21 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X36 source.t20 plus.t17 drain_left.t18 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.7
X37 source.t38 minus.t15 drain_right.t4 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X38 drain_left.t11 plus.t18 source.t19 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X39 source.t16 minus.t16 drain_right.t3 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X40 source.t1 minus.t17 drain_right.t2 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X41 source.t18 plus.t19 drain_left.t10 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X42 source.t11 minus.t18 drain_right.t1 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
X43 drain_right.t0 minus.t19 source.t13 a_n2982_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.7
R0 plus.n9 plus.t7 597.941
R1 plus.n43 plus.t2 597.941
R2 plus.n32 plus.t5 572.548
R3 plus.n30 plus.t19 572.548
R4 plus.n2 plus.t10 572.548
R5 plus.n24 plus.t1 572.548
R6 plus.n4 plus.t12 572.548
R7 plus.n18 plus.t6 572.548
R8 plus.n6 plus.t11 572.548
R9 plus.n12 plus.t4 572.548
R10 plus.n8 plus.t15 572.548
R11 plus.n66 plus.t17 572.548
R12 plus.n64 plus.t16 572.548
R13 plus.n36 plus.t0 572.548
R14 plus.n58 plus.t9 572.548
R15 plus.n38 plus.t8 572.548
R16 plus.n52 plus.t14 572.548
R17 plus.n40 plus.t13 572.548
R18 plus.n46 plus.t18 572.548
R19 plus.n42 plus.t3 572.548
R20 plus.n11 plus.n10 161.3
R21 plus.n12 plus.n7 161.3
R22 plus.n14 plus.n13 161.3
R23 plus.n15 plus.n6 161.3
R24 plus.n17 plus.n16 161.3
R25 plus.n18 plus.n5 161.3
R26 plus.n20 plus.n19 161.3
R27 plus.n21 plus.n4 161.3
R28 plus.n23 plus.n22 161.3
R29 plus.n24 plus.n3 161.3
R30 plus.n26 plus.n25 161.3
R31 plus.n27 plus.n2 161.3
R32 plus.n29 plus.n28 161.3
R33 plus.n30 plus.n1 161.3
R34 plus.n31 plus.n0 161.3
R35 plus.n33 plus.n32 161.3
R36 plus.n45 plus.n44 161.3
R37 plus.n46 plus.n41 161.3
R38 plus.n48 plus.n47 161.3
R39 plus.n49 plus.n40 161.3
R40 plus.n51 plus.n50 161.3
R41 plus.n52 plus.n39 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n55 plus.n38 161.3
R44 plus.n57 plus.n56 161.3
R45 plus.n58 plus.n37 161.3
R46 plus.n60 plus.n59 161.3
R47 plus.n61 plus.n36 161.3
R48 plus.n63 plus.n62 161.3
R49 plus.n64 plus.n35 161.3
R50 plus.n65 plus.n34 161.3
R51 plus.n67 plus.n66 161.3
R52 plus.n10 plus.n9 45.0031
R53 plus.n44 plus.n43 45.0031
R54 plus.n32 plus.n31 41.6278
R55 plus.n66 plus.n65 41.6278
R56 plus.n30 plus.n29 37.246
R57 plus.n11 plus.n8 37.246
R58 plus.n64 plus.n63 37.246
R59 plus.n45 plus.n42 37.246
R60 plus plus.n67 35.6013
R61 plus.n25 plus.n2 32.8641
R62 plus.n13 plus.n12 32.8641
R63 plus.n59 plus.n36 32.8641
R64 plus.n47 plus.n46 32.8641
R65 plus.n24 plus.n23 28.4823
R66 plus.n17 plus.n6 28.4823
R67 plus.n58 plus.n57 28.4823
R68 plus.n51 plus.n40 28.4823
R69 plus.n19 plus.n18 24.1005
R70 plus.n19 plus.n4 24.1005
R71 plus.n53 plus.n38 24.1005
R72 plus.n53 plus.n52 24.1005
R73 plus.n23 plus.n4 19.7187
R74 plus.n18 plus.n17 19.7187
R75 plus.n57 plus.n38 19.7187
R76 plus.n52 plus.n51 19.7187
R77 plus.n9 plus.n8 15.6319
R78 plus.n43 plus.n42 15.6319
R79 plus.n25 plus.n24 15.3369
R80 plus.n13 plus.n6 15.3369
R81 plus.n59 plus.n58 15.3369
R82 plus.n47 plus.n40 15.3369
R83 plus plus.n33 13.4475
R84 plus.n29 plus.n2 10.955
R85 plus.n12 plus.n11 10.955
R86 plus.n63 plus.n36 10.955
R87 plus.n46 plus.n45 10.955
R88 plus.n31 plus.n30 6.57323
R89 plus.n65 plus.n64 6.57323
R90 plus.n10 plus.n7 0.189894
R91 plus.n14 plus.n7 0.189894
R92 plus.n15 plus.n14 0.189894
R93 plus.n16 plus.n15 0.189894
R94 plus.n16 plus.n5 0.189894
R95 plus.n20 plus.n5 0.189894
R96 plus.n21 plus.n20 0.189894
R97 plus.n22 plus.n21 0.189894
R98 plus.n22 plus.n3 0.189894
R99 plus.n26 plus.n3 0.189894
R100 plus.n27 plus.n26 0.189894
R101 plus.n28 plus.n27 0.189894
R102 plus.n28 plus.n1 0.189894
R103 plus.n1 plus.n0 0.189894
R104 plus.n33 plus.n0 0.189894
R105 plus.n67 plus.n34 0.189894
R106 plus.n35 plus.n34 0.189894
R107 plus.n62 plus.n35 0.189894
R108 plus.n62 plus.n61 0.189894
R109 plus.n61 plus.n60 0.189894
R110 plus.n60 plus.n37 0.189894
R111 plus.n56 plus.n37 0.189894
R112 plus.n56 plus.n55 0.189894
R113 plus.n55 plus.n54 0.189894
R114 plus.n54 plus.n39 0.189894
R115 plus.n50 plus.n39 0.189894
R116 plus.n50 plus.n49 0.189894
R117 plus.n49 plus.n48 0.189894
R118 plus.n48 plus.n41 0.189894
R119 plus.n44 plus.n41 0.189894
R120 drain_left.n10 drain_left.n8 61.7677
R121 drain_left.n6 drain_left.n4 61.7675
R122 drain_left.n2 drain_left.n0 61.7675
R123 drain_left.n14 drain_left.n13 60.8798
R124 drain_left.n12 drain_left.n11 60.8798
R125 drain_left.n10 drain_left.n9 60.8798
R126 drain_left.n16 drain_left.n15 60.8796
R127 drain_left.n7 drain_left.n3 60.8796
R128 drain_left.n6 drain_left.n5 60.8796
R129 drain_left.n2 drain_left.n1 60.8796
R130 drain_left drain_left.n7 36.7433
R131 drain_left drain_left.n16 6.54115
R132 drain_left.n3 drain_left.t1 1.3205
R133 drain_left.n3 drain_left.t9 1.3205
R134 drain_left.n4 drain_left.t12 1.3205
R135 drain_left.n4 drain_left.t13 1.3205
R136 drain_left.n5 drain_left.t4 1.3205
R137 drain_left.n5 drain_left.t11 1.3205
R138 drain_left.n1 drain_left.t7 1.3205
R139 drain_left.n1 drain_left.t0 1.3205
R140 drain_left.n0 drain_left.t18 1.3205
R141 drain_left.n0 drain_left.t19 1.3205
R142 drain_left.n15 drain_left.t10 1.3205
R143 drain_left.n15 drain_left.t14 1.3205
R144 drain_left.n13 drain_left.t6 1.3205
R145 drain_left.n13 drain_left.t17 1.3205
R146 drain_left.n11 drain_left.t3 1.3205
R147 drain_left.n11 drain_left.t5 1.3205
R148 drain_left.n9 drain_left.t15 1.3205
R149 drain_left.n9 drain_left.t16 1.3205
R150 drain_left.n8 drain_left.t2 1.3205
R151 drain_left.n8 drain_left.t8 1.3205
R152 drain_left.n12 drain_left.n10 0.888431
R153 drain_left.n14 drain_left.n12 0.888431
R154 drain_left.n16 drain_left.n14 0.888431
R155 drain_left.n7 drain_left.n6 0.833085
R156 drain_left.n7 drain_left.n2 0.833085
R157 source.n9 source.t30 45.521
R158 source.n10 source.t4 45.521
R159 source.n19 source.t9 45.521
R160 source.n39 source.t15 45.5208
R161 source.n30 source.t14 45.5208
R162 source.n29 source.t35 45.5208
R163 source.n20 source.t20 45.5208
R164 source.n0 source.t32 45.5208
R165 source.n2 source.n1 44.201
R166 source.n4 source.n3 44.201
R167 source.n6 source.n5 44.201
R168 source.n8 source.n7 44.201
R169 source.n12 source.n11 44.201
R170 source.n14 source.n13 44.201
R171 source.n16 source.n15 44.201
R172 source.n18 source.n17 44.201
R173 source.n38 source.n37 44.2008
R174 source.n36 source.n35 44.2008
R175 source.n34 source.n33 44.2008
R176 source.n32 source.n31 44.2008
R177 source.n28 source.n27 44.2008
R178 source.n26 source.n25 44.2008
R179 source.n24 source.n23 44.2008
R180 source.n22 source.n21 44.2008
R181 source.n20 source.n19 24.4484
R182 source.n40 source.n0 18.7415
R183 source.n40 source.n39 5.7074
R184 source.n37 source.t39 1.3205
R185 source.n37 source.t12 1.3205
R186 source.n35 source.t13 1.3205
R187 source.n35 source.t11 1.3205
R188 source.n33 source.t8 1.3205
R189 source.n33 source.t2 1.3205
R190 source.n31 source.t6 1.3205
R191 source.n31 source.t3 1.3205
R192 source.n27 source.t19 1.3205
R193 source.n27 source.t34 1.3205
R194 source.n25 source.t23 1.3205
R195 source.n25 source.t24 1.3205
R196 source.n23 source.t28 1.3205
R197 source.n23 source.t29 1.3205
R198 source.n21 source.t21 1.3205
R199 source.n21 source.t37 1.3205
R200 source.n1 source.t27 1.3205
R201 source.n1 source.t18 1.3205
R202 source.n3 source.t25 1.3205
R203 source.n3 source.t36 1.3205
R204 source.n5 source.t26 1.3205
R205 source.n5 source.t31 1.3205
R206 source.n7 source.t22 1.3205
R207 source.n7 source.t33 1.3205
R208 source.n11 source.t17 1.3205
R209 source.n11 source.t7 1.3205
R210 source.n13 source.t5 1.3205
R211 source.n13 source.t16 1.3205
R212 source.n15 source.t10 1.3205
R213 source.n15 source.t1 1.3205
R214 source.n17 source.t0 1.3205
R215 source.n17 source.t38 1.3205
R216 source.n19 source.n18 0.888431
R217 source.n18 source.n16 0.888431
R218 source.n16 source.n14 0.888431
R219 source.n14 source.n12 0.888431
R220 source.n12 source.n10 0.888431
R221 source.n9 source.n8 0.888431
R222 source.n8 source.n6 0.888431
R223 source.n6 source.n4 0.888431
R224 source.n4 source.n2 0.888431
R225 source.n2 source.n0 0.888431
R226 source.n22 source.n20 0.888431
R227 source.n24 source.n22 0.888431
R228 source.n26 source.n24 0.888431
R229 source.n28 source.n26 0.888431
R230 source.n29 source.n28 0.888431
R231 source.n32 source.n30 0.888431
R232 source.n34 source.n32 0.888431
R233 source.n36 source.n34 0.888431
R234 source.n38 source.n36 0.888431
R235 source.n39 source.n38 0.888431
R236 source.n10 source.n9 0.470328
R237 source.n30 source.n29 0.470328
R238 source source.n40 0.188
R239 minus.n9 minus.t11 597.941
R240 minus.n43 minus.t5 597.941
R241 minus.n8 minus.t1 572.548
R242 minus.n12 minus.t10 572.548
R243 minus.n14 minus.t16 572.548
R244 minus.n18 minus.t8 572.548
R245 minus.n20 minus.t17 572.548
R246 minus.n24 minus.t7 572.548
R247 minus.n26 minus.t15 572.548
R248 minus.n30 minus.t4 572.548
R249 minus.n32 minus.t12 572.548
R250 minus.n42 minus.t6 572.548
R251 minus.n46 minus.t0 572.548
R252 minus.n48 minus.t2 572.548
R253 minus.n52 minus.t3 572.548
R254 minus.n54 minus.t19 572.548
R255 minus.n58 minus.t18 572.548
R256 minus.n60 minus.t13 572.548
R257 minus.n64 minus.t14 572.548
R258 minus.n66 minus.t9 572.548
R259 minus.n33 minus.n32 161.3
R260 minus.n31 minus.n0 161.3
R261 minus.n30 minus.n29 161.3
R262 minus.n28 minus.n1 161.3
R263 minus.n27 minus.n26 161.3
R264 minus.n25 minus.n2 161.3
R265 minus.n24 minus.n23 161.3
R266 minus.n22 minus.n3 161.3
R267 minus.n21 minus.n20 161.3
R268 minus.n19 minus.n4 161.3
R269 minus.n18 minus.n17 161.3
R270 minus.n16 minus.n5 161.3
R271 minus.n15 minus.n14 161.3
R272 minus.n13 minus.n6 161.3
R273 minus.n12 minus.n11 161.3
R274 minus.n10 minus.n7 161.3
R275 minus.n67 minus.n66 161.3
R276 minus.n65 minus.n34 161.3
R277 minus.n64 minus.n63 161.3
R278 minus.n62 minus.n35 161.3
R279 minus.n61 minus.n60 161.3
R280 minus.n59 minus.n36 161.3
R281 minus.n58 minus.n57 161.3
R282 minus.n56 minus.n37 161.3
R283 minus.n55 minus.n54 161.3
R284 minus.n53 minus.n38 161.3
R285 minus.n52 minus.n51 161.3
R286 minus.n50 minus.n39 161.3
R287 minus.n49 minus.n48 161.3
R288 minus.n47 minus.n40 161.3
R289 minus.n46 minus.n45 161.3
R290 minus.n44 minus.n41 161.3
R291 minus.n10 minus.n9 45.0031
R292 minus.n44 minus.n43 45.0031
R293 minus.n68 minus.n33 42.8566
R294 minus.n32 minus.n31 41.6278
R295 minus.n66 minus.n65 41.6278
R296 minus.n8 minus.n7 37.246
R297 minus.n30 minus.n1 37.246
R298 minus.n42 minus.n41 37.246
R299 minus.n64 minus.n35 37.246
R300 minus.n13 minus.n12 32.8641
R301 minus.n26 minus.n25 32.8641
R302 minus.n47 minus.n46 32.8641
R303 minus.n60 minus.n59 32.8641
R304 minus.n14 minus.n5 28.4823
R305 minus.n24 minus.n3 28.4823
R306 minus.n48 minus.n39 28.4823
R307 minus.n58 minus.n37 28.4823
R308 minus.n20 minus.n19 24.1005
R309 minus.n19 minus.n18 24.1005
R310 minus.n53 minus.n52 24.1005
R311 minus.n54 minus.n53 24.1005
R312 minus.n18 minus.n5 19.7187
R313 minus.n20 minus.n3 19.7187
R314 minus.n52 minus.n39 19.7187
R315 minus.n54 minus.n37 19.7187
R316 minus.n9 minus.n8 15.6319
R317 minus.n43 minus.n42 15.6319
R318 minus.n14 minus.n13 15.3369
R319 minus.n25 minus.n24 15.3369
R320 minus.n48 minus.n47 15.3369
R321 minus.n59 minus.n58 15.3369
R322 minus.n12 minus.n7 10.955
R323 minus.n26 minus.n1 10.955
R324 minus.n46 minus.n41 10.955
R325 minus.n60 minus.n35 10.955
R326 minus.n68 minus.n67 6.66717
R327 minus.n31 minus.n30 6.57323
R328 minus.n65 minus.n64 6.57323
R329 minus.n33 minus.n0 0.189894
R330 minus.n29 minus.n0 0.189894
R331 minus.n29 minus.n28 0.189894
R332 minus.n28 minus.n27 0.189894
R333 minus.n27 minus.n2 0.189894
R334 minus.n23 minus.n2 0.189894
R335 minus.n23 minus.n22 0.189894
R336 minus.n22 minus.n21 0.189894
R337 minus.n21 minus.n4 0.189894
R338 minus.n17 minus.n4 0.189894
R339 minus.n17 minus.n16 0.189894
R340 minus.n16 minus.n15 0.189894
R341 minus.n15 minus.n6 0.189894
R342 minus.n11 minus.n6 0.189894
R343 minus.n11 minus.n10 0.189894
R344 minus.n45 minus.n44 0.189894
R345 minus.n45 minus.n40 0.189894
R346 minus.n49 minus.n40 0.189894
R347 minus.n50 minus.n49 0.189894
R348 minus.n51 minus.n50 0.189894
R349 minus.n51 minus.n38 0.189894
R350 minus.n55 minus.n38 0.189894
R351 minus.n56 minus.n55 0.189894
R352 minus.n57 minus.n56 0.189894
R353 minus.n57 minus.n36 0.189894
R354 minus.n61 minus.n36 0.189894
R355 minus.n62 minus.n61 0.189894
R356 minus.n63 minus.n62 0.189894
R357 minus.n63 minus.n34 0.189894
R358 minus.n67 minus.n34 0.189894
R359 minus minus.n68 0.188
R360 drain_right.n10 drain_right.n8 61.7676
R361 drain_right.n6 drain_right.n4 61.7675
R362 drain_right.n2 drain_right.n0 61.7675
R363 drain_right.n10 drain_right.n9 60.8798
R364 drain_right.n12 drain_right.n11 60.8798
R365 drain_right.n14 drain_right.n13 60.8798
R366 drain_right.n16 drain_right.n15 60.8798
R367 drain_right.n7 drain_right.n3 60.8796
R368 drain_right.n6 drain_right.n5 60.8796
R369 drain_right.n2 drain_right.n1 60.8796
R370 drain_right drain_right.n7 36.19
R371 drain_right drain_right.n16 6.54115
R372 drain_right.n3 drain_right.t16 1.3205
R373 drain_right.n3 drain_right.t0 1.3205
R374 drain_right.n4 drain_right.t5 1.3205
R375 drain_right.n4 drain_right.t10 1.3205
R376 drain_right.n5 drain_right.t1 1.3205
R377 drain_right.n5 drain_right.t6 1.3205
R378 drain_right.n1 drain_right.t19 1.3205
R379 drain_right.n1 drain_right.t17 1.3205
R380 drain_right.n0 drain_right.t14 1.3205
R381 drain_right.n0 drain_right.t13 1.3205
R382 drain_right.n8 drain_right.t18 1.3205
R383 drain_right.n8 drain_right.t8 1.3205
R384 drain_right.n9 drain_right.t3 1.3205
R385 drain_right.n9 drain_right.t9 1.3205
R386 drain_right.n11 drain_right.t2 1.3205
R387 drain_right.n11 drain_right.t11 1.3205
R388 drain_right.n13 drain_right.t4 1.3205
R389 drain_right.n13 drain_right.t12 1.3205
R390 drain_right.n15 drain_right.t7 1.3205
R391 drain_right.n15 drain_right.t15 1.3205
R392 drain_right.n16 drain_right.n14 0.888431
R393 drain_right.n14 drain_right.n12 0.888431
R394 drain_right.n12 drain_right.n10 0.888431
R395 drain_right.n7 drain_right.n6 0.833085
R396 drain_right.n7 drain_right.n2 0.833085
C0 drain_left minus 0.173554f
C1 plus minus 7.42109f
C2 source drain_right 29.06f
C3 drain_left plus 15.8639f
C4 source minus 15.6064f
C5 drain_right minus 15.566401f
C6 source drain_left 29.0576f
C7 drain_left drain_right 1.59885f
C8 source plus 15.620501f
C9 plus drain_right 0.454687f
C10 drain_right a_n2982_n3888# 7.88675f
C11 drain_left a_n2982_n3888# 8.30361f
C12 source a_n2982_n3888# 11.100306f
C13 minus a_n2982_n3888# 12.203388f
C14 plus a_n2982_n3888# 14.16684f
C15 drain_right.t14 a_n2982_n3888# 0.322669f
C16 drain_right.t13 a_n2982_n3888# 0.322669f
C17 drain_right.n0 a_n2982_n3888# 2.92215f
C18 drain_right.t19 a_n2982_n3888# 0.322669f
C19 drain_right.t17 a_n2982_n3888# 0.322669f
C20 drain_right.n1 a_n2982_n3888# 2.91655f
C21 drain_right.n2 a_n2982_n3888# 0.758722f
C22 drain_right.t16 a_n2982_n3888# 0.322669f
C23 drain_right.t0 a_n2982_n3888# 0.322669f
C24 drain_right.n3 a_n2982_n3888# 2.91655f
C25 drain_right.t5 a_n2982_n3888# 0.322669f
C26 drain_right.t10 a_n2982_n3888# 0.322669f
C27 drain_right.n4 a_n2982_n3888# 2.92215f
C28 drain_right.t1 a_n2982_n3888# 0.322669f
C29 drain_right.t6 a_n2982_n3888# 0.322669f
C30 drain_right.n5 a_n2982_n3888# 2.91655f
C31 drain_right.n6 a_n2982_n3888# 0.758722f
C32 drain_right.n7 a_n2982_n3888# 2.1213f
C33 drain_right.t18 a_n2982_n3888# 0.322669f
C34 drain_right.t8 a_n2982_n3888# 0.322669f
C35 drain_right.n8 a_n2982_n3888# 2.92214f
C36 drain_right.t3 a_n2982_n3888# 0.322669f
C37 drain_right.t9 a_n2982_n3888# 0.322669f
C38 drain_right.n9 a_n2982_n3888# 2.91655f
C39 drain_right.n10 a_n2982_n3888# 0.762824f
C40 drain_right.t2 a_n2982_n3888# 0.322669f
C41 drain_right.t11 a_n2982_n3888# 0.322669f
C42 drain_right.n11 a_n2982_n3888# 2.91655f
C43 drain_right.n12 a_n2982_n3888# 0.378726f
C44 drain_right.t4 a_n2982_n3888# 0.322669f
C45 drain_right.t12 a_n2982_n3888# 0.322669f
C46 drain_right.n13 a_n2982_n3888# 2.91655f
C47 drain_right.n14 a_n2982_n3888# 0.378726f
C48 drain_right.t7 a_n2982_n3888# 0.322669f
C49 drain_right.t15 a_n2982_n3888# 0.322669f
C50 drain_right.n15 a_n2982_n3888# 2.91655f
C51 drain_right.n16 a_n2982_n3888# 0.619502f
C52 minus.n0 a_n2982_n3888# 0.039575f
C53 minus.n1 a_n2982_n3888# 0.00898f
C54 minus.t4 a_n2982_n3888# 1.18082f
C55 minus.n2 a_n2982_n3888# 0.039575f
C56 minus.n3 a_n2982_n3888# 0.00898f
C57 minus.t7 a_n2982_n3888# 1.18082f
C58 minus.n4 a_n2982_n3888# 0.039575f
C59 minus.n5 a_n2982_n3888# 0.00898f
C60 minus.t8 a_n2982_n3888# 1.18082f
C61 minus.n6 a_n2982_n3888# 0.039575f
C62 minus.n7 a_n2982_n3888# 0.00898f
C63 minus.t10 a_n2982_n3888# 1.18082f
C64 minus.t11 a_n2982_n3888# 1.20019f
C65 minus.t1 a_n2982_n3888# 1.18082f
C66 minus.n8 a_n2982_n3888# 0.462301f
C67 minus.n9 a_n2982_n3888# 0.439154f
C68 minus.n10 a_n2982_n3888# 0.16892f
C69 minus.n11 a_n2982_n3888# 0.039575f
C70 minus.n12 a_n2982_n3888# 0.455682f
C71 minus.n13 a_n2982_n3888# 0.00898f
C72 minus.t16 a_n2982_n3888# 1.18082f
C73 minus.n14 a_n2982_n3888# 0.455682f
C74 minus.n15 a_n2982_n3888# 0.039575f
C75 minus.n16 a_n2982_n3888# 0.039575f
C76 minus.n17 a_n2982_n3888# 0.039575f
C77 minus.n18 a_n2982_n3888# 0.455682f
C78 minus.n19 a_n2982_n3888# 0.00898f
C79 minus.t17 a_n2982_n3888# 1.18082f
C80 minus.n20 a_n2982_n3888# 0.455682f
C81 minus.n21 a_n2982_n3888# 0.039575f
C82 minus.n22 a_n2982_n3888# 0.039575f
C83 minus.n23 a_n2982_n3888# 0.039575f
C84 minus.n24 a_n2982_n3888# 0.455682f
C85 minus.n25 a_n2982_n3888# 0.00898f
C86 minus.t15 a_n2982_n3888# 1.18082f
C87 minus.n26 a_n2982_n3888# 0.455682f
C88 minus.n27 a_n2982_n3888# 0.039575f
C89 minus.n28 a_n2982_n3888# 0.039575f
C90 minus.n29 a_n2982_n3888# 0.039575f
C91 minus.n30 a_n2982_n3888# 0.455682f
C92 minus.n31 a_n2982_n3888# 0.00898f
C93 minus.t12 a_n2982_n3888# 1.18082f
C94 minus.n32 a_n2982_n3888# 0.455316f
C95 minus.n33 a_n2982_n3888# 1.80961f
C96 minus.n34 a_n2982_n3888# 0.039575f
C97 minus.n35 a_n2982_n3888# 0.00898f
C98 minus.n36 a_n2982_n3888# 0.039575f
C99 minus.n37 a_n2982_n3888# 0.00898f
C100 minus.n38 a_n2982_n3888# 0.039575f
C101 minus.n39 a_n2982_n3888# 0.00898f
C102 minus.n40 a_n2982_n3888# 0.039575f
C103 minus.n41 a_n2982_n3888# 0.00898f
C104 minus.t5 a_n2982_n3888# 1.20019f
C105 minus.t6 a_n2982_n3888# 1.18082f
C106 minus.n42 a_n2982_n3888# 0.462301f
C107 minus.n43 a_n2982_n3888# 0.439154f
C108 minus.n44 a_n2982_n3888# 0.16892f
C109 minus.n45 a_n2982_n3888# 0.039575f
C110 minus.t0 a_n2982_n3888# 1.18082f
C111 minus.n46 a_n2982_n3888# 0.455682f
C112 minus.n47 a_n2982_n3888# 0.00898f
C113 minus.t2 a_n2982_n3888# 1.18082f
C114 minus.n48 a_n2982_n3888# 0.455682f
C115 minus.n49 a_n2982_n3888# 0.039575f
C116 minus.n50 a_n2982_n3888# 0.039575f
C117 minus.n51 a_n2982_n3888# 0.039575f
C118 minus.t3 a_n2982_n3888# 1.18082f
C119 minus.n52 a_n2982_n3888# 0.455682f
C120 minus.n53 a_n2982_n3888# 0.00898f
C121 minus.t19 a_n2982_n3888# 1.18082f
C122 minus.n54 a_n2982_n3888# 0.455682f
C123 minus.n55 a_n2982_n3888# 0.039575f
C124 minus.n56 a_n2982_n3888# 0.039575f
C125 minus.n57 a_n2982_n3888# 0.039575f
C126 minus.t18 a_n2982_n3888# 1.18082f
C127 minus.n58 a_n2982_n3888# 0.455682f
C128 minus.n59 a_n2982_n3888# 0.00898f
C129 minus.t13 a_n2982_n3888# 1.18082f
C130 minus.n60 a_n2982_n3888# 0.455682f
C131 minus.n61 a_n2982_n3888# 0.039575f
C132 minus.n62 a_n2982_n3888# 0.039575f
C133 minus.n63 a_n2982_n3888# 0.039575f
C134 minus.t14 a_n2982_n3888# 1.18082f
C135 minus.n64 a_n2982_n3888# 0.455682f
C136 minus.n65 a_n2982_n3888# 0.00898f
C137 minus.t9 a_n2982_n3888# 1.18082f
C138 minus.n66 a_n2982_n3888# 0.455316f
C139 minus.n67 a_n2982_n3888# 0.274193f
C140 minus.n68 a_n2982_n3888# 2.15234f
C141 source.t32 a_n2982_n3888# 3.16483f
C142 source.n0 a_n2982_n3888# 1.50856f
C143 source.t27 a_n2982_n3888# 0.282407f
C144 source.t18 a_n2982_n3888# 0.282407f
C145 source.n1 a_n2982_n3888# 2.48071f
C146 source.n2 a_n2982_n3888# 0.371009f
C147 source.t25 a_n2982_n3888# 0.282407f
C148 source.t36 a_n2982_n3888# 0.282407f
C149 source.n3 a_n2982_n3888# 2.48071f
C150 source.n4 a_n2982_n3888# 0.371009f
C151 source.t26 a_n2982_n3888# 0.282407f
C152 source.t31 a_n2982_n3888# 0.282407f
C153 source.n5 a_n2982_n3888# 2.48071f
C154 source.n6 a_n2982_n3888# 0.371009f
C155 source.t22 a_n2982_n3888# 0.282407f
C156 source.t33 a_n2982_n3888# 0.282407f
C157 source.n7 a_n2982_n3888# 2.48071f
C158 source.n8 a_n2982_n3888# 0.371009f
C159 source.t30 a_n2982_n3888# 3.16483f
C160 source.n9 a_n2982_n3888# 0.424992f
C161 source.t4 a_n2982_n3888# 3.16483f
C162 source.n10 a_n2982_n3888# 0.424992f
C163 source.t17 a_n2982_n3888# 0.282407f
C164 source.t7 a_n2982_n3888# 0.282407f
C165 source.n11 a_n2982_n3888# 2.48071f
C166 source.n12 a_n2982_n3888# 0.371009f
C167 source.t5 a_n2982_n3888# 0.282407f
C168 source.t16 a_n2982_n3888# 0.282407f
C169 source.n13 a_n2982_n3888# 2.48071f
C170 source.n14 a_n2982_n3888# 0.371009f
C171 source.t10 a_n2982_n3888# 0.282407f
C172 source.t1 a_n2982_n3888# 0.282407f
C173 source.n15 a_n2982_n3888# 2.48071f
C174 source.n16 a_n2982_n3888# 0.371009f
C175 source.t0 a_n2982_n3888# 0.282407f
C176 source.t38 a_n2982_n3888# 0.282407f
C177 source.n17 a_n2982_n3888# 2.48071f
C178 source.n18 a_n2982_n3888# 0.371009f
C179 source.t9 a_n2982_n3888# 3.16483f
C180 source.n19 a_n2982_n3888# 1.91494f
C181 source.t20 a_n2982_n3888# 3.16483f
C182 source.n20 a_n2982_n3888# 1.91494f
C183 source.t21 a_n2982_n3888# 0.282407f
C184 source.t37 a_n2982_n3888# 0.282407f
C185 source.n21 a_n2982_n3888# 2.48071f
C186 source.n22 a_n2982_n3888# 0.371013f
C187 source.t28 a_n2982_n3888# 0.282407f
C188 source.t29 a_n2982_n3888# 0.282407f
C189 source.n23 a_n2982_n3888# 2.48071f
C190 source.n24 a_n2982_n3888# 0.371013f
C191 source.t23 a_n2982_n3888# 0.282407f
C192 source.t24 a_n2982_n3888# 0.282407f
C193 source.n25 a_n2982_n3888# 2.48071f
C194 source.n26 a_n2982_n3888# 0.371013f
C195 source.t19 a_n2982_n3888# 0.282407f
C196 source.t34 a_n2982_n3888# 0.282407f
C197 source.n27 a_n2982_n3888# 2.48071f
C198 source.n28 a_n2982_n3888# 0.371013f
C199 source.t35 a_n2982_n3888# 3.16483f
C200 source.n29 a_n2982_n3888# 0.424996f
C201 source.t14 a_n2982_n3888# 3.16483f
C202 source.n30 a_n2982_n3888# 0.424996f
C203 source.t6 a_n2982_n3888# 0.282407f
C204 source.t3 a_n2982_n3888# 0.282407f
C205 source.n31 a_n2982_n3888# 2.48071f
C206 source.n32 a_n2982_n3888# 0.371013f
C207 source.t8 a_n2982_n3888# 0.282407f
C208 source.t2 a_n2982_n3888# 0.282407f
C209 source.n33 a_n2982_n3888# 2.48071f
C210 source.n34 a_n2982_n3888# 0.371013f
C211 source.t13 a_n2982_n3888# 0.282407f
C212 source.t11 a_n2982_n3888# 0.282407f
C213 source.n35 a_n2982_n3888# 2.48071f
C214 source.n36 a_n2982_n3888# 0.371013f
C215 source.t39 a_n2982_n3888# 0.282407f
C216 source.t12 a_n2982_n3888# 0.282407f
C217 source.n37 a_n2982_n3888# 2.48071f
C218 source.n38 a_n2982_n3888# 0.371013f
C219 source.t15 a_n2982_n3888# 3.16483f
C220 source.n39 a_n2982_n3888# 0.580407f
C221 source.n40 a_n2982_n3888# 1.75787f
C222 drain_left.t18 a_n2982_n3888# 0.324063f
C223 drain_left.t19 a_n2982_n3888# 0.324063f
C224 drain_left.n0 a_n2982_n3888# 2.93477f
C225 drain_left.t7 a_n2982_n3888# 0.324063f
C226 drain_left.t0 a_n2982_n3888# 0.324063f
C227 drain_left.n1 a_n2982_n3888# 2.92915f
C228 drain_left.n2 a_n2982_n3888# 0.761999f
C229 drain_left.t1 a_n2982_n3888# 0.324063f
C230 drain_left.t9 a_n2982_n3888# 0.324063f
C231 drain_left.n3 a_n2982_n3888# 2.92915f
C232 drain_left.t12 a_n2982_n3888# 0.324063f
C233 drain_left.t13 a_n2982_n3888# 0.324063f
C234 drain_left.n4 a_n2982_n3888# 2.93477f
C235 drain_left.t4 a_n2982_n3888# 0.324063f
C236 drain_left.t11 a_n2982_n3888# 0.324063f
C237 drain_left.n5 a_n2982_n3888# 2.92915f
C238 drain_left.n6 a_n2982_n3888# 0.761999f
C239 drain_left.n7 a_n2982_n3888# 2.18638f
C240 drain_left.t2 a_n2982_n3888# 0.324063f
C241 drain_left.t8 a_n2982_n3888# 0.324063f
C242 drain_left.n8 a_n2982_n3888# 2.93477f
C243 drain_left.t15 a_n2982_n3888# 0.324063f
C244 drain_left.t16 a_n2982_n3888# 0.324063f
C245 drain_left.n9 a_n2982_n3888# 2.92915f
C246 drain_left.n10 a_n2982_n3888# 0.766109f
C247 drain_left.t3 a_n2982_n3888# 0.324063f
C248 drain_left.t5 a_n2982_n3888# 0.324063f
C249 drain_left.n11 a_n2982_n3888# 2.92915f
C250 drain_left.n12 a_n2982_n3888# 0.380362f
C251 drain_left.t6 a_n2982_n3888# 0.324063f
C252 drain_left.t17 a_n2982_n3888# 0.324063f
C253 drain_left.n13 a_n2982_n3888# 2.92915f
C254 drain_left.n14 a_n2982_n3888# 0.380362f
C255 drain_left.t10 a_n2982_n3888# 0.324063f
C256 drain_left.t14 a_n2982_n3888# 0.324063f
C257 drain_left.n15 a_n2982_n3888# 2.92914f
C258 drain_left.n16 a_n2982_n3888# 0.622188f
C259 plus.n0 a_n2982_n3888# 0.039965f
C260 plus.t5 a_n2982_n3888# 1.19247f
C261 plus.t19 a_n2982_n3888# 1.19247f
C262 plus.n1 a_n2982_n3888# 0.039965f
C263 plus.t10 a_n2982_n3888# 1.19247f
C264 plus.n2 a_n2982_n3888# 0.460178f
C265 plus.n3 a_n2982_n3888# 0.039965f
C266 plus.t1 a_n2982_n3888# 1.19247f
C267 plus.t12 a_n2982_n3888# 1.19247f
C268 plus.n4 a_n2982_n3888# 0.460178f
C269 plus.n5 a_n2982_n3888# 0.039965f
C270 plus.t6 a_n2982_n3888# 1.19247f
C271 plus.t11 a_n2982_n3888# 1.19247f
C272 plus.n6 a_n2982_n3888# 0.460178f
C273 plus.n7 a_n2982_n3888# 0.039965f
C274 plus.t4 a_n2982_n3888# 1.19247f
C275 plus.t15 a_n2982_n3888# 1.19247f
C276 plus.n8 a_n2982_n3888# 0.466862f
C277 plus.t7 a_n2982_n3888# 1.21203f
C278 plus.n9 a_n2982_n3888# 0.443487f
C279 plus.n10 a_n2982_n3888# 0.170587f
C280 plus.n11 a_n2982_n3888# 0.009069f
C281 plus.n12 a_n2982_n3888# 0.460178f
C282 plus.n13 a_n2982_n3888# 0.009069f
C283 plus.n14 a_n2982_n3888# 0.039965f
C284 plus.n15 a_n2982_n3888# 0.039965f
C285 plus.n16 a_n2982_n3888# 0.039965f
C286 plus.n17 a_n2982_n3888# 0.009069f
C287 plus.n18 a_n2982_n3888# 0.460178f
C288 plus.n19 a_n2982_n3888# 0.009069f
C289 plus.n20 a_n2982_n3888# 0.039965f
C290 plus.n21 a_n2982_n3888# 0.039965f
C291 plus.n22 a_n2982_n3888# 0.039965f
C292 plus.n23 a_n2982_n3888# 0.009069f
C293 plus.n24 a_n2982_n3888# 0.460178f
C294 plus.n25 a_n2982_n3888# 0.009069f
C295 plus.n26 a_n2982_n3888# 0.039965f
C296 plus.n27 a_n2982_n3888# 0.039965f
C297 plus.n28 a_n2982_n3888# 0.039965f
C298 plus.n29 a_n2982_n3888# 0.009069f
C299 plus.n30 a_n2982_n3888# 0.460178f
C300 plus.n31 a_n2982_n3888# 0.009069f
C301 plus.n32 a_n2982_n3888# 0.459808f
C302 plus.n33 a_n2982_n3888# 0.52071f
C303 plus.n34 a_n2982_n3888# 0.039965f
C304 plus.t17 a_n2982_n3888# 1.19247f
C305 plus.n35 a_n2982_n3888# 0.039965f
C306 plus.t16 a_n2982_n3888# 1.19247f
C307 plus.t0 a_n2982_n3888# 1.19247f
C308 plus.n36 a_n2982_n3888# 0.460178f
C309 plus.n37 a_n2982_n3888# 0.039965f
C310 plus.t9 a_n2982_n3888# 1.19247f
C311 plus.t8 a_n2982_n3888# 1.19247f
C312 plus.n38 a_n2982_n3888# 0.460178f
C313 plus.n39 a_n2982_n3888# 0.039965f
C314 plus.t14 a_n2982_n3888# 1.19247f
C315 plus.t13 a_n2982_n3888# 1.19247f
C316 plus.n40 a_n2982_n3888# 0.460178f
C317 plus.n41 a_n2982_n3888# 0.039965f
C318 plus.t18 a_n2982_n3888# 1.19247f
C319 plus.t3 a_n2982_n3888# 1.19247f
C320 plus.n42 a_n2982_n3888# 0.466862f
C321 plus.t2 a_n2982_n3888# 1.21203f
C322 plus.n43 a_n2982_n3888# 0.443487f
C323 plus.n44 a_n2982_n3888# 0.170587f
C324 plus.n45 a_n2982_n3888# 0.009069f
C325 plus.n46 a_n2982_n3888# 0.460178f
C326 plus.n47 a_n2982_n3888# 0.009069f
C327 plus.n48 a_n2982_n3888# 0.039965f
C328 plus.n49 a_n2982_n3888# 0.039965f
C329 plus.n50 a_n2982_n3888# 0.039965f
C330 plus.n51 a_n2982_n3888# 0.009069f
C331 plus.n52 a_n2982_n3888# 0.460178f
C332 plus.n53 a_n2982_n3888# 0.009069f
C333 plus.n54 a_n2982_n3888# 0.039965f
C334 plus.n55 a_n2982_n3888# 0.039965f
C335 plus.n56 a_n2982_n3888# 0.039965f
C336 plus.n57 a_n2982_n3888# 0.009069f
C337 plus.n58 a_n2982_n3888# 0.460178f
C338 plus.n59 a_n2982_n3888# 0.009069f
C339 plus.n60 a_n2982_n3888# 0.039965f
C340 plus.n61 a_n2982_n3888# 0.039965f
C341 plus.n62 a_n2982_n3888# 0.039965f
C342 plus.n63 a_n2982_n3888# 0.009069f
C343 plus.n64 a_n2982_n3888# 0.460178f
C344 plus.n65 a_n2982_n3888# 0.009069f
C345 plus.n66 a_n2982_n3888# 0.459808f
C346 plus.n67 a_n2982_n3888# 1.52641f
.ends

