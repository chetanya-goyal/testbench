* NGSPICE file created from diffpair574.ext - technology: sky130A

.subckt diffpair574 minus drain_right drain_left source plus
X0 drain_left.t9 plus.t0 source.t13 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X1 drain_left.t8 plus.t1 source.t19 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X2 a_n1352_n4888# a_n1352_n4888# a_n1352_n4888# a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.2
X3 drain_right.t9 minus.t0 source.t6 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X4 source.t11 plus.t2 drain_left.t7 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X5 source.t12 plus.t3 drain_left.t6 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X6 drain_right.t8 minus.t1 source.t4 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X7 drain_right.t7 minus.t2 source.t9 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X8 source.t1 minus.t3 drain_right.t6 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X9 source.t5 minus.t4 drain_right.t5 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X10 source.t8 minus.t5 drain_right.t4 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X11 drain_left.t5 plus.t4 source.t10 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X12 drain_right.t3 minus.t6 source.t7 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X13 drain_right.t2 minus.t7 source.t0 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X14 drain_right.t1 minus.t8 source.t3 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X15 a_n1352_n4888# a_n1352_n4888# a_n1352_n4888# a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X16 drain_left.t4 plus.t5 source.t17 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X17 source.t16 plus.t6 drain_left.t3 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X18 a_n1352_n4888# a_n1352_n4888# a_n1352_n4888# a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X19 source.t2 minus.t9 drain_right.t0 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X20 source.t15 plus.t7 drain_left.t2 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X21 a_n1352_n4888# a_n1352_n4888# a_n1352_n4888# a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X22 drain_left.t1 plus.t8 source.t14 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X23 drain_left.t0 plus.t9 source.t18 a_n1352_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
R0 plus.n2 plus.t4 2611.93
R1 plus.n8 plus.t5 2611.93
R2 plus.n12 plus.t0 2611.93
R3 plus.n18 plus.t9 2611.93
R4 plus.n1 plus.t3 2566.65
R5 plus.n5 plus.t8 2566.65
R6 plus.n7 plus.t6 2566.65
R7 plus.n11 plus.t2 2566.65
R8 plus.n15 plus.t1 2566.65
R9 plus.n17 plus.t7 2566.65
R10 plus.n3 plus.n2 161.489
R11 plus.n13 plus.n12 161.489
R12 plus.n4 plus.n3 161.3
R13 plus.n6 plus.n0 161.3
R14 plus.n9 plus.n8 161.3
R15 plus.n14 plus.n13 161.3
R16 plus.n16 plus.n10 161.3
R17 plus.n19 plus.n18 161.3
R18 plus.n4 plus.n1 40.8975
R19 plus.n7 plus.n6 40.8975
R20 plus.n17 plus.n16 40.8975
R21 plus.n14 plus.n11 40.8975
R22 plus.n5 plus.n4 36.5157
R23 plus.n6 plus.n5 36.5157
R24 plus.n16 plus.n15 36.5157
R25 plus.n15 plus.n14 36.5157
R26 plus.n2 plus.n1 32.1338
R27 plus.n8 plus.n7 32.1338
R28 plus.n18 plus.n17 32.1338
R29 plus.n12 plus.n11 32.1338
R30 plus plus.n19 31.1032
R31 plus plus.n9 15.1236
R32 plus.n3 plus.n0 0.189894
R33 plus.n9 plus.n0 0.189894
R34 plus.n19 plus.n10 0.189894
R35 plus.n13 plus.n10 0.189894
R36 source.n0 source.t17 44.1297
R37 source.n5 source.t7 44.1296
R38 source.n19 source.t3 44.1295
R39 source.n14 source.t13 44.1295
R40 source.n2 source.n1 43.1397
R41 source.n4 source.n3 43.1397
R42 source.n7 source.n6 43.1397
R43 source.n9 source.n8 43.1397
R44 source.n18 source.n17 43.1396
R45 source.n16 source.n15 43.1396
R46 source.n13 source.n12 43.1396
R47 source.n11 source.n10 43.1396
R48 source.n11 source.n9 28.2621
R49 source.n20 source.n0 22.3138
R50 source.n20 source.n19 5.49188
R51 source.n17 source.t4 0.9905
R52 source.n17 source.t5 0.9905
R53 source.n15 source.t9 0.9905
R54 source.n15 source.t8 0.9905
R55 source.n12 source.t19 0.9905
R56 source.n12 source.t11 0.9905
R57 source.n10 source.t18 0.9905
R58 source.n10 source.t15 0.9905
R59 source.n1 source.t14 0.9905
R60 source.n1 source.t16 0.9905
R61 source.n3 source.t10 0.9905
R62 source.n3 source.t12 0.9905
R63 source.n6 source.t6 0.9905
R64 source.n6 source.t1 0.9905
R65 source.n8 source.t0 0.9905
R66 source.n8 source.t2 0.9905
R67 source.n5 source.n4 0.698776
R68 source.n16 source.n14 0.698776
R69 source.n9 source.n7 0.457397
R70 source.n7 source.n5 0.457397
R71 source.n4 source.n2 0.457397
R72 source.n2 source.n0 0.457397
R73 source.n13 source.n11 0.457397
R74 source.n14 source.n13 0.457397
R75 source.n18 source.n16 0.457397
R76 source.n19 source.n18 0.457397
R77 source source.n20 0.188
R78 drain_left.n5 drain_left.t5 61.2653
R79 drain_left.n1 drain_left.t0 61.2652
R80 drain_left.n3 drain_left.n2 60.1057
R81 drain_left.n7 drain_left.n6 59.8185
R82 drain_left.n5 drain_left.n4 59.8185
R83 drain_left.n1 drain_left.n0 59.8184
R84 drain_left drain_left.n3 35.3695
R85 drain_left drain_left.n7 6.11011
R86 drain_left.n2 drain_left.t7 0.9905
R87 drain_left.n2 drain_left.t9 0.9905
R88 drain_left.n0 drain_left.t2 0.9905
R89 drain_left.n0 drain_left.t8 0.9905
R90 drain_left.n6 drain_left.t3 0.9905
R91 drain_left.n6 drain_left.t4 0.9905
R92 drain_left.n4 drain_left.t6 0.9905
R93 drain_left.n4 drain_left.t1 0.9905
R94 drain_left.n7 drain_left.n5 0.457397
R95 drain_left.n3 drain_left.n1 0.0593781
R96 minus.n8 minus.t7 2611.93
R97 minus.n2 minus.t6 2611.93
R98 minus.n18 minus.t8 2611.93
R99 minus.n12 minus.t2 2611.93
R100 minus.n7 minus.t9 2566.65
R101 minus.n5 minus.t0 2566.65
R102 minus.n1 minus.t3 2566.65
R103 minus.n17 minus.t4 2566.65
R104 minus.n15 minus.t1 2566.65
R105 minus.n11 minus.t5 2566.65
R106 minus.n3 minus.n2 161.489
R107 minus.n13 minus.n12 161.489
R108 minus.n9 minus.n8 161.3
R109 minus.n6 minus.n0 161.3
R110 minus.n4 minus.n3 161.3
R111 minus.n19 minus.n18 161.3
R112 minus.n16 minus.n10 161.3
R113 minus.n14 minus.n13 161.3
R114 minus.n7 minus.n6 40.8975
R115 minus.n4 minus.n1 40.8975
R116 minus.n14 minus.n11 40.8975
R117 minus.n17 minus.n16 40.8975
R118 minus.n20 minus.n9 40.2524
R119 minus.n6 minus.n5 36.5157
R120 minus.n5 minus.n4 36.5157
R121 minus.n15 minus.n14 36.5157
R122 minus.n16 minus.n15 36.5157
R123 minus.n8 minus.n7 32.1338
R124 minus.n2 minus.n1 32.1338
R125 minus.n12 minus.n11 32.1338
R126 minus.n18 minus.n17 32.1338
R127 minus.n20 minus.n19 6.44936
R128 minus.n9 minus.n0 0.189894
R129 minus.n3 minus.n0 0.189894
R130 minus.n13 minus.n10 0.189894
R131 minus.n19 minus.n10 0.189894
R132 minus minus.n20 0.188
R133 drain_right.n1 drain_right.t7 61.2652
R134 drain_right.n7 drain_right.t2 60.8084
R135 drain_right.n6 drain_right.n4 60.2753
R136 drain_right.n3 drain_right.n2 60.1057
R137 drain_right.n6 drain_right.n5 59.8185
R138 drain_right.n1 drain_right.n0 59.8184
R139 drain_right drain_right.n3 34.8163
R140 drain_right drain_right.n7 5.88166
R141 drain_right.n2 drain_right.t5 0.9905
R142 drain_right.n2 drain_right.t1 0.9905
R143 drain_right.n0 drain_right.t4 0.9905
R144 drain_right.n0 drain_right.t8 0.9905
R145 drain_right.n4 drain_right.t6 0.9905
R146 drain_right.n4 drain_right.t3 0.9905
R147 drain_right.n5 drain_right.t0 0.9905
R148 drain_right.n5 drain_right.t9 0.9905
R149 drain_right.n7 drain_right.n6 0.457397
R150 drain_right.n3 drain_right.n1 0.0593781
C0 drain_left minus 0.170748f
C1 drain_right minus 4.87423f
C2 drain_left source 40.1497f
C3 drain_right source 40.130398f
C4 drain_left plus 4.997221f
C5 drain_right plus 0.285178f
C6 drain_left drain_right 0.666424f
C7 minus source 4.04997f
C8 plus minus 6.32203f
C9 plus source 4.06518f
C10 drain_right a_n1352_n4888# 9.585141f
C11 drain_left a_n1352_n4888# 9.80033f
C12 source a_n1352_n4888# 8.697069f
C13 minus a_n1352_n4888# 5.752514f
C14 plus a_n1352_n4888# 8.45726f
C15 drain_right.t7 a_n1352_n4888# 6.226f
C16 drain_right.t4 a_n1352_n4888# 0.532197f
C17 drain_right.t8 a_n1352_n4888# 0.532197f
C18 drain_right.n0 a_n1352_n4888# 4.86546f
C19 drain_right.n1 a_n1352_n4888# 0.791581f
C20 drain_right.t5 a_n1352_n4888# 0.532197f
C21 drain_right.t1 a_n1352_n4888# 0.532197f
C22 drain_right.n2 a_n1352_n4888# 4.86728f
C23 drain_right.n3 a_n1352_n4888# 2.43114f
C24 drain_right.t6 a_n1352_n4888# 0.532197f
C25 drain_right.t3 a_n1352_n4888# 0.532197f
C26 drain_right.n4 a_n1352_n4888# 4.86846f
C27 drain_right.t0 a_n1352_n4888# 0.532197f
C28 drain_right.t9 a_n1352_n4888# 0.532197f
C29 drain_right.n5 a_n1352_n4888# 4.86545f
C30 drain_right.n6 a_n1352_n4888# 0.777181f
C31 drain_right.t2 a_n1352_n4888# 6.22273f
C32 drain_right.n7 a_n1352_n4888# 0.715162f
C33 minus.n0 a_n1352_n4888# 0.057735f
C34 minus.t7 a_n1352_n4888# 0.65474f
C35 minus.t9 a_n1352_n4888# 0.650442f
C36 minus.t0 a_n1352_n4888# 0.650442f
C37 minus.t3 a_n1352_n4888# 0.650442f
C38 minus.n1 a_n1352_n4888# 0.247556f
C39 minus.t6 a_n1352_n4888# 0.65474f
C40 minus.n2 a_n1352_n4888# 0.263916f
C41 minus.n3 a_n1352_n4888# 0.12678f
C42 minus.n4 a_n1352_n4888# 0.020221f
C43 minus.n5 a_n1352_n4888# 0.247556f
C44 minus.n6 a_n1352_n4888# 0.020221f
C45 minus.n7 a_n1352_n4888# 0.247556f
C46 minus.n8 a_n1352_n4888# 0.263835f
C47 minus.n9 a_n1352_n4888# 2.39853f
C48 minus.n10 a_n1352_n4888# 0.057735f
C49 minus.t4 a_n1352_n4888# 0.650442f
C50 minus.t1 a_n1352_n4888# 0.650442f
C51 minus.t5 a_n1352_n4888# 0.650442f
C52 minus.n11 a_n1352_n4888# 0.247556f
C53 minus.t2 a_n1352_n4888# 0.65474f
C54 minus.n12 a_n1352_n4888# 0.263916f
C55 minus.n13 a_n1352_n4888# 0.12678f
C56 minus.n14 a_n1352_n4888# 0.020221f
C57 minus.n15 a_n1352_n4888# 0.247556f
C58 minus.n16 a_n1352_n4888# 0.020221f
C59 minus.n17 a_n1352_n4888# 0.247556f
C60 minus.t8 a_n1352_n4888# 0.65474f
C61 minus.n18 a_n1352_n4888# 0.263835f
C62 minus.n19 a_n1352_n4888# 0.370555f
C63 minus.n20 a_n1352_n4888# 2.88063f
C64 drain_left.t0 a_n1352_n4888# 6.22162f
C65 drain_left.t2 a_n1352_n4888# 0.531823f
C66 drain_left.t8 a_n1352_n4888# 0.531823f
C67 drain_left.n0 a_n1352_n4888# 4.86204f
C68 drain_left.n1 a_n1352_n4888# 0.791025f
C69 drain_left.t7 a_n1352_n4888# 0.531823f
C70 drain_left.t9 a_n1352_n4888# 0.531823f
C71 drain_left.n2 a_n1352_n4888# 4.86386f
C72 drain_left.n3 a_n1352_n4888# 2.5f
C73 drain_left.t5 a_n1352_n4888# 6.22165f
C74 drain_left.t6 a_n1352_n4888# 0.531823f
C75 drain_left.t1 a_n1352_n4888# 0.531823f
C76 drain_left.n4 a_n1352_n4888# 4.86203f
C77 drain_left.n5 a_n1352_n4888# 0.820914f
C78 drain_left.t3 a_n1352_n4888# 0.531823f
C79 drain_left.t4 a_n1352_n4888# 0.531823f
C80 drain_left.n6 a_n1352_n4888# 4.86203f
C81 drain_left.n7 a_n1352_n4888# 0.658436f
C82 source.t17 a_n1352_n4888# 6.14392f
C83 source.n0 a_n1352_n4888# 2.59832f
C84 source.t14 a_n1352_n4888# 0.537602f
C85 source.t16 a_n1352_n4888# 0.537602f
C86 source.n1 a_n1352_n4888# 4.80639f
C87 source.n2 a_n1352_n4888# 0.44945f
C88 source.t10 a_n1352_n4888# 0.537602f
C89 source.t12 a_n1352_n4888# 0.537602f
C90 source.n3 a_n1352_n4888# 4.80639f
C91 source.n4 a_n1352_n4888# 0.475906f
C92 source.t7 a_n1352_n4888# 6.14393f
C93 source.n5 a_n1352_n4888# 0.604552f
C94 source.t6 a_n1352_n4888# 0.537602f
C95 source.t1 a_n1352_n4888# 0.537602f
C96 source.n6 a_n1352_n4888# 4.80639f
C97 source.n7 a_n1352_n4888# 0.44945f
C98 source.t0 a_n1352_n4888# 0.537602f
C99 source.t2 a_n1352_n4888# 0.537602f
C100 source.n8 a_n1352_n4888# 4.80639f
C101 source.n9 a_n1352_n4888# 3.11855f
C102 source.t18 a_n1352_n4888# 0.537602f
C103 source.t15 a_n1352_n4888# 0.537602f
C104 source.n10 a_n1352_n4888# 4.8064f
C105 source.n11 a_n1352_n4888# 3.11854f
C106 source.t19 a_n1352_n4888# 0.537602f
C107 source.t11 a_n1352_n4888# 0.537602f
C108 source.n12 a_n1352_n4888# 4.8064f
C109 source.n13 a_n1352_n4888# 0.44944f
C110 source.t13 a_n1352_n4888# 6.1439f
C111 source.n14 a_n1352_n4888# 0.604586f
C112 source.t9 a_n1352_n4888# 0.537602f
C113 source.t8 a_n1352_n4888# 0.537602f
C114 source.n15 a_n1352_n4888# 4.8064f
C115 source.n16 a_n1352_n4888# 0.475897f
C116 source.t4 a_n1352_n4888# 0.537602f
C117 source.t5 a_n1352_n4888# 0.537602f
C118 source.n17 a_n1352_n4888# 4.8064f
C119 source.n18 a_n1352_n4888# 0.44944f
C120 source.t3 a_n1352_n4888# 6.1439f
C121 source.n19 a_n1352_n4888# 0.76399f
C122 source.n20 a_n1352_n4888# 3.05616f
C123 plus.n0 a_n1352_n4888# 0.058948f
C124 plus.t6 a_n1352_n4888# 0.664102f
C125 plus.t8 a_n1352_n4888# 0.664102f
C126 plus.t3 a_n1352_n4888# 0.664102f
C127 plus.n1 a_n1352_n4888# 0.252755f
C128 plus.t4 a_n1352_n4888# 0.66849f
C129 plus.n2 a_n1352_n4888# 0.269459f
C130 plus.n3 a_n1352_n4888# 0.129443f
C131 plus.n4 a_n1352_n4888# 0.020645f
C132 plus.n5 a_n1352_n4888# 0.252755f
C133 plus.n6 a_n1352_n4888# 0.020645f
C134 plus.n7 a_n1352_n4888# 0.252755f
C135 plus.t5 a_n1352_n4888# 0.66849f
C136 plus.n8 a_n1352_n4888# 0.269376f
C137 plus.n9 a_n1352_n4888# 0.888211f
C138 plus.n10 a_n1352_n4888# 0.058948f
C139 plus.t9 a_n1352_n4888# 0.66849f
C140 plus.t7 a_n1352_n4888# 0.664102f
C141 plus.t1 a_n1352_n4888# 0.664102f
C142 plus.t2 a_n1352_n4888# 0.664102f
C143 plus.n11 a_n1352_n4888# 0.252755f
C144 plus.t0 a_n1352_n4888# 0.66849f
C145 plus.n12 a_n1352_n4888# 0.269459f
C146 plus.n13 a_n1352_n4888# 0.129443f
C147 plus.n14 a_n1352_n4888# 0.020645f
C148 plus.n15 a_n1352_n4888# 0.252755f
C149 plus.n16 a_n1352_n4888# 0.020645f
C150 plus.n17 a_n1352_n4888# 0.252755f
C151 plus.n18 a_n1352_n4888# 0.269376f
C152 plus.n19 a_n1352_n4888# 1.92212f
.ends

