* NGSPICE file created from diffpair633.ext - technology: sky130A

.subckt diffpair633 minus drain_right drain_left source plus
X0 a_n1846_n4888# a_n1846_n4888# a_n1846_n4888# a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.8
X1 drain_left.t7 plus.t0 source.t8 a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X2 source.t1 minus.t0 drain_right.t7 a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X3 a_n1846_n4888# a_n1846_n4888# a_n1846_n4888# a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X4 a_n1846_n4888# a_n1846_n4888# a_n1846_n4888# a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X5 drain_right.t6 minus.t1 source.t3 a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X6 source.t10 plus.t1 drain_left.t6 a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X7 drain_right.t5 minus.t2 source.t0 a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X8 source.t7 minus.t3 drain_right.t4 a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X9 source.t9 plus.t2 drain_left.t5 a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X10 drain_right.t3 minus.t4 source.t6 a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X11 drain_right.t2 minus.t5 source.t5 a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X12 source.t2 minus.t6 drain_right.t1 a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
X13 a_n1846_n4888# a_n1846_n4888# a_n1846_n4888# a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.8
X14 drain_left.t4 plus.t3 source.t14 a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.8
X15 source.t15 plus.t4 drain_left.t3 a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X16 drain_left.t2 plus.t5 source.t11 a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X17 drain_left.t1 plus.t6 source.t12 a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X18 source.t4 minus.t7 drain_right.t0 a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.8
X19 source.t13 plus.t7 drain_left.t0 a_n1846_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.8
R0 plus.n2 plus.t7 672.207
R1 plus.n10 plus.t0 672.207
R2 plus.n6 plus.t3 651.605
R3 plus.n4 plus.t4 651.605
R4 plus.n3 plus.t6 651.605
R5 plus.n14 plus.t1 651.605
R6 plus.n12 plus.t5 651.605
R7 plus.n11 plus.t2 651.605
R8 plus.n5 plus.n0 161.3
R9 plus.n7 plus.n6 161.3
R10 plus.n13 plus.n8 161.3
R11 plus.n15 plus.n14 161.3
R12 plus.n4 plus.n1 80.6037
R13 plus.n12 plus.n9 80.6037
R14 plus.n4 plus.n3 48.2005
R15 plus.n12 plus.n11 48.2005
R16 plus.n5 plus.n4 41.6278
R17 plus.n13 plus.n12 41.6278
R18 plus plus.n15 33.1771
R19 plus.n2 plus.n1 31.6158
R20 plus.n10 plus.n9 31.6158
R21 plus.n3 plus.n2 17.6494
R22 plus.n11 plus.n10 17.6494
R23 plus plus.n7 15.3263
R24 plus.n6 plus.n5 6.57323
R25 plus.n14 plus.n13 6.57323
R26 plus.n1 plus.n0 0.285035
R27 plus.n9 plus.n8 0.285035
R28 plus.n7 plus.n0 0.189894
R29 plus.n15 plus.n8 0.189894
R30 source.n0 source.t14 44.1297
R31 source.n3 source.t13 44.1296
R32 source.n4 source.t6 44.1296
R33 source.n7 source.t2 44.1296
R34 source.n15 source.t3 44.1295
R35 source.n12 source.t1 44.1295
R36 source.n11 source.t8 44.1295
R37 source.n8 source.t10 44.1295
R38 source.n2 source.n1 43.1397
R39 source.n6 source.n5 43.1397
R40 source.n14 source.n13 43.1396
R41 source.n10 source.n9 43.1396
R42 source.n8 source.n7 28.3225
R43 source.n16 source.n0 22.5725
R44 source.n16 source.n15 5.7505
R45 source.n13 source.t5 0.9905
R46 source.n13 source.t4 0.9905
R47 source.n9 source.t11 0.9905
R48 source.n9 source.t9 0.9905
R49 source.n1 source.t12 0.9905
R50 source.n1 source.t15 0.9905
R51 source.n5 source.t0 0.9905
R52 source.n5 source.t7 0.9905
R53 source.n7 source.n6 0.974638
R54 source.n6 source.n4 0.974638
R55 source.n3 source.n2 0.974638
R56 source.n2 source.n0 0.974638
R57 source.n10 source.n8 0.974638
R58 source.n11 source.n10 0.974638
R59 source.n14 source.n12 0.974638
R60 source.n15 source.n14 0.974638
R61 source.n4 source.n3 0.470328
R62 source.n12 source.n11 0.470328
R63 source source.n16 0.188
R64 drain_left.n5 drain_left.n3 60.7926
R65 drain_left.n2 drain_left.n1 60.2501
R66 drain_left.n2 drain_left.n0 60.2501
R67 drain_left.n5 drain_left.n4 59.8185
R68 drain_left drain_left.n2 36.8372
R69 drain_left drain_left.n5 6.62735
R70 drain_left.n1 drain_left.t5 0.9905
R71 drain_left.n1 drain_left.t7 0.9905
R72 drain_left.n0 drain_left.t6 0.9905
R73 drain_left.n0 drain_left.t2 0.9905
R74 drain_left.n4 drain_left.t3 0.9905
R75 drain_left.n4 drain_left.t4 0.9905
R76 drain_left.n3 drain_left.t0 0.9905
R77 drain_left.n3 drain_left.t1 0.9905
R78 minus.n2 minus.t4 672.207
R79 minus.n10 minus.t0 672.207
R80 minus.n1 minus.t3 651.605
R81 minus.n4 minus.t2 651.605
R82 minus.n6 minus.t6 651.605
R83 minus.n9 minus.t5 651.605
R84 minus.n12 minus.t7 651.605
R85 minus.n14 minus.t1 651.605
R86 minus.n7 minus.n6 161.3
R87 minus.n5 minus.n0 161.3
R88 minus.n15 minus.n14 161.3
R89 minus.n13 minus.n8 161.3
R90 minus.n4 minus.n3 80.6037
R91 minus.n12 minus.n11 80.6037
R92 minus.n4 minus.n1 48.2005
R93 minus.n12 minus.n9 48.2005
R94 minus.n16 minus.n7 42.3263
R95 minus.n5 minus.n4 41.6278
R96 minus.n13 minus.n12 41.6278
R97 minus.n3 minus.n2 31.6158
R98 minus.n11 minus.n10 31.6158
R99 minus.n2 minus.n1 17.6494
R100 minus.n10 minus.n9 17.6494
R101 minus.n16 minus.n15 6.65202
R102 minus.n6 minus.n5 6.57323
R103 minus.n14 minus.n13 6.57323
R104 minus.n3 minus.n0 0.285035
R105 minus.n11 minus.n8 0.285035
R106 minus.n7 minus.n0 0.189894
R107 minus.n15 minus.n8 0.189894
R108 minus minus.n16 0.188
R109 drain_right.n5 drain_right.n3 60.7926
R110 drain_right.n2 drain_right.n1 60.2501
R111 drain_right.n2 drain_right.n0 60.2501
R112 drain_right.n5 drain_right.n4 59.8185
R113 drain_right drain_right.n2 36.2839
R114 drain_right drain_right.n5 6.62735
R115 drain_right.n1 drain_right.t0 0.9905
R116 drain_right.n1 drain_right.t6 0.9905
R117 drain_right.n0 drain_right.t7 0.9905
R118 drain_right.n0 drain_right.t2 0.9905
R119 drain_right.n3 drain_right.t4 0.9905
R120 drain_right.n3 drain_right.t3 0.9905
R121 drain_right.n4 drain_right.t1 0.9905
R122 drain_right.n4 drain_right.t5 0.9905
C0 minus drain_left 0.17159f
C1 drain_right drain_left 0.873724f
C2 drain_left plus 9.76114f
C3 source drain_left 16.164501f
C4 minus drain_right 9.58189f
C5 minus plus 6.92473f
C6 source minus 9.05562f
C7 drain_right plus 0.333957f
C8 source drain_right 16.1668f
C9 source plus 9.069651f
C10 drain_right a_n1846_n4888# 7.21735f
C11 drain_left a_n1846_n4888# 7.48736f
C12 source a_n1846_n4888# 13.63161f
C13 minus a_n1846_n4888# 7.695901f
C14 plus a_n1846_n4888# 9.72678f
C15 drain_right.t7 a_n1846_n4888# 0.422192f
C16 drain_right.t2 a_n1846_n4888# 0.422192f
C17 drain_right.n0 a_n1846_n4888# 3.86235f
C18 drain_right.t0 a_n1846_n4888# 0.422192f
C19 drain_right.t6 a_n1846_n4888# 0.422192f
C20 drain_right.n1 a_n1846_n4888# 3.86235f
C21 drain_right.n2 a_n1846_n4888# 2.52042f
C22 drain_right.t4 a_n1846_n4888# 0.422192f
C23 drain_right.t3 a_n1846_n4888# 0.422192f
C24 drain_right.n3 a_n1846_n4888# 3.86624f
C25 drain_right.t1 a_n1846_n4888# 0.422192f
C26 drain_right.t5 a_n1846_n4888# 0.422192f
C27 drain_right.n4 a_n1846_n4888# 3.85977f
C28 drain_right.n5 a_n1846_n4888# 1.03008f
C29 minus.n0 a_n1846_n4888# 0.055211f
C30 minus.t3 a_n1846_n4888# 1.87475f
C31 minus.n1 a_n1846_n4888# 0.707536f
C32 minus.t2 a_n1846_n4888# 1.87475f
C33 minus.t4 a_n1846_n4888# 1.89617f
C34 minus.n2 a_n1846_n4888# 0.681099f
C35 minus.n3 a_n1846_n4888# 0.236808f
C36 minus.n4 a_n1846_n4888# 0.706862f
C37 minus.n5 a_n1846_n4888# 0.009389f
C38 minus.t6 a_n1846_n4888# 1.87475f
C39 minus.n6 a_n1846_n4888# 0.691351f
C40 minus.n7 a_n1846_n4888# 1.8575f
C41 minus.n8 a_n1846_n4888# 0.055211f
C42 minus.t5 a_n1846_n4888# 1.87475f
C43 minus.n9 a_n1846_n4888# 0.707536f
C44 minus.t0 a_n1846_n4888# 1.89617f
C45 minus.n10 a_n1846_n4888# 0.681099f
C46 minus.n11 a_n1846_n4888# 0.236808f
C47 minus.t7 a_n1846_n4888# 1.87475f
C48 minus.n12 a_n1846_n4888# 0.706862f
C49 minus.n13 a_n1846_n4888# 0.009389f
C50 minus.t1 a_n1846_n4888# 1.87475f
C51 minus.n14 a_n1846_n4888# 0.691351f
C52 minus.n15 a_n1846_n4888# 0.285217f
C53 minus.n16 a_n1846_n4888# 2.21276f
C54 drain_left.t6 a_n1846_n4888# 0.423749f
C55 drain_left.t2 a_n1846_n4888# 0.423749f
C56 drain_left.n0 a_n1846_n4888# 3.87658f
C57 drain_left.t5 a_n1846_n4888# 0.423749f
C58 drain_left.t7 a_n1846_n4888# 0.423749f
C59 drain_left.n1 a_n1846_n4888# 3.87658f
C60 drain_left.n2 a_n1846_n4888# 2.58554f
C61 drain_left.t0 a_n1846_n4888# 0.423749f
C62 drain_left.t1 a_n1846_n4888# 0.423749f
C63 drain_left.n3 a_n1846_n4888# 3.8805f
C64 drain_left.t3 a_n1846_n4888# 0.423749f
C65 drain_left.t4 a_n1846_n4888# 0.423749f
C66 drain_left.n4 a_n1846_n4888# 3.874f
C67 drain_left.n5 a_n1846_n4888# 1.03388f
C68 source.t14 a_n1846_n4888# 3.42391f
C69 source.n0 a_n1846_n4888# 1.49779f
C70 source.t12 a_n1846_n4888# 0.299597f
C71 source.t15 a_n1846_n4888# 0.299597f
C72 source.n1 a_n1846_n4888# 2.67853f
C73 source.n2 a_n1846_n4888# 0.313659f
C74 source.t13 a_n1846_n4888# 3.42392f
C75 source.n3 a_n1846_n4888# 0.354547f
C76 source.t6 a_n1846_n4888# 3.42392f
C77 source.n4 a_n1846_n4888# 0.354547f
C78 source.t0 a_n1846_n4888# 0.299597f
C79 source.t7 a_n1846_n4888# 0.299597f
C80 source.n5 a_n1846_n4888# 2.67853f
C81 source.n6 a_n1846_n4888# 0.313659f
C82 source.t2 a_n1846_n4888# 3.42392f
C83 source.n7 a_n1846_n4888# 1.84489f
C84 source.t10 a_n1846_n4888# 3.4239f
C85 source.n8 a_n1846_n4888# 1.84491f
C86 source.t11 a_n1846_n4888# 0.299597f
C87 source.t9 a_n1846_n4888# 0.299597f
C88 source.n9 a_n1846_n4888# 2.67853f
C89 source.n10 a_n1846_n4888# 0.313654f
C90 source.t8 a_n1846_n4888# 3.4239f
C91 source.n11 a_n1846_n4888# 0.354566f
C92 source.t1 a_n1846_n4888# 3.4239f
C93 source.n12 a_n1846_n4888# 0.354566f
C94 source.t5 a_n1846_n4888# 0.299597f
C95 source.t4 a_n1846_n4888# 0.299597f
C96 source.n13 a_n1846_n4888# 2.67853f
C97 source.n14 a_n1846_n4888# 0.313654f
C98 source.t3 a_n1846_n4888# 3.4239f
C99 source.n15 a_n1846_n4888# 0.482323f
C100 source.n16 a_n1846_n4888# 1.72317f
C101 plus.n0 a_n1846_n4888# 0.055825f
C102 plus.t3 a_n1846_n4888# 1.89559f
C103 plus.t4 a_n1846_n4888# 1.89559f
C104 plus.n1 a_n1846_n4888# 0.239441f
C105 plus.t6 a_n1846_n4888# 1.89559f
C106 plus.t7 a_n1846_n4888# 1.91725f
C107 plus.n2 a_n1846_n4888# 0.688671f
C108 plus.n3 a_n1846_n4888# 0.715402f
C109 plus.n4 a_n1846_n4888# 0.714721f
C110 plus.n5 a_n1846_n4888# 0.009493f
C111 plus.n6 a_n1846_n4888# 0.699037f
C112 plus.n7 a_n1846_n4888# 0.649834f
C113 plus.n8 a_n1846_n4888# 0.055825f
C114 plus.t1 a_n1846_n4888# 1.89559f
C115 plus.n9 a_n1846_n4888# 0.239441f
C116 plus.t5 a_n1846_n4888# 1.89559f
C117 plus.t0 a_n1846_n4888# 1.91725f
C118 plus.n10 a_n1846_n4888# 0.688671f
C119 plus.t2 a_n1846_n4888# 1.89559f
C120 plus.n11 a_n1846_n4888# 0.715402f
C121 plus.n12 a_n1846_n4888# 0.714721f
C122 plus.n13 a_n1846_n4888# 0.009493f
C123 plus.n14 a_n1846_n4888# 0.699037f
C124 plus.n15 a_n1846_n4888# 1.48842f
.ends

