* NGSPICE file created from diffpair93.ext - technology: sky130A

.subckt diffpair93 minus drain_right drain_left source plus
X0 drain_right.t7 minus.t0 source.t10 a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X1 source.t6 plus.t0 drain_left.t7 a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X2 drain_right.t6 minus.t1 source.t11 a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X3 source.t4 plus.t1 drain_left.t6 a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X4 a_n1246_n1288# a_n1246_n1288# a_n1246_n1288# a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.2
X5 drain_left.t5 plus.t2 source.t5 a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X6 a_n1246_n1288# a_n1246_n1288# a_n1246_n1288# a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X7 source.t9 minus.t2 drain_right.t5 a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X8 source.t2 plus.t3 drain_left.t4 a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X9 a_n1246_n1288# a_n1246_n1288# a_n1246_n1288# a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X10 source.t8 minus.t3 drain_right.t4 a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X11 drain_left.t3 plus.t4 source.t3 a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
X12 drain_right.t3 minus.t4 source.t14 a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X13 drain_left.t2 plus.t5 source.t7 a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X14 a_n1246_n1288# a_n1246_n1288# a_n1246_n1288# a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.2
X15 drain_right.t2 minus.t5 source.t12 a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X16 source.t13 minus.t6 drain_right.t1 a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X17 source.t15 minus.t7 drain_right.t0 a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.2
X18 drain_left.t1 plus.t6 source.t1 a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.2
X19 source.t0 plus.t7 drain_left.t0 a_n1246_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.2
R0 minus.n5 minus.t6 440.738
R1 minus.n1 minus.t4 440.738
R2 minus.n12 minus.t5 440.738
R3 minus.n8 minus.t7 440.738
R4 minus.n4 minus.t1 397.651
R5 minus.n2 minus.t2 397.651
R6 minus.n11 minus.t3 397.651
R7 minus.n9 minus.t0 397.651
R8 minus.n1 minus.n0 161.489
R9 minus.n8 minus.n7 161.489
R10 minus.n6 minus.n5 161.3
R11 minus.n3 minus.n0 161.3
R12 minus.n13 minus.n12 161.3
R13 minus.n10 minus.n7 161.3
R14 minus.n4 minus.n3 38.7066
R15 minus.n3 minus.n2 38.7066
R16 minus.n10 minus.n9 38.7066
R17 minus.n11 minus.n10 38.7066
R18 minus.n5 minus.n4 34.3247
R19 minus.n2 minus.n1 34.3247
R20 minus.n9 minus.n8 34.3247
R21 minus.n12 minus.n11 34.3247
R22 minus.n14 minus.n6 26.2088
R23 minus.n14 minus.n13 6.44368
R24 minus.n6 minus.n0 0.189894
R25 minus.n13 minus.n7 0.189894
R26 minus minus.n14 0.188
R27 source.n66 source.n64 289.615
R28 source.n56 source.n54 289.615
R29 source.n48 source.n46 289.615
R30 source.n38 source.n36 289.615
R31 source.n2 source.n0 289.615
R32 source.n12 source.n10 289.615
R33 source.n20 source.n18 289.615
R34 source.n30 source.n28 289.615
R35 source.n67 source.n66 185
R36 source.n57 source.n56 185
R37 source.n49 source.n48 185
R38 source.n39 source.n38 185
R39 source.n3 source.n2 185
R40 source.n13 source.n12 185
R41 source.n21 source.n20 185
R42 source.n31 source.n30 185
R43 source.t12 source.n65 167.117
R44 source.t15 source.n55 167.117
R45 source.t1 source.n47 167.117
R46 source.t6 source.n37 167.117
R47 source.t7 source.n1 167.117
R48 source.t2 source.n11 167.117
R49 source.t14 source.n19 167.117
R50 source.t13 source.n29 167.117
R51 source.n9 source.n8 84.1169
R52 source.n27 source.n26 84.1169
R53 source.n63 source.n62 84.1168
R54 source.n45 source.n44 84.1168
R55 source.n66 source.t12 52.3082
R56 source.n56 source.t15 52.3082
R57 source.n48 source.t1 52.3082
R58 source.n38 source.t6 52.3082
R59 source.n2 source.t7 52.3082
R60 source.n12 source.t2 52.3082
R61 source.n20 source.t14 52.3082
R62 source.n30 source.t13 52.3082
R63 source.n71 source.n70 31.4096
R64 source.n61 source.n60 31.4096
R65 source.n53 source.n52 31.4096
R66 source.n43 source.n42 31.4096
R67 source.n7 source.n6 31.4096
R68 source.n17 source.n16 31.4096
R69 source.n25 source.n24 31.4096
R70 source.n35 source.n34 31.4096
R71 source.n43 source.n35 14.1689
R72 source.n62 source.t10 9.9005
R73 source.n62 source.t8 9.9005
R74 source.n44 source.t3 9.9005
R75 source.n44 source.t4 9.9005
R76 source.n8 source.t5 9.9005
R77 source.n8 source.t0 9.9005
R78 source.n26 source.t11 9.9005
R79 source.n26 source.t9 9.9005
R80 source.n67 source.n65 9.71174
R81 source.n57 source.n55 9.71174
R82 source.n49 source.n47 9.71174
R83 source.n39 source.n37 9.71174
R84 source.n3 source.n1 9.71174
R85 source.n13 source.n11 9.71174
R86 source.n21 source.n19 9.71174
R87 source.n31 source.n29 9.71174
R88 source.n70 source.n69 9.45567
R89 source.n60 source.n59 9.45567
R90 source.n52 source.n51 9.45567
R91 source.n42 source.n41 9.45567
R92 source.n6 source.n5 9.45567
R93 source.n16 source.n15 9.45567
R94 source.n24 source.n23 9.45567
R95 source.n34 source.n33 9.45567
R96 source.n69 source.n68 9.3005
R97 source.n59 source.n58 9.3005
R98 source.n51 source.n50 9.3005
R99 source.n41 source.n40 9.3005
R100 source.n5 source.n4 9.3005
R101 source.n15 source.n14 9.3005
R102 source.n23 source.n22 9.3005
R103 source.n33 source.n32 9.3005
R104 source.n72 source.n7 8.67749
R105 source.n70 source.n64 8.14595
R106 source.n60 source.n54 8.14595
R107 source.n52 source.n46 8.14595
R108 source.n42 source.n36 8.14595
R109 source.n6 source.n0 8.14595
R110 source.n16 source.n10 8.14595
R111 source.n24 source.n18 8.14595
R112 source.n34 source.n28 8.14595
R113 source.n68 source.n67 7.3702
R114 source.n58 source.n57 7.3702
R115 source.n50 source.n49 7.3702
R116 source.n40 source.n39 7.3702
R117 source.n4 source.n3 7.3702
R118 source.n14 source.n13 7.3702
R119 source.n22 source.n21 7.3702
R120 source.n32 source.n31 7.3702
R121 source.n68 source.n64 5.81868
R122 source.n58 source.n54 5.81868
R123 source.n50 source.n46 5.81868
R124 source.n40 source.n36 5.81868
R125 source.n4 source.n0 5.81868
R126 source.n14 source.n10 5.81868
R127 source.n22 source.n18 5.81868
R128 source.n32 source.n28 5.81868
R129 source.n72 source.n71 5.49188
R130 source.n69 source.n65 3.44771
R131 source.n59 source.n55 3.44771
R132 source.n51 source.n47 3.44771
R133 source.n41 source.n37 3.44771
R134 source.n5 source.n1 3.44771
R135 source.n15 source.n11 3.44771
R136 source.n23 source.n19 3.44771
R137 source.n33 source.n29 3.44771
R138 source.n25 source.n17 0.470328
R139 source.n61 source.n53 0.470328
R140 source.n35 source.n27 0.457397
R141 source.n27 source.n25 0.457397
R142 source.n17 source.n9 0.457397
R143 source.n9 source.n7 0.457397
R144 source.n45 source.n43 0.457397
R145 source.n53 source.n45 0.457397
R146 source.n63 source.n61 0.457397
R147 source.n71 source.n63 0.457397
R148 source source.n72 0.188
R149 drain_right.n5 drain_right.n3 101.252
R150 drain_right.n2 drain_right.n1 100.969
R151 drain_right.n2 drain_right.n0 100.969
R152 drain_right.n5 drain_right.n4 100.796
R153 drain_right drain_right.n2 20.8372
R154 drain_right.n1 drain_right.t4 9.9005
R155 drain_right.n1 drain_right.t2 9.9005
R156 drain_right.n0 drain_right.t0 9.9005
R157 drain_right.n0 drain_right.t7 9.9005
R158 drain_right.n3 drain_right.t5 9.9005
R159 drain_right.n3 drain_right.t3 9.9005
R160 drain_right.n4 drain_right.t1 9.9005
R161 drain_right.n4 drain_right.t6 9.9005
R162 drain_right drain_right.n5 6.11011
R163 plus.n1 plus.t3 440.738
R164 plus.n5 plus.t5 440.738
R165 plus.n8 plus.t6 440.738
R166 plus.n12 plus.t0 440.738
R167 plus.n2 plus.t2 397.651
R168 plus.n4 plus.t7 397.651
R169 plus.n9 plus.t1 397.651
R170 plus.n11 plus.t4 397.651
R171 plus.n1 plus.n0 161.489
R172 plus.n8 plus.n7 161.489
R173 plus.n3 plus.n0 161.3
R174 plus.n6 plus.n5 161.3
R175 plus.n10 plus.n7 161.3
R176 plus.n13 plus.n12 161.3
R177 plus.n3 plus.n2 38.7066
R178 plus.n4 plus.n3 38.7066
R179 plus.n11 plus.n10 38.7066
R180 plus.n10 plus.n9 38.7066
R181 plus.n2 plus.n1 34.3247
R182 plus.n5 plus.n4 34.3247
R183 plus.n12 plus.n11 34.3247
R184 plus.n9 plus.n8 34.3247
R185 plus plus.n13 23.8778
R186 plus plus.n6 8.29974
R187 plus.n6 plus.n0 0.189894
R188 plus.n13 plus.n7 0.189894
R189 drain_left.n5 drain_left.n3 101.252
R190 drain_left.n2 drain_left.n1 100.969
R191 drain_left.n2 drain_left.n0 100.969
R192 drain_left.n5 drain_left.n4 100.796
R193 drain_left drain_left.n2 21.3905
R194 drain_left.n1 drain_left.t6 9.9005
R195 drain_left.n1 drain_left.t1 9.9005
R196 drain_left.n0 drain_left.t7 9.9005
R197 drain_left.n0 drain_left.t3 9.9005
R198 drain_left.n4 drain_left.t0 9.9005
R199 drain_left.n4 drain_left.t2 9.9005
R200 drain_left.n3 drain_left.t4 9.9005
R201 drain_left.n3 drain_left.t5 9.9005
R202 drain_left drain_left.n5 6.11011
C0 source drain_left 4.74531f
C1 minus drain_right 0.72879f
C2 plus source 0.766089f
C3 plus drain_left 0.845608f
C4 drain_right source 4.74389f
C5 drain_right drain_left 0.58123f
C6 plus drain_right 0.27616f
C7 minus source 0.752126f
C8 minus drain_left 0.175947f
C9 plus minus 2.86409f
C10 drain_right a_n1246_n1288# 3.13501f
C11 drain_left a_n1246_n1288# 3.28964f
C12 source a_n1246_n1288# 2.828752f
C13 minus a_n1246_n1288# 4.003915f
C14 plus a_n1246_n1288# 4.767689f
C15 drain_left.t7 a_n1246_n1288# 0.042668f
C16 drain_left.t3 a_n1246_n1288# 0.042668f
C17 drain_left.n0 a_n1246_n1288# 0.268527f
C18 drain_left.t6 a_n1246_n1288# 0.042668f
C19 drain_left.t1 a_n1246_n1288# 0.042668f
C20 drain_left.n1 a_n1246_n1288# 0.268527f
C21 drain_left.n2 a_n1246_n1288# 1.15563f
C22 drain_left.t4 a_n1246_n1288# 0.042668f
C23 drain_left.t5 a_n1246_n1288# 0.042668f
C24 drain_left.n3 a_n1246_n1288# 0.269395f
C25 drain_left.t0 a_n1246_n1288# 0.042668f
C26 drain_left.t2 a_n1246_n1288# 0.042668f
C27 drain_left.n4 a_n1246_n1288# 0.268055f
C28 drain_left.n5 a_n1246_n1288# 0.802731f
C29 plus.n0 a_n1246_n1288# 0.085312f
C30 plus.t7 a_n1246_n1288# 0.046117f
C31 plus.t2 a_n1246_n1288# 0.046117f
C32 plus.t3 a_n1246_n1288# 0.049648f
C33 plus.n1 a_n1246_n1288# 0.04636f
C34 plus.n2 a_n1246_n1288# 0.036235f
C35 plus.n3 a_n1246_n1288# 0.013722f
C36 plus.n4 a_n1246_n1288# 0.036235f
C37 plus.t5 a_n1246_n1288# 0.049648f
C38 plus.n5 a_n1246_n1288# 0.046306f
C39 plus.n6 a_n1246_n1288# 0.274608f
C40 plus.n7 a_n1246_n1288# 0.085312f
C41 plus.t0 a_n1246_n1288# 0.049648f
C42 plus.t4 a_n1246_n1288# 0.046117f
C43 plus.t1 a_n1246_n1288# 0.046117f
C44 plus.t6 a_n1246_n1288# 0.049648f
C45 plus.n8 a_n1246_n1288# 0.04636f
C46 plus.n9 a_n1246_n1288# 0.036235f
C47 plus.n10 a_n1246_n1288# 0.013722f
C48 plus.n11 a_n1246_n1288# 0.036235f
C49 plus.n12 a_n1246_n1288# 0.046306f
C50 plus.n13 a_n1246_n1288# 0.769515f
C51 drain_right.t0 a_n1246_n1288# 0.043649f
C52 drain_right.t7 a_n1246_n1288# 0.043649f
C53 drain_right.n0 a_n1246_n1288# 0.274699f
C54 drain_right.t4 a_n1246_n1288# 0.043649f
C55 drain_right.t2 a_n1246_n1288# 0.043649f
C56 drain_right.n1 a_n1246_n1288# 0.274699f
C57 drain_right.n2 a_n1246_n1288# 1.12776f
C58 drain_right.t5 a_n1246_n1288# 0.043649f
C59 drain_right.t3 a_n1246_n1288# 0.043649f
C60 drain_right.n3 a_n1246_n1288# 0.275588f
C61 drain_right.t1 a_n1246_n1288# 0.043649f
C62 drain_right.t6 a_n1246_n1288# 0.043649f
C63 drain_right.n4 a_n1246_n1288# 0.274217f
C64 drain_right.n5 a_n1246_n1288# 0.821183f
C65 source.n0 a_n1246_n1288# 0.0381f
C66 source.n1 a_n1246_n1288# 0.084302f
C67 source.t7 a_n1246_n1288# 0.063264f
C68 source.n2 a_n1246_n1288# 0.065978f
C69 source.n3 a_n1246_n1288# 0.021269f
C70 source.n4 a_n1246_n1288# 0.014027f
C71 source.n5 a_n1246_n1288# 0.185822f
C72 source.n6 a_n1246_n1288# 0.041767f
C73 source.n7 a_n1246_n1288# 0.381233f
C74 source.t5 a_n1246_n1288# 0.041256f
C75 source.t0 a_n1246_n1288# 0.041256f
C76 source.n8 a_n1246_n1288# 0.220556f
C77 source.n9 a_n1246_n1288# 0.279809f
C78 source.n10 a_n1246_n1288# 0.0381f
C79 source.n11 a_n1246_n1288# 0.084302f
C80 source.t2 a_n1246_n1288# 0.063264f
C81 source.n12 a_n1246_n1288# 0.065978f
C82 source.n13 a_n1246_n1288# 0.021269f
C83 source.n14 a_n1246_n1288# 0.014027f
C84 source.n15 a_n1246_n1288# 0.185822f
C85 source.n16 a_n1246_n1288# 0.041767f
C86 source.n17 a_n1246_n1288# 0.09944f
C87 source.n18 a_n1246_n1288# 0.0381f
C88 source.n19 a_n1246_n1288# 0.084302f
C89 source.t14 a_n1246_n1288# 0.063264f
C90 source.n20 a_n1246_n1288# 0.065978f
C91 source.n21 a_n1246_n1288# 0.021269f
C92 source.n22 a_n1246_n1288# 0.014027f
C93 source.n23 a_n1246_n1288# 0.185822f
C94 source.n24 a_n1246_n1288# 0.041767f
C95 source.n25 a_n1246_n1288# 0.09944f
C96 source.t11 a_n1246_n1288# 0.041256f
C97 source.t9 a_n1246_n1288# 0.041256f
C98 source.n26 a_n1246_n1288# 0.220556f
C99 source.n27 a_n1246_n1288# 0.279809f
C100 source.n28 a_n1246_n1288# 0.0381f
C101 source.n29 a_n1246_n1288# 0.084302f
C102 source.t13 a_n1246_n1288# 0.063264f
C103 source.n30 a_n1246_n1288# 0.065978f
C104 source.n31 a_n1246_n1288# 0.021269f
C105 source.n32 a_n1246_n1288# 0.014027f
C106 source.n33 a_n1246_n1288# 0.185822f
C107 source.n34 a_n1246_n1288# 0.041767f
C108 source.n35 a_n1246_n1288# 0.622995f
C109 source.n36 a_n1246_n1288# 0.0381f
C110 source.n37 a_n1246_n1288# 0.084302f
C111 source.t6 a_n1246_n1288# 0.063264f
C112 source.n38 a_n1246_n1288# 0.065978f
C113 source.n39 a_n1246_n1288# 0.021269f
C114 source.n40 a_n1246_n1288# 0.014027f
C115 source.n41 a_n1246_n1288# 0.185822f
C116 source.n42 a_n1246_n1288# 0.041767f
C117 source.n43 a_n1246_n1288# 0.622995f
C118 source.t3 a_n1246_n1288# 0.041256f
C119 source.t4 a_n1246_n1288# 0.041256f
C120 source.n44 a_n1246_n1288# 0.220554f
C121 source.n45 a_n1246_n1288# 0.27981f
C122 source.n46 a_n1246_n1288# 0.0381f
C123 source.n47 a_n1246_n1288# 0.084302f
C124 source.t1 a_n1246_n1288# 0.063264f
C125 source.n48 a_n1246_n1288# 0.065978f
C126 source.n49 a_n1246_n1288# 0.021269f
C127 source.n50 a_n1246_n1288# 0.014027f
C128 source.n51 a_n1246_n1288# 0.185822f
C129 source.n52 a_n1246_n1288# 0.041767f
C130 source.n53 a_n1246_n1288# 0.09944f
C131 source.n54 a_n1246_n1288# 0.0381f
C132 source.n55 a_n1246_n1288# 0.084302f
C133 source.t15 a_n1246_n1288# 0.063264f
C134 source.n56 a_n1246_n1288# 0.065978f
C135 source.n57 a_n1246_n1288# 0.021269f
C136 source.n58 a_n1246_n1288# 0.014027f
C137 source.n59 a_n1246_n1288# 0.185822f
C138 source.n60 a_n1246_n1288# 0.041767f
C139 source.n61 a_n1246_n1288# 0.09944f
C140 source.t10 a_n1246_n1288# 0.041256f
C141 source.t8 a_n1246_n1288# 0.041256f
C142 source.n62 a_n1246_n1288# 0.220554f
C143 source.n63 a_n1246_n1288# 0.27981f
C144 source.n64 a_n1246_n1288# 0.0381f
C145 source.n65 a_n1246_n1288# 0.084302f
C146 source.t12 a_n1246_n1288# 0.063264f
C147 source.n66 a_n1246_n1288# 0.065978f
C148 source.n67 a_n1246_n1288# 0.021269f
C149 source.n68 a_n1246_n1288# 0.014027f
C150 source.n69 a_n1246_n1288# 0.185822f
C151 source.n70 a_n1246_n1288# 0.041767f
C152 source.n71 a_n1246_n1288# 0.240984f
C153 source.n72 a_n1246_n1288# 0.642341f
C154 minus.n0 a_n1246_n1288# 0.083044f
C155 minus.t6 a_n1246_n1288# 0.048327f
C156 minus.t1 a_n1246_n1288# 0.044891f
C157 minus.t2 a_n1246_n1288# 0.044891f
C158 minus.t4 a_n1246_n1288# 0.048327f
C159 minus.n1 a_n1246_n1288# 0.045127f
C160 minus.n2 a_n1246_n1288# 0.035271f
C161 minus.n3 a_n1246_n1288# 0.013357f
C162 minus.n4 a_n1246_n1288# 0.035271f
C163 minus.n5 a_n1246_n1288# 0.045074f
C164 minus.n6 a_n1246_n1288# 0.77884f
C165 minus.n7 a_n1246_n1288# 0.083044f
C166 minus.t3 a_n1246_n1288# 0.044891f
C167 minus.t0 a_n1246_n1288# 0.044891f
C168 minus.t7 a_n1246_n1288# 0.048327f
C169 minus.n8 a_n1246_n1288# 0.045127f
C170 minus.n9 a_n1246_n1288# 0.035271f
C171 minus.n10 a_n1246_n1288# 0.013357f
C172 minus.n11 a_n1246_n1288# 0.035271f
C173 minus.t5 a_n1246_n1288# 0.048327f
C174 minus.n12 a_n1246_n1288# 0.045074f
C175 minus.n13 a_n1246_n1288# 0.244267f
C176 minus.n14 a_n1246_n1288# 0.96469f
.ends

