* NGSPICE file created from diffpair183.ext - technology: sky130A

.subckt diffpair183 minus drain_right drain_left source plus
X0 a_n1296_n1488# a_n1296_n1488# a_n1296_n1488# a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.25
X1 drain_left.t7 plus.t0 source.t6 a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X2 drain_left.t6 plus.t1 source.t7 a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X3 source.t14 minus.t0 drain_right.t7 a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X4 source.t3 minus.t1 drain_right.t6 a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X5 source.t8 plus.t2 drain_left.t5 a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X6 source.t13 plus.t3 drain_left.t4 a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X7 drain_left.t3 plus.t4 source.t10 a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X8 a_n1296_n1488# a_n1296_n1488# a_n1296_n1488# a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X9 a_n1296_n1488# a_n1296_n1488# a_n1296_n1488# a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X10 drain_left.t2 plus.t5 source.t11 a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X11 source.t9 plus.t6 drain_left.t1 a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X12 source.t12 plus.t7 drain_left.t0 a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
X13 drain_right.t5 minus.t2 source.t0 a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X14 drain_right.t4 minus.t3 source.t15 a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X15 drain_right.t3 minus.t4 source.t1 a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X16 a_n1296_n1488# a_n1296_n1488# a_n1296_n1488# a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.25
X17 drain_right.t2 minus.t5 source.t2 a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.25
X18 source.t5 minus.t6 drain_right.t1 a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.25
X19 source.t4 minus.t7 drain_right.t0 a_n1296_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.25
R0 plus.n1 plus.t2 468.562
R1 plus.n5 plus.t0 468.562
R2 plus.n8 plus.t4 468.562
R3 plus.n12 plus.t7 468.562
R4 plus.n2 plus.t1 414.521
R5 plus.n4 plus.t6 414.521
R6 plus.n9 plus.t3 414.521
R7 plus.n11 plus.t5 414.521
R8 plus.n1 plus.n0 161.489
R9 plus.n8 plus.n7 161.489
R10 plus.n3 plus.n0 161.3
R11 plus.n6 plus.n5 161.3
R12 plus.n10 plus.n7 161.3
R13 plus.n13 plus.n12 161.3
R14 plus.n3 plus.n2 42.3581
R15 plus.n4 plus.n3 42.3581
R16 plus.n11 plus.n10 42.3581
R17 plus.n10 plus.n9 42.3581
R18 plus.n2 plus.n1 30.6732
R19 plus.n5 plus.n4 30.6732
R20 plus.n12 plus.n11 30.6732
R21 plus.n9 plus.n8 30.6732
R22 plus plus.n13 24.5028
R23 plus plus.n6 8.73535
R24 plus.n6 plus.n0 0.189894
R25 plus.n13 plus.n7 0.189894
R26 source.n0 source.t6 69.6943
R27 source.n3 source.t8 69.6943
R28 source.n4 source.t15 69.6943
R29 source.n7 source.t14 69.6943
R30 source.n15 source.t2 69.6942
R31 source.n12 source.t4 69.6942
R32 source.n11 source.t10 69.6942
R33 source.n8 source.t12 69.6942
R34 source.n2 source.n1 63.0943
R35 source.n6 source.n5 63.0943
R36 source.n14 source.n13 63.0942
R37 source.n10 source.n9 63.0942
R38 source.n8 source.n7 14.9695
R39 source.n16 source.n0 9.45661
R40 source.n13 source.t1 6.6005
R41 source.n13 source.t5 6.6005
R42 source.n9 source.t11 6.6005
R43 source.n9 source.t13 6.6005
R44 source.n1 source.t7 6.6005
R45 source.n1 source.t9 6.6005
R46 source.n5 source.t0 6.6005
R47 source.n5 source.t3 6.6005
R48 source.n16 source.n15 5.51343
R49 source.n7 source.n6 0.5005
R50 source.n6 source.n4 0.5005
R51 source.n3 source.n2 0.5005
R52 source.n2 source.n0 0.5005
R53 source.n10 source.n8 0.5005
R54 source.n11 source.n10 0.5005
R55 source.n14 source.n12 0.5005
R56 source.n15 source.n14 0.5005
R57 source.n4 source.n3 0.470328
R58 source.n12 source.n11 0.470328
R59 source source.n16 0.188
R60 drain_left.n5 drain_left.n3 80.2731
R61 drain_left.n2 drain_left.n1 79.9677
R62 drain_left.n2 drain_left.n0 79.9677
R63 drain_left.n5 drain_left.n4 79.7731
R64 drain_left drain_left.n2 22.2989
R65 drain_left.n1 drain_left.t4 6.6005
R66 drain_left.n1 drain_left.t3 6.6005
R67 drain_left.n0 drain_left.t0 6.6005
R68 drain_left.n0 drain_left.t2 6.6005
R69 drain_left.n4 drain_left.t1 6.6005
R70 drain_left.n4 drain_left.t7 6.6005
R71 drain_left.n3 drain_left.t5 6.6005
R72 drain_left.n3 drain_left.t6 6.6005
R73 drain_left drain_left.n5 6.15322
R74 minus.n5 minus.t0 468.562
R75 minus.n1 minus.t3 468.562
R76 minus.n12 minus.t5 468.562
R77 minus.n8 minus.t7 468.562
R78 minus.n4 minus.t2 414.521
R79 minus.n2 minus.t1 414.521
R80 minus.n11 minus.t6 414.521
R81 minus.n9 minus.t4 414.521
R82 minus.n1 minus.n0 161.489
R83 minus.n8 minus.n7 161.489
R84 minus.n6 minus.n5 161.3
R85 minus.n3 minus.n0 161.3
R86 minus.n13 minus.n12 161.3
R87 minus.n10 minus.n7 161.3
R88 minus.n4 minus.n3 42.3581
R89 minus.n3 minus.n2 42.3581
R90 minus.n10 minus.n9 42.3581
R91 minus.n11 minus.n10 42.3581
R92 minus.n5 minus.n4 30.6732
R93 minus.n2 minus.n1 30.6732
R94 minus.n9 minus.n8 30.6732
R95 minus.n12 minus.n11 30.6732
R96 minus.n14 minus.n6 27.2126
R97 minus.n14 minus.n13 6.5005
R98 minus.n6 minus.n0 0.189894
R99 minus.n13 minus.n7 0.189894
R100 minus minus.n14 0.188
R101 drain_right.n5 drain_right.n3 80.2731
R102 drain_right.n2 drain_right.n1 79.9677
R103 drain_right.n2 drain_right.n0 79.9677
R104 drain_right.n5 drain_right.n4 79.7731
R105 drain_right drain_right.n2 21.7457
R106 drain_right.n1 drain_right.t1 6.6005
R107 drain_right.n1 drain_right.t2 6.6005
R108 drain_right.n0 drain_right.t0 6.6005
R109 drain_right.n0 drain_right.t3 6.6005
R110 drain_right.n3 drain_right.t6 6.6005
R111 drain_right.n3 drain_right.t4 6.6005
R112 drain_right.n4 drain_right.t7 6.6005
R113 drain_right.n4 drain_right.t5 6.6005
R114 drain_right drain_right.n5 6.15322
C0 drain_right plus 0.280621f
C1 drain_right minus 1.01365f
C2 source drain_left 5.8266f
C3 drain_left plus 1.13567f
C4 drain_left minus 0.175359f
C5 source plus 1.02114f
C6 source minus 1.00714f
C7 minus plus 3.10595f
C8 drain_right drain_left 0.605638f
C9 drain_right source 5.82547f
C10 drain_right a_n1296_n1488# 3.37659f
C11 drain_left a_n1296_n1488# 3.53871f
C12 source a_n1296_n1488# 3.419357f
C13 minus a_n1296_n1488# 4.269279f
C14 plus a_n1296_n1488# 5.002267f
C15 drain_right.t0 a_n1296_n1488# 0.063917f
C16 drain_right.t3 a_n1296_n1488# 0.063917f
C17 drain_right.n0 a_n1296_n1488# 0.46167f
C18 drain_right.t1 a_n1296_n1488# 0.063917f
C19 drain_right.t2 a_n1296_n1488# 0.063917f
C20 drain_right.n1 a_n1296_n1488# 0.46167f
C21 drain_right.n2 a_n1296_n1488# 1.19071f
C22 drain_right.t6 a_n1296_n1488# 0.063917f
C23 drain_right.t4 a_n1296_n1488# 0.063917f
C24 drain_right.n3 a_n1296_n1488# 0.462918f
C25 drain_right.t7 a_n1296_n1488# 0.063917f
C26 drain_right.t5 a_n1296_n1488# 0.063917f
C27 drain_right.n4 a_n1296_n1488# 0.460965f
C28 drain_right.n5 a_n1296_n1488# 0.836844f
C29 minus.n0 a_n1296_n1488# 0.078121f
C30 minus.t0 a_n1296_n1488# 0.079182f
C31 minus.t2 a_n1296_n1488# 0.073752f
C32 minus.t1 a_n1296_n1488# 0.073752f
C33 minus.t3 a_n1296_n1488# 0.079182f
C34 minus.n1 a_n1296_n1488# 0.054642f
C35 minus.n2 a_n1296_n1488# 0.044569f
C36 minus.n3 a_n1296_n1488# 0.01294f
C37 minus.n4 a_n1296_n1488# 0.044569f
C38 minus.n5 a_n1296_n1488# 0.05459f
C39 minus.n6 a_n1296_n1488# 0.744663f
C40 minus.n7 a_n1296_n1488# 0.078121f
C41 minus.t6 a_n1296_n1488# 0.073752f
C42 minus.t4 a_n1296_n1488# 0.073752f
C43 minus.t7 a_n1296_n1488# 0.079182f
C44 minus.n8 a_n1296_n1488# 0.054642f
C45 minus.n9 a_n1296_n1488# 0.044569f
C46 minus.n10 a_n1296_n1488# 0.01294f
C47 minus.n11 a_n1296_n1488# 0.044569f
C48 minus.t5 a_n1296_n1488# 0.079182f
C49 minus.n12 a_n1296_n1488# 0.05459f
C50 minus.n13 a_n1296_n1488# 0.222044f
C51 minus.n14 a_n1296_n1488# 0.920396f
C52 drain_left.t0 a_n1296_n1488# 0.062776f
C53 drain_left.t2 a_n1296_n1488# 0.062776f
C54 drain_left.n0 a_n1296_n1488# 0.453424f
C55 drain_left.t4 a_n1296_n1488# 0.062776f
C56 drain_left.t3 a_n1296_n1488# 0.062776f
C57 drain_left.n1 a_n1296_n1488# 0.453424f
C58 drain_left.n2 a_n1296_n1488# 1.22228f
C59 drain_left.t5 a_n1296_n1488# 0.062776f
C60 drain_left.t6 a_n1296_n1488# 0.062776f
C61 drain_left.n3 a_n1296_n1488# 0.454651f
C62 drain_left.t1 a_n1296_n1488# 0.062776f
C63 drain_left.t7 a_n1296_n1488# 0.062776f
C64 drain_left.n4 a_n1296_n1488# 0.452733f
C65 drain_left.n5 a_n1296_n1488# 0.821898f
C66 source.t6 a_n1296_n1488# 0.466686f
C67 source.n0 a_n1296_n1488# 0.630915f
C68 source.t7 a_n1296_n1488# 0.056201f
C69 source.t9 a_n1296_n1488# 0.056201f
C70 source.n1 a_n1296_n1488# 0.356349f
C71 source.n2 a_n1296_n1488# 0.282905f
C72 source.t8 a_n1296_n1488# 0.466686f
C73 source.n3 a_n1296_n1488# 0.323539f
C74 source.t15 a_n1296_n1488# 0.466686f
C75 source.n4 a_n1296_n1488# 0.323539f
C76 source.t0 a_n1296_n1488# 0.056201f
C77 source.t3 a_n1296_n1488# 0.056201f
C78 source.n5 a_n1296_n1488# 0.356349f
C79 source.n6 a_n1296_n1488# 0.282905f
C80 source.t14 a_n1296_n1488# 0.466686f
C81 source.n7 a_n1296_n1488# 0.877241f
C82 source.t12 a_n1296_n1488# 0.466683f
C83 source.n8 a_n1296_n1488# 0.877244f
C84 source.t11 a_n1296_n1488# 0.056201f
C85 source.t13 a_n1296_n1488# 0.056201f
C86 source.n9 a_n1296_n1488# 0.356346f
C87 source.n10 a_n1296_n1488# 0.282907f
C88 source.t10 a_n1296_n1488# 0.466683f
C89 source.n11 a_n1296_n1488# 0.323541f
C90 source.t4 a_n1296_n1488# 0.466683f
C91 source.n12 a_n1296_n1488# 0.323541f
C92 source.t1 a_n1296_n1488# 0.056201f
C93 source.t5 a_n1296_n1488# 0.056201f
C94 source.n13 a_n1296_n1488# 0.356346f
C95 source.n14 a_n1296_n1488# 0.282907f
C96 source.t2 a_n1296_n1488# 0.466683f
C97 source.n15 a_n1296_n1488# 0.45473f
C98 source.n16 a_n1296_n1488# 0.685702f
C99 plus.n0 a_n1296_n1488# 0.079891f
C100 plus.t6 a_n1296_n1488# 0.075423f
C101 plus.t1 a_n1296_n1488# 0.075423f
C102 plus.t2 a_n1296_n1488# 0.080976f
C103 plus.n1 a_n1296_n1488# 0.05588f
C104 plus.n2 a_n1296_n1488# 0.045578f
C105 plus.n3 a_n1296_n1488# 0.013233f
C106 plus.n4 a_n1296_n1488# 0.045578f
C107 plus.t0 a_n1296_n1488# 0.080976f
C108 plus.n5 a_n1296_n1488# 0.055827f
C109 plus.n6 a_n1296_n1488# 0.259446f
C110 plus.n7 a_n1296_n1488# 0.079891f
C111 plus.t7 a_n1296_n1488# 0.080976f
C112 plus.t5 a_n1296_n1488# 0.075423f
C113 plus.t3 a_n1296_n1488# 0.075423f
C114 plus.t4 a_n1296_n1488# 0.080976f
C115 plus.n8 a_n1296_n1488# 0.05588f
C116 plus.n9 a_n1296_n1488# 0.045578f
C117 plus.n10 a_n1296_n1488# 0.013233f
C118 plus.n11 a_n1296_n1488# 0.045578f
C119 plus.n12 a_n1296_n1488# 0.055827f
C120 plus.n13 a_n1296_n1488# 0.720017f
.ends

