* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 a_n1352_n1088# a_n1352_n1088# a_n1352_n1088# a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.2
X1 drain_right.t9 minus.t0 source.t11 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X2 drain_right.t8 minus.t1 source.t15 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X3 drain_left.t9 plus.t0 source.t9 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X4 source.t5 plus.t1 drain_left.t8 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X5 a_n1352_n1088# a_n1352_n1088# a_n1352_n1088# a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.2
X6 source.t12 minus.t2 drain_right.t7 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X7 source.t18 minus.t3 drain_right.t6 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X8 drain_left.t7 plus.t2 source.t1 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.2
X9 drain_right.t5 minus.t4 source.t16 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.2
X10 drain_left.t6 plus.t3 source.t8 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.2
X11 drain_right.t4 minus.t5 source.t17 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.2
X12 drain_right.t3 minus.t6 source.t13 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.2
X13 drain_right.t2 minus.t7 source.t10 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.2
X14 source.t14 minus.t8 drain_right.t1 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X15 source.t2 plus.t4 drain_left.t5 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X16 drain_left.t4 plus.t5 source.t7 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.2
X17 source.t6 plus.t6 drain_left.t3 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X18 source.t3 plus.t7 drain_left.t2 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X19 source.t19 minus.t9 drain_right.t0 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
X20 a_n1352_n1088# a_n1352_n1088# a_n1352_n1088# a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.2
X21 a_n1352_n1088# a_n1352_n1088# a_n1352_n1088# a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.2
X22 drain_left.t1 plus.t8 source.t4 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.2
X23 drain_left.t0 plus.t9 source.t0 a_n1352_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.2
R0 minus.n8 minus.t6 322.43
R1 minus.n2 minus.t5 322.43
R2 minus.n18 minus.t7 322.43
R3 minus.n12 minus.t4 322.43
R4 minus.n7 minus.t9 277.151
R5 minus.n5 minus.t0 277.151
R6 minus.n1 minus.t2 277.151
R7 minus.n17 minus.t3 277.151
R8 minus.n15 minus.t1 277.151
R9 minus.n11 minus.t8 277.151
R10 minus.n3 minus.n2 161.489
R11 minus.n13 minus.n12 161.489
R12 minus.n9 minus.n8 161.3
R13 minus.n6 minus.n0 161.3
R14 minus.n4 minus.n3 161.3
R15 minus.n19 minus.n18 161.3
R16 minus.n16 minus.n10 161.3
R17 minus.n14 minus.n13 161.3
R18 minus.n7 minus.n6 40.8975
R19 minus.n4 minus.n1 40.8975
R20 minus.n14 minus.n11 40.8975
R21 minus.n17 minus.n16 40.8975
R22 minus.n6 minus.n5 36.5157
R23 minus.n5 minus.n4 36.5157
R24 minus.n15 minus.n14 36.5157
R25 minus.n16 minus.n15 36.5157
R26 minus.n8 minus.n7 32.1338
R27 minus.n2 minus.n1 32.1338
R28 minus.n12 minus.n11 32.1338
R29 minus.n18 minus.n17 32.1338
R30 minus.n20 minus.n9 25.8585
R31 minus.n20 minus.n19 6.44936
R32 minus.n9 minus.n0 0.189894
R33 minus.n3 minus.n0 0.189894
R34 minus.n13 minus.n10 0.189894
R35 minus.n19 minus.n10 0.189894
R36 minus minus.n20 0.188
R37 source.n0 source.t7 243.255
R38 source.n5 source.t17 243.255
R39 source.n19 source.t10 243.254
R40 source.n14 source.t8 243.254
R41 source.n2 source.n1 223.454
R42 source.n4 source.n3 223.454
R43 source.n7 source.n6 223.454
R44 source.n9 source.n8 223.454
R45 source.n18 source.n17 223.453
R46 source.n16 source.n15 223.453
R47 source.n13 source.n12 223.453
R48 source.n11 source.n10 223.453
R49 source.n17 source.t15 19.8005
R50 source.n17 source.t18 19.8005
R51 source.n15 source.t16 19.8005
R52 source.n15 source.t14 19.8005
R53 source.n12 source.t9 19.8005
R54 source.n12 source.t3 19.8005
R55 source.n10 source.t4 19.8005
R56 source.n10 source.t2 19.8005
R57 source.n1 source.t0 19.8005
R58 source.n1 source.t6 19.8005
R59 source.n3 source.t1 19.8005
R60 source.n3 source.t5 19.8005
R61 source.n6 source.t11 19.8005
R62 source.n6 source.t12 19.8005
R63 source.n8 source.t13 19.8005
R64 source.n8 source.t19 19.8005
R65 source.n11 source.n9 13.8682
R66 source.n20 source.n0 7.91991
R67 source.n20 source.n19 5.49188
R68 source.n5 source.n4 0.698776
R69 source.n16 source.n14 0.698776
R70 source.n9 source.n7 0.457397
R71 source.n7 source.n5 0.457397
R72 source.n4 source.n2 0.457397
R73 source.n2 source.n0 0.457397
R74 source.n13 source.n11 0.457397
R75 source.n14 source.n13 0.457397
R76 source.n18 source.n16 0.457397
R77 source.n19 source.n18 0.457397
R78 source source.n20 0.188
R79 drain_right.n1 drain_right.t5 260.389
R80 drain_right.n7 drain_right.t3 259.933
R81 drain_right.n6 drain_right.n4 240.589
R82 drain_right.n3 drain_right.n2 240.419
R83 drain_right.n6 drain_right.n5 240.132
R84 drain_right.n1 drain_right.n0 240.131
R85 drain_right drain_right.n3 20.4223
R86 drain_right.n2 drain_right.t6 19.8005
R87 drain_right.n2 drain_right.t2 19.8005
R88 drain_right.n0 drain_right.t1 19.8005
R89 drain_right.n0 drain_right.t8 19.8005
R90 drain_right.n4 drain_right.t7 19.8005
R91 drain_right.n4 drain_right.t4 19.8005
R92 drain_right.n5 drain_right.t0 19.8005
R93 drain_right.n5 drain_right.t9 19.8005
R94 drain_right drain_right.n7 5.88166
R95 drain_right.n7 drain_right.n6 0.457397
R96 drain_right.n3 drain_right.n1 0.0593781
R97 plus.n2 plus.t2 322.43
R98 plus.n8 plus.t5 322.43
R99 plus.n12 plus.t3 322.43
R100 plus.n18 plus.t8 322.43
R101 plus.n1 plus.t1 277.151
R102 plus.n5 plus.t9 277.151
R103 plus.n7 plus.t6 277.151
R104 plus.n11 plus.t7 277.151
R105 plus.n15 plus.t0 277.151
R106 plus.n17 plus.t4 277.151
R107 plus.n3 plus.n2 161.489
R108 plus.n13 plus.n12 161.489
R109 plus.n4 plus.n3 161.3
R110 plus.n6 plus.n0 161.3
R111 plus.n9 plus.n8 161.3
R112 plus.n14 plus.n13 161.3
R113 plus.n16 plus.n10 161.3
R114 plus.n19 plus.n18 161.3
R115 plus.n4 plus.n1 40.8975
R116 plus.n7 plus.n6 40.8975
R117 plus.n17 plus.n16 40.8975
R118 plus.n14 plus.n11 40.8975
R119 plus.n5 plus.n4 36.5157
R120 plus.n6 plus.n5 36.5157
R121 plus.n16 plus.n15 36.5157
R122 plus.n15 plus.n14 36.5157
R123 plus.n2 plus.n1 32.1338
R124 plus.n8 plus.n7 32.1338
R125 plus.n18 plus.n17 32.1338
R126 plus.n12 plus.n11 32.1338
R127 plus plus.n19 23.9062
R128 plus plus.n9 7.92664
R129 plus.n3 plus.n0 0.189894
R130 plus.n9 plus.n0 0.189894
R131 plus.n19 plus.n10 0.189894
R132 plus.n13 plus.n10 0.189894
R133 drain_left.n5 drain_left.t7 260.389
R134 drain_left.n1 drain_left.t1 260.389
R135 drain_left.n3 drain_left.n2 240.419
R136 drain_left.n7 drain_left.n6 240.132
R137 drain_left.n5 drain_left.n4 240.132
R138 drain_left.n1 drain_left.n0 240.131
R139 drain_left drain_left.n3 20.9755
R140 drain_left.n2 drain_left.t2 19.8005
R141 drain_left.n2 drain_left.t6 19.8005
R142 drain_left.n0 drain_left.t5 19.8005
R143 drain_left.n0 drain_left.t9 19.8005
R144 drain_left.n6 drain_left.t3 19.8005
R145 drain_left.n6 drain_left.t4 19.8005
R146 drain_left.n4 drain_left.t8 19.8005
R147 drain_left.n4 drain_left.t0 19.8005
R148 drain_left drain_left.n7 6.11011
R149 drain_left.n7 drain_left.n5 0.457397
R150 drain_left.n3 drain_left.n1 0.0593781
C0 drain_left minus 0.178307f
C1 drain_right minus 0.606675f
C2 drain_left source 3.97779f
C3 drain_right source 3.97491f
C4 drain_left plus 0.734329f
C5 drain_right plus 0.29013f
C6 drain_left drain_right 0.658344f
C7 minus source 0.749509f
C8 plus minus 2.8128f
C9 plus source 0.763431f
C10 drain_right a_n1352_n1088# 3.14687f
C11 drain_left a_n1352_n1088# 3.32399f
C12 source a_n1352_n1088# 1.980342f
C13 minus a_n1352_n1088# 4.318577f
C14 plus a_n1352_n1088# 5.044781f
C15 drain_left.t1 a_n1352_n1088# 0.121868f
C16 drain_left.t5 a_n1352_n1088# 0.019638f
C17 drain_left.t9 a_n1352_n1088# 0.019638f
C18 drain_left.n0 a_n1352_n1088# 0.076306f
C19 drain_left.n1 a_n1352_n1088# 0.45324f
C20 drain_left.t2 a_n1352_n1088# 0.019638f
C21 drain_left.t6 a_n1352_n1088# 0.019638f
C22 drain_left.n2 a_n1352_n1088# 0.076599f
C23 drain_left.n3 a_n1352_n1088# 0.783469f
C24 drain_left.t7 a_n1352_n1088# 0.121869f
C25 drain_left.t8 a_n1352_n1088# 0.019638f
C26 drain_left.t0 a_n1352_n1088# 0.019638f
C27 drain_left.n4 a_n1352_n1088# 0.076306f
C28 drain_left.n5 a_n1352_n1088# 0.475326f
C29 drain_left.t3 a_n1352_n1088# 0.019638f
C30 drain_left.t4 a_n1352_n1088# 0.019638f
C31 drain_left.n6 a_n1352_n1088# 0.076306f
C32 drain_left.n7 a_n1352_n1088# 0.450332f
C33 plus.n0 a_n1352_n1088# 0.038675f
C34 plus.t6 a_n1352_n1088# 0.023845f
C35 plus.t9 a_n1352_n1088# 0.023845f
C36 plus.t1 a_n1352_n1088# 0.023845f
C37 plus.n1 a_n1352_n1088# 0.028541f
C38 plus.t2 a_n1352_n1088# 0.027886f
C39 plus.n2 a_n1352_n1088# 0.038337f
C40 plus.n3 a_n1352_n1088# 0.084925f
C41 plus.n4 a_n1352_n1088# 0.013545f
C42 plus.n5 a_n1352_n1088# 0.028541f
C43 plus.n6 a_n1352_n1088# 0.013545f
C44 plus.n7 a_n1352_n1088# 0.028541f
C45 plus.t5 a_n1352_n1088# 0.027886f
C46 plus.n8 a_n1352_n1088# 0.038283f
C47 plus.n9 a_n1352_n1088# 0.26028f
C48 plus.n10 a_n1352_n1088# 0.038675f
C49 plus.t8 a_n1352_n1088# 0.027886f
C50 plus.t4 a_n1352_n1088# 0.023845f
C51 plus.t0 a_n1352_n1088# 0.023845f
C52 plus.t7 a_n1352_n1088# 0.023845f
C53 plus.n11 a_n1352_n1088# 0.028541f
C54 plus.t3 a_n1352_n1088# 0.027886f
C55 plus.n12 a_n1352_n1088# 0.038337f
C56 plus.n13 a_n1352_n1088# 0.084925f
C57 plus.n14 a_n1352_n1088# 0.013545f
C58 plus.n15 a_n1352_n1088# 0.028541f
C59 plus.n16 a_n1352_n1088# 0.013545f
C60 plus.n17 a_n1352_n1088# 0.028541f
C61 plus.n18 a_n1352_n1088# 0.038283f
C62 plus.n19 a_n1352_n1088# 0.7527f
C63 drain_right.t5 a_n1352_n1088# 0.124904f
C64 drain_right.t1 a_n1352_n1088# 0.020127f
C65 drain_right.t8 a_n1352_n1088# 0.020127f
C66 drain_right.n0 a_n1352_n1088# 0.078207f
C67 drain_right.n1 a_n1352_n1088# 0.464529f
C68 drain_right.t6 a_n1352_n1088# 0.020127f
C69 drain_right.t2 a_n1352_n1088# 0.020127f
C70 drain_right.n2 a_n1352_n1088# 0.078507f
C71 drain_right.n3 a_n1352_n1088# 0.7536f
C72 drain_right.t7 a_n1352_n1088# 0.020127f
C73 drain_right.t4 a_n1352_n1088# 0.020127f
C74 drain_right.n4 a_n1352_n1088# 0.078707f
C75 drain_right.t0 a_n1352_n1088# 0.020127f
C76 drain_right.t9 a_n1352_n1088# 0.020127f
C77 drain_right.n5 a_n1352_n1088# 0.078207f
C78 drain_right.n6 a_n1352_n1088# 0.515968f
C79 drain_right.t3 a_n1352_n1088# 0.124493f
C80 drain_right.n7 a_n1352_n1088# 0.441482f
C81 source.t7 a_n1352_n1088# 0.148309f
C82 source.n0 a_n1352_n1088# 0.620016f
C83 source.t0 a_n1352_n1088# 0.026646f
C84 source.t6 a_n1352_n1088# 0.026646f
C85 source.n1 a_n1352_n1088# 0.086418f
C86 source.n2 a_n1352_n1088# 0.30638f
C87 source.t1 a_n1352_n1088# 0.026646f
C88 source.t5 a_n1352_n1088# 0.026646f
C89 source.n3 a_n1352_n1088# 0.086418f
C90 source.n4 a_n1352_n1088# 0.332606f
C91 source.t17 a_n1352_n1088# 0.148309f
C92 source.n5 a_n1352_n1088# 0.343386f
C93 source.t11 a_n1352_n1088# 0.026646f
C94 source.t12 a_n1352_n1088# 0.026646f
C95 source.n6 a_n1352_n1088# 0.086418f
C96 source.n7 a_n1352_n1088# 0.30638f
C97 source.t13 a_n1352_n1088# 0.026646f
C98 source.t19 a_n1352_n1088# 0.026646f
C99 source.n8 a_n1352_n1088# 0.086418f
C100 source.n9 a_n1352_n1088# 0.927139f
C101 source.t4 a_n1352_n1088# 0.026646f
C102 source.t2 a_n1352_n1088# 0.026646f
C103 source.n10 a_n1352_n1088# 0.086418f
C104 source.n11 a_n1352_n1088# 0.927139f
C105 source.t9 a_n1352_n1088# 0.026646f
C106 source.t3 a_n1352_n1088# 0.026646f
C107 source.n12 a_n1352_n1088# 0.086418f
C108 source.n13 a_n1352_n1088# 0.30638f
C109 source.t8 a_n1352_n1088# 0.148309f
C110 source.n14 a_n1352_n1088# 0.343386f
C111 source.t16 a_n1352_n1088# 0.026646f
C112 source.t14 a_n1352_n1088# 0.026646f
C113 source.n15 a_n1352_n1088# 0.086418f
C114 source.n16 a_n1352_n1088# 0.332606f
C115 source.t15 a_n1352_n1088# 0.026646f
C116 source.t18 a_n1352_n1088# 0.026646f
C117 source.n17 a_n1352_n1088# 0.086418f
C118 source.n18 a_n1352_n1088# 0.30638f
C119 source.t10 a_n1352_n1088# 0.148309f
C120 source.n19 a_n1352_n1088# 0.501403f
C121 source.n20 a_n1352_n1088# 0.67912f
C122 minus.n0 a_n1352_n1088# 0.037624f
C123 minus.t6 a_n1352_n1088# 0.027128f
C124 minus.t9 a_n1352_n1088# 0.023197f
C125 minus.t0 a_n1352_n1088# 0.023197f
C126 minus.t2 a_n1352_n1088# 0.023197f
C127 minus.n1 a_n1352_n1088# 0.027766f
C128 minus.t5 a_n1352_n1088# 0.027128f
C129 minus.n2 a_n1352_n1088# 0.037296f
C130 minus.n3 a_n1352_n1088# 0.082617f
C131 minus.n4 a_n1352_n1088# 0.013177f
C132 minus.n5 a_n1352_n1088# 0.027766f
C133 minus.n6 a_n1352_n1088# 0.013177f
C134 minus.n7 a_n1352_n1088# 0.027766f
C135 minus.n8 a_n1352_n1088# 0.037243f
C136 minus.n9 a_n1352_n1088# 0.749641f
C137 minus.n10 a_n1352_n1088# 0.037624f
C138 minus.t3 a_n1352_n1088# 0.023197f
C139 minus.t1 a_n1352_n1088# 0.023197f
C140 minus.t8 a_n1352_n1088# 0.023197f
C141 minus.n11 a_n1352_n1088# 0.027766f
C142 minus.t4 a_n1352_n1088# 0.027128f
C143 minus.n12 a_n1352_n1088# 0.037296f
C144 minus.n13 a_n1352_n1088# 0.082617f
C145 minus.n14 a_n1352_n1088# 0.013177f
C146 minus.n15 a_n1352_n1088# 0.027766f
C147 minus.n16 a_n1352_n1088# 0.013177f
C148 minus.n17 a_n1352_n1088# 0.027766f
C149 minus.t7 a_n1352_n1088# 0.027128f
C150 minus.n18 a_n1352_n1088# 0.037243f
C151 minus.n19 a_n1352_n1088# 0.241475f
C152 minus.n20 a_n1352_n1088# 0.927624f
.ends

