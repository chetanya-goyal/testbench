* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t29 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X1 source.t30 plus.t1 drain_left.t18 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X2 source.t25 plus.t2 drain_left.t17 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X3 source.t24 plus.t3 drain_left.t16 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X4 source.t2 minus.t0 drain_right.t19 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X5 source.t0 minus.t1 drain_right.t18 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X6 drain_right.t17 minus.t2 source.t1 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X7 drain_left.t15 plus.t4 source.t26 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X8 a_n2982_n1288# a_n2982_n1288# a_n2982_n1288# a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.7
X9 drain_left.t14 plus.t5 source.t20 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X10 source.t31 plus.t6 drain_left.t13 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X11 source.t34 plus.t7 drain_left.t12 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X12 drain_right.t16 minus.t3 source.t4 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X13 a_n2982_n1288# a_n2982_n1288# a_n2982_n1288# a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X14 source.t9 minus.t4 drain_right.t15 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X15 drain_right.t14 minus.t5 source.t5 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X16 drain_left.t11 plus.t8 source.t22 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X17 source.t23 plus.t9 drain_left.t10 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X18 drain_right.t13 minus.t6 source.t16 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X19 drain_right.t12 minus.t7 source.t18 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X20 drain_left.t9 plus.t10 source.t39 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X21 drain_right.t11 minus.t8 source.t6 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X22 drain_left.t8 plus.t11 source.t33 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X23 drain_left.t7 plus.t12 source.t36 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X24 source.t28 plus.t13 drain_left.t6 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X25 drain_left.t5 plus.t14 source.t35 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X26 drain_right.t10 minus.t9 source.t12 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X27 drain_right.t9 minus.t10 source.t15 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X28 source.t3 minus.t11 drain_right.t8 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X29 drain_left.t4 plus.t15 source.t37 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X30 a_n2982_n1288# a_n2982_n1288# a_n2982_n1288# a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X31 source.t14 minus.t12 drain_right.t7 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X32 a_n2982_n1288# a_n2982_n1288# a_n2982_n1288# a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X33 source.t27 plus.t16 drain_left.t3 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X34 drain_right.t6 minus.t13 source.t7 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X35 source.t19 minus.t14 drain_right.t5 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X36 source.t10 minus.t15 drain_right.t4 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X37 drain_right.t3 minus.t16 source.t13 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X38 source.t17 minus.t17 drain_right.t2 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X39 source.t38 plus.t17 drain_left.t2 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X40 drain_left.t1 plus.t18 source.t32 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X41 source.t8 minus.t18 drain_right.t1 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X42 source.t11 minus.t19 drain_right.t0 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X43 source.t21 plus.t19 drain_left.t0 a_n2982_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
R0 plus.n11 plus.n10 161.3
R1 plus.n12 plus.n7 161.3
R2 plus.n14 plus.n13 161.3
R3 plus.n15 plus.n6 161.3
R4 plus.n17 plus.n16 161.3
R5 plus.n18 plus.n5 161.3
R6 plus.n20 plus.n19 161.3
R7 plus.n21 plus.n4 161.3
R8 plus.n23 plus.n22 161.3
R9 plus.n24 plus.n3 161.3
R10 plus.n26 plus.n25 161.3
R11 plus.n27 plus.n2 161.3
R12 plus.n29 plus.n28 161.3
R13 plus.n30 plus.n1 161.3
R14 plus.n31 plus.n0 161.3
R15 plus.n33 plus.n32 161.3
R16 plus.n45 plus.n44 161.3
R17 plus.n46 plus.n41 161.3
R18 plus.n48 plus.n47 161.3
R19 plus.n49 plus.n40 161.3
R20 plus.n51 plus.n50 161.3
R21 plus.n52 plus.n39 161.3
R22 plus.n54 plus.n53 161.3
R23 plus.n55 plus.n38 161.3
R24 plus.n57 plus.n56 161.3
R25 plus.n58 plus.n37 161.3
R26 plus.n60 plus.n59 161.3
R27 plus.n61 plus.n36 161.3
R28 plus.n63 plus.n62 161.3
R29 plus.n64 plus.n35 161.3
R30 plus.n65 plus.n34 161.3
R31 plus.n67 plus.n66 161.3
R32 plus.n9 plus.t7 150.369
R33 plus.n43 plus.t18 150.369
R34 plus.n32 plus.t5 124.977
R35 plus.n30 plus.t19 124.977
R36 plus.n2 plus.t10 124.977
R37 plus.n24 plus.t2 124.977
R38 plus.n4 plus.t14 124.977
R39 plus.n18 plus.t6 124.977
R40 plus.n6 plus.t12 124.977
R41 plus.n12 plus.t3 124.977
R42 plus.n8 plus.t15 124.977
R43 plus.n66 plus.t1 124.977
R44 plus.n64 plus.t0 124.977
R45 plus.n36 plus.t16 124.977
R46 plus.n58 plus.t11 124.977
R47 plus.n38 plus.t13 124.977
R48 plus.n52 plus.t8 124.977
R49 plus.n40 plus.t9 124.977
R50 plus.n46 plus.t4 124.977
R51 plus.n42 plus.t17 124.977
R52 plus.n10 plus.n9 45.0031
R53 plus.n44 plus.n43 45.0031
R54 plus.n32 plus.n31 41.6278
R55 plus.n66 plus.n65 41.6278
R56 plus.n30 plus.n29 37.246
R57 plus.n11 plus.n8 37.246
R58 plus.n64 plus.n63 37.246
R59 plus.n45 plus.n42 37.246
R60 plus.n25 plus.n2 32.8641
R61 plus.n13 plus.n12 32.8641
R62 plus.n59 plus.n36 32.8641
R63 plus.n47 plus.n46 32.8641
R64 plus plus.n67 30.6771
R65 plus.n24 plus.n23 28.4823
R66 plus.n17 plus.n6 28.4823
R67 plus.n58 plus.n57 28.4823
R68 plus.n51 plus.n40 28.4823
R69 plus.n19 plus.n18 24.1005
R70 plus.n19 plus.n4 24.1005
R71 plus.n53 plus.n38 24.1005
R72 plus.n53 plus.n52 24.1005
R73 plus.n23 plus.n4 19.7187
R74 plus.n18 plus.n17 19.7187
R75 plus.n57 plus.n38 19.7187
R76 plus.n52 plus.n51 19.7187
R77 plus.n9 plus.n8 15.6319
R78 plus.n43 plus.n42 15.6319
R79 plus.n25 plus.n24 15.3369
R80 plus.n13 plus.n6 15.3369
R81 plus.n59 plus.n58 15.3369
R82 plus.n47 plus.n40 15.3369
R83 plus.n29 plus.n2 10.955
R84 plus.n12 plus.n11 10.955
R85 plus.n63 plus.n36 10.955
R86 plus.n46 plus.n45 10.955
R87 plus plus.n33 8.52323
R88 plus.n31 plus.n30 6.57323
R89 plus.n65 plus.n64 6.57323
R90 plus.n10 plus.n7 0.189894
R91 plus.n14 plus.n7 0.189894
R92 plus.n15 plus.n14 0.189894
R93 plus.n16 plus.n15 0.189894
R94 plus.n16 plus.n5 0.189894
R95 plus.n20 plus.n5 0.189894
R96 plus.n21 plus.n20 0.189894
R97 plus.n22 plus.n21 0.189894
R98 plus.n22 plus.n3 0.189894
R99 plus.n26 plus.n3 0.189894
R100 plus.n27 plus.n26 0.189894
R101 plus.n28 plus.n27 0.189894
R102 plus.n28 plus.n1 0.189894
R103 plus.n1 plus.n0 0.189894
R104 plus.n33 plus.n0 0.189894
R105 plus.n67 plus.n34 0.189894
R106 plus.n35 plus.n34 0.189894
R107 plus.n62 plus.n35 0.189894
R108 plus.n62 plus.n61 0.189894
R109 plus.n61 plus.n60 0.189894
R110 plus.n60 plus.n37 0.189894
R111 plus.n56 plus.n37 0.189894
R112 plus.n56 plus.n55 0.189894
R113 plus.n55 plus.n54 0.189894
R114 plus.n54 plus.n39 0.189894
R115 plus.n50 plus.n39 0.189894
R116 plus.n50 plus.n49 0.189894
R117 plus.n49 plus.n48 0.189894
R118 plus.n48 plus.n41 0.189894
R119 plus.n44 plus.n41 0.189894
R120 source.n90 source.n88 289.615
R121 source.n74 source.n72 289.615
R122 source.n66 source.n64 289.615
R123 source.n50 source.n48 289.615
R124 source.n2 source.n0 289.615
R125 source.n18 source.n16 289.615
R126 source.n26 source.n24 289.615
R127 source.n42 source.n40 289.615
R128 source.n91 source.n90 185
R129 source.n75 source.n74 185
R130 source.n67 source.n66 185
R131 source.n51 source.n50 185
R132 source.n3 source.n2 185
R133 source.n19 source.n18 185
R134 source.n27 source.n26 185
R135 source.n43 source.n42 185
R136 source.t13 source.n89 167.117
R137 source.t3 source.n73 167.117
R138 source.t32 source.n65 167.117
R139 source.t30 source.n49 167.117
R140 source.t20 source.n1 167.117
R141 source.t34 source.n17 167.117
R142 source.t15 source.n25 167.117
R143 source.t14 source.n41 167.117
R144 source.n9 source.n8 84.1169
R145 source.n11 source.n10 84.1169
R146 source.n13 source.n12 84.1169
R147 source.n15 source.n14 84.1169
R148 source.n33 source.n32 84.1169
R149 source.n35 source.n34 84.1169
R150 source.n37 source.n36 84.1169
R151 source.n39 source.n38 84.1169
R152 source.n87 source.n86 84.1168
R153 source.n85 source.n84 84.1168
R154 source.n83 source.n82 84.1168
R155 source.n81 source.n80 84.1168
R156 source.n63 source.n62 84.1168
R157 source.n61 source.n60 84.1168
R158 source.n59 source.n58 84.1168
R159 source.n57 source.n56 84.1168
R160 source.n90 source.t13 52.3082
R161 source.n74 source.t3 52.3082
R162 source.n66 source.t32 52.3082
R163 source.n50 source.t30 52.3082
R164 source.n2 source.t20 52.3082
R165 source.n18 source.t34 52.3082
R166 source.n26 source.t15 52.3082
R167 source.n42 source.t14 52.3082
R168 source.n95 source.n94 31.4096
R169 source.n79 source.n78 31.4096
R170 source.n71 source.n70 31.4096
R171 source.n55 source.n54 31.4096
R172 source.n7 source.n6 31.4096
R173 source.n23 source.n22 31.4096
R174 source.n31 source.n30 31.4096
R175 source.n47 source.n46 31.4096
R176 source.n55 source.n47 14.5999
R177 source.n86 source.t5 9.9005
R178 source.n86 source.t9 9.9005
R179 source.n84 source.t1 9.9005
R180 source.n84 source.t0 9.9005
R181 source.n82 source.t7 9.9005
R182 source.n82 source.t17 9.9005
R183 source.n80 source.t12 9.9005
R184 source.n80 source.t10 9.9005
R185 source.n62 source.t26 9.9005
R186 source.n62 source.t38 9.9005
R187 source.n60 source.t22 9.9005
R188 source.n60 source.t23 9.9005
R189 source.n58 source.t33 9.9005
R190 source.n58 source.t28 9.9005
R191 source.n56 source.t29 9.9005
R192 source.n56 source.t27 9.9005
R193 source.n8 source.t39 9.9005
R194 source.n8 source.t21 9.9005
R195 source.n10 source.t35 9.9005
R196 source.n10 source.t25 9.9005
R197 source.n12 source.t36 9.9005
R198 source.n12 source.t31 9.9005
R199 source.n14 source.t37 9.9005
R200 source.n14 source.t24 9.9005
R201 source.n32 source.t6 9.9005
R202 source.n32 source.t2 9.9005
R203 source.n34 source.t18 9.9005
R204 source.n34 source.t8 9.9005
R205 source.n36 source.t16 9.9005
R206 source.n36 source.t11 9.9005
R207 source.n38 source.t4 9.9005
R208 source.n38 source.t19 9.9005
R209 source.n91 source.n89 9.71174
R210 source.n75 source.n73 9.71174
R211 source.n67 source.n65 9.71174
R212 source.n51 source.n49 9.71174
R213 source.n3 source.n1 9.71174
R214 source.n19 source.n17 9.71174
R215 source.n27 source.n25 9.71174
R216 source.n43 source.n41 9.71174
R217 source.n94 source.n93 9.45567
R218 source.n78 source.n77 9.45567
R219 source.n70 source.n69 9.45567
R220 source.n54 source.n53 9.45567
R221 source.n6 source.n5 9.45567
R222 source.n22 source.n21 9.45567
R223 source.n30 source.n29 9.45567
R224 source.n46 source.n45 9.45567
R225 source.n93 source.n92 9.3005
R226 source.n77 source.n76 9.3005
R227 source.n69 source.n68 9.3005
R228 source.n53 source.n52 9.3005
R229 source.n5 source.n4 9.3005
R230 source.n21 source.n20 9.3005
R231 source.n29 source.n28 9.3005
R232 source.n45 source.n44 9.3005
R233 source.n96 source.n7 8.893
R234 source.n94 source.n88 8.14595
R235 source.n78 source.n72 8.14595
R236 source.n70 source.n64 8.14595
R237 source.n54 source.n48 8.14595
R238 source.n6 source.n0 8.14595
R239 source.n22 source.n16 8.14595
R240 source.n30 source.n24 8.14595
R241 source.n46 source.n40 8.14595
R242 source.n92 source.n91 7.3702
R243 source.n76 source.n75 7.3702
R244 source.n68 source.n67 7.3702
R245 source.n52 source.n51 7.3702
R246 source.n4 source.n3 7.3702
R247 source.n20 source.n19 7.3702
R248 source.n28 source.n27 7.3702
R249 source.n44 source.n43 7.3702
R250 source.n92 source.n88 5.81868
R251 source.n76 source.n72 5.81868
R252 source.n68 source.n64 5.81868
R253 source.n52 source.n48 5.81868
R254 source.n4 source.n0 5.81868
R255 source.n20 source.n16 5.81868
R256 source.n28 source.n24 5.81868
R257 source.n44 source.n40 5.81868
R258 source.n96 source.n95 5.7074
R259 source.n93 source.n89 3.44771
R260 source.n77 source.n73 3.44771
R261 source.n69 source.n65 3.44771
R262 source.n53 source.n49 3.44771
R263 source.n5 source.n1 3.44771
R264 source.n21 source.n17 3.44771
R265 source.n29 source.n25 3.44771
R266 source.n45 source.n41 3.44771
R267 source.n47 source.n39 0.888431
R268 source.n39 source.n37 0.888431
R269 source.n37 source.n35 0.888431
R270 source.n35 source.n33 0.888431
R271 source.n33 source.n31 0.888431
R272 source.n23 source.n15 0.888431
R273 source.n15 source.n13 0.888431
R274 source.n13 source.n11 0.888431
R275 source.n11 source.n9 0.888431
R276 source.n9 source.n7 0.888431
R277 source.n57 source.n55 0.888431
R278 source.n59 source.n57 0.888431
R279 source.n61 source.n59 0.888431
R280 source.n63 source.n61 0.888431
R281 source.n71 source.n63 0.888431
R282 source.n81 source.n79 0.888431
R283 source.n83 source.n81 0.888431
R284 source.n85 source.n83 0.888431
R285 source.n87 source.n85 0.888431
R286 source.n95 source.n87 0.888431
R287 source.n31 source.n23 0.470328
R288 source.n79 source.n71 0.470328
R289 source source.n96 0.188
R290 drain_left.n10 drain_left.n8 101.683
R291 drain_left.n6 drain_left.n4 101.683
R292 drain_left.n2 drain_left.n0 101.683
R293 drain_left.n16 drain_left.n15 100.796
R294 drain_left.n14 drain_left.n13 100.796
R295 drain_left.n12 drain_left.n11 100.796
R296 drain_left.n10 drain_left.n9 100.796
R297 drain_left.n7 drain_left.n3 100.796
R298 drain_left.n6 drain_left.n5 100.796
R299 drain_left.n2 drain_left.n1 100.796
R300 drain_left drain_left.n7 26.8948
R301 drain_left.n3 drain_left.t6 9.9005
R302 drain_left.n3 drain_left.t11 9.9005
R303 drain_left.n4 drain_left.t2 9.9005
R304 drain_left.n4 drain_left.t1 9.9005
R305 drain_left.n5 drain_left.t10 9.9005
R306 drain_left.n5 drain_left.t15 9.9005
R307 drain_left.n1 drain_left.t3 9.9005
R308 drain_left.n1 drain_left.t8 9.9005
R309 drain_left.n0 drain_left.t18 9.9005
R310 drain_left.n0 drain_left.t19 9.9005
R311 drain_left.n15 drain_left.t0 9.9005
R312 drain_left.n15 drain_left.t14 9.9005
R313 drain_left.n13 drain_left.t17 9.9005
R314 drain_left.n13 drain_left.t9 9.9005
R315 drain_left.n11 drain_left.t13 9.9005
R316 drain_left.n11 drain_left.t5 9.9005
R317 drain_left.n9 drain_left.t16 9.9005
R318 drain_left.n9 drain_left.t7 9.9005
R319 drain_left.n8 drain_left.t12 9.9005
R320 drain_left.n8 drain_left.t4 9.9005
R321 drain_left drain_left.n16 6.54115
R322 drain_left.n12 drain_left.n10 0.888431
R323 drain_left.n14 drain_left.n12 0.888431
R324 drain_left.n16 drain_left.n14 0.888431
R325 drain_left.n7 drain_left.n6 0.833085
R326 drain_left.n7 drain_left.n2 0.833085
R327 minus.n33 minus.n32 161.3
R328 minus.n31 minus.n0 161.3
R329 minus.n30 minus.n29 161.3
R330 minus.n28 minus.n1 161.3
R331 minus.n27 minus.n26 161.3
R332 minus.n25 minus.n2 161.3
R333 minus.n24 minus.n23 161.3
R334 minus.n22 minus.n3 161.3
R335 minus.n21 minus.n20 161.3
R336 minus.n19 minus.n4 161.3
R337 minus.n18 minus.n17 161.3
R338 minus.n16 minus.n5 161.3
R339 minus.n15 minus.n14 161.3
R340 minus.n13 minus.n6 161.3
R341 minus.n12 minus.n11 161.3
R342 minus.n10 minus.n7 161.3
R343 minus.n67 minus.n66 161.3
R344 minus.n65 minus.n34 161.3
R345 minus.n64 minus.n63 161.3
R346 minus.n62 minus.n35 161.3
R347 minus.n61 minus.n60 161.3
R348 minus.n59 minus.n36 161.3
R349 minus.n58 minus.n57 161.3
R350 minus.n56 minus.n37 161.3
R351 minus.n55 minus.n54 161.3
R352 minus.n53 minus.n38 161.3
R353 minus.n52 minus.n51 161.3
R354 minus.n50 minus.n39 161.3
R355 minus.n49 minus.n48 161.3
R356 minus.n47 minus.n40 161.3
R357 minus.n46 minus.n45 161.3
R358 minus.n44 minus.n41 161.3
R359 minus.n9 minus.t10 150.369
R360 minus.n43 minus.t11 150.369
R361 minus.n8 minus.t0 124.977
R362 minus.n12 minus.t8 124.977
R363 minus.n14 minus.t18 124.977
R364 minus.n18 minus.t7 124.977
R365 minus.n20 minus.t19 124.977
R366 minus.n24 minus.t6 124.977
R367 minus.n26 minus.t14 124.977
R368 minus.n30 minus.t3 124.977
R369 minus.n32 minus.t12 124.977
R370 minus.n42 minus.t9 124.977
R371 minus.n46 minus.t15 124.977
R372 minus.n48 minus.t13 124.977
R373 minus.n52 minus.t17 124.977
R374 minus.n54 minus.t2 124.977
R375 minus.n58 minus.t1 124.977
R376 minus.n60 minus.t5 124.977
R377 minus.n64 minus.t4 124.977
R378 minus.n66 minus.t16 124.977
R379 minus.n10 minus.n9 45.0031
R380 minus.n44 minus.n43 45.0031
R381 minus.n32 minus.n31 41.6278
R382 minus.n66 minus.n65 41.6278
R383 minus.n8 minus.n7 37.246
R384 minus.n30 minus.n1 37.246
R385 minus.n42 minus.n41 37.246
R386 minus.n64 minus.n35 37.246
R387 minus.n68 minus.n33 33.0081
R388 minus.n13 minus.n12 32.8641
R389 minus.n26 minus.n25 32.8641
R390 minus.n47 minus.n46 32.8641
R391 minus.n60 minus.n59 32.8641
R392 minus.n14 minus.n5 28.4823
R393 minus.n24 minus.n3 28.4823
R394 minus.n48 minus.n39 28.4823
R395 minus.n58 minus.n37 28.4823
R396 minus.n20 minus.n19 24.1005
R397 minus.n19 minus.n18 24.1005
R398 minus.n53 minus.n52 24.1005
R399 minus.n54 minus.n53 24.1005
R400 minus.n18 minus.n5 19.7187
R401 minus.n20 minus.n3 19.7187
R402 minus.n52 minus.n39 19.7187
R403 minus.n54 minus.n37 19.7187
R404 minus.n9 minus.n8 15.6319
R405 minus.n43 minus.n42 15.6319
R406 minus.n14 minus.n13 15.3369
R407 minus.n25 minus.n24 15.3369
R408 minus.n48 minus.n47 15.3369
R409 minus.n59 minus.n58 15.3369
R410 minus.n12 minus.n7 10.955
R411 minus.n26 minus.n1 10.955
R412 minus.n46 minus.n41 10.955
R413 minus.n60 minus.n35 10.955
R414 minus.n68 minus.n67 6.66717
R415 minus.n31 minus.n30 6.57323
R416 minus.n65 minus.n64 6.57323
R417 minus.n33 minus.n0 0.189894
R418 minus.n29 minus.n0 0.189894
R419 minus.n29 minus.n28 0.189894
R420 minus.n28 minus.n27 0.189894
R421 minus.n27 minus.n2 0.189894
R422 minus.n23 minus.n2 0.189894
R423 minus.n23 minus.n22 0.189894
R424 minus.n22 minus.n21 0.189894
R425 minus.n21 minus.n4 0.189894
R426 minus.n17 minus.n4 0.189894
R427 minus.n17 minus.n16 0.189894
R428 minus.n16 minus.n15 0.189894
R429 minus.n15 minus.n6 0.189894
R430 minus.n11 minus.n6 0.189894
R431 minus.n11 minus.n10 0.189894
R432 minus.n45 minus.n44 0.189894
R433 minus.n45 minus.n40 0.189894
R434 minus.n49 minus.n40 0.189894
R435 minus.n50 minus.n49 0.189894
R436 minus.n51 minus.n50 0.189894
R437 minus.n51 minus.n38 0.189894
R438 minus.n55 minus.n38 0.189894
R439 minus.n56 minus.n55 0.189894
R440 minus.n57 minus.n56 0.189894
R441 minus.n57 minus.n36 0.189894
R442 minus.n61 minus.n36 0.189894
R443 minus.n62 minus.n61 0.189894
R444 minus.n63 minus.n62 0.189894
R445 minus.n63 minus.n34 0.189894
R446 minus.n67 minus.n34 0.189894
R447 minus minus.n68 0.188
R448 drain_right.n10 drain_right.n8 101.683
R449 drain_right.n6 drain_right.n4 101.683
R450 drain_right.n2 drain_right.n0 101.683
R451 drain_right.n10 drain_right.n9 100.796
R452 drain_right.n12 drain_right.n11 100.796
R453 drain_right.n14 drain_right.n13 100.796
R454 drain_right.n16 drain_right.n15 100.796
R455 drain_right.n7 drain_right.n3 100.796
R456 drain_right.n6 drain_right.n5 100.796
R457 drain_right.n2 drain_right.n1 100.796
R458 drain_right drain_right.n7 26.3415
R459 drain_right.n3 drain_right.t2 9.9005
R460 drain_right.n3 drain_right.t17 9.9005
R461 drain_right.n4 drain_right.t15 9.9005
R462 drain_right.n4 drain_right.t3 9.9005
R463 drain_right.n5 drain_right.t18 9.9005
R464 drain_right.n5 drain_right.t14 9.9005
R465 drain_right.n1 drain_right.t4 9.9005
R466 drain_right.n1 drain_right.t6 9.9005
R467 drain_right.n0 drain_right.t8 9.9005
R468 drain_right.n0 drain_right.t10 9.9005
R469 drain_right.n8 drain_right.t19 9.9005
R470 drain_right.n8 drain_right.t9 9.9005
R471 drain_right.n9 drain_right.t1 9.9005
R472 drain_right.n9 drain_right.t11 9.9005
R473 drain_right.n11 drain_right.t0 9.9005
R474 drain_right.n11 drain_right.t12 9.9005
R475 drain_right.n13 drain_right.t5 9.9005
R476 drain_right.n13 drain_right.t13 9.9005
R477 drain_right.n15 drain_right.t7 9.9005
R478 drain_right.n15 drain_right.t16 9.9005
R479 drain_right drain_right.n16 6.54115
R480 drain_right.n16 drain_right.n14 0.888431
R481 drain_right.n14 drain_right.n12 0.888431
R482 drain_right.n12 drain_right.n10 0.888431
R483 drain_right.n7 drain_right.n6 0.833085
R484 drain_right.n7 drain_right.n2 0.833085
C0 drain_left drain_right 1.5991f
C1 minus drain_left 0.179545f
C2 source drain_left 7.43075f
C3 minus drain_right 2.67697f
C4 source drain_right 7.43312f
C5 minus source 3.40933f
C6 plus drain_left 2.97438f
C7 plus drain_right 0.461602f
C8 minus plus 5.02172f
C9 source plus 3.4233f
C10 drain_right a_n2982_n1288# 5.39428f
C11 drain_left a_n2982_n1288# 5.83446f
C12 source a_n2982_n1288# 3.51404f
C13 minus a_n2982_n1288# 11.158289f
C14 plus a_n2982_n1288# 12.530611f
C15 drain_right.t8 a_n2982_n1288# 0.042347f
C16 drain_right.t10 a_n2982_n1288# 0.042347f
C17 drain_right.n0 a_n2982_n1288# 0.269261f
C18 drain_right.t4 a_n2982_n1288# 0.042347f
C19 drain_right.t6 a_n2982_n1288# 0.042347f
C20 drain_right.n1 a_n2982_n1288# 0.266037f
C21 drain_right.n2 a_n2982_n1288# 0.72034f
C22 drain_right.t2 a_n2982_n1288# 0.042347f
C23 drain_right.t17 a_n2982_n1288# 0.042347f
C24 drain_right.n3 a_n2982_n1288# 0.266037f
C25 drain_right.t15 a_n2982_n1288# 0.042347f
C26 drain_right.t3 a_n2982_n1288# 0.042347f
C27 drain_right.n4 a_n2982_n1288# 0.269261f
C28 drain_right.t18 a_n2982_n1288# 0.042347f
C29 drain_right.t14 a_n2982_n1288# 0.042347f
C30 drain_right.n5 a_n2982_n1288# 0.266037f
C31 drain_right.n6 a_n2982_n1288# 0.72034f
C32 drain_right.n7 a_n2982_n1288# 1.32282f
C33 drain_right.t19 a_n2982_n1288# 0.042347f
C34 drain_right.t9 a_n2982_n1288# 0.042347f
C35 drain_right.n8 a_n2982_n1288# 0.269262f
C36 drain_right.t1 a_n2982_n1288# 0.042347f
C37 drain_right.t11 a_n2982_n1288# 0.042347f
C38 drain_right.n9 a_n2982_n1288# 0.266038f
C39 drain_right.n10 a_n2982_n1288# 0.72437f
C40 drain_right.t0 a_n2982_n1288# 0.042347f
C41 drain_right.t12 a_n2982_n1288# 0.042347f
C42 drain_right.n11 a_n2982_n1288# 0.266038f
C43 drain_right.n12 a_n2982_n1288# 0.358401f
C44 drain_right.t5 a_n2982_n1288# 0.042347f
C45 drain_right.t13 a_n2982_n1288# 0.042347f
C46 drain_right.n13 a_n2982_n1288# 0.266038f
C47 drain_right.n14 a_n2982_n1288# 0.358401f
C48 drain_right.t7 a_n2982_n1288# 0.042347f
C49 drain_right.t16 a_n2982_n1288# 0.042347f
C50 drain_right.n15 a_n2982_n1288# 0.266038f
C51 drain_right.n16 a_n2982_n1288# 0.595396f
C52 minus.n0 a_n2982_n1288# 0.042166f
C53 minus.n1 a_n2982_n1288# 0.009568f
C54 minus.t3 a_n2982_n1288# 0.182805f
C55 minus.n2 a_n2982_n1288# 0.042166f
C56 minus.n3 a_n2982_n1288# 0.009568f
C57 minus.t6 a_n2982_n1288# 0.182805f
C58 minus.n4 a_n2982_n1288# 0.042166f
C59 minus.n5 a_n2982_n1288# 0.009568f
C60 minus.t7 a_n2982_n1288# 0.182805f
C61 minus.n6 a_n2982_n1288# 0.042166f
C62 minus.n7 a_n2982_n1288# 0.009568f
C63 minus.t8 a_n2982_n1288# 0.182805f
C64 minus.t10 a_n2982_n1288# 0.204338f
C65 minus.t0 a_n2982_n1288# 0.182805f
C66 minus.n8 a_n2982_n1288# 0.134127f
C67 minus.n9 a_n2982_n1288# 0.108569f
C68 minus.n10 a_n2982_n1288# 0.17998f
C69 minus.n11 a_n2982_n1288# 0.042166f
C70 minus.n12 a_n2982_n1288# 0.127074f
C71 minus.n13 a_n2982_n1288# 0.009568f
C72 minus.t18 a_n2982_n1288# 0.182805f
C73 minus.n14 a_n2982_n1288# 0.127074f
C74 minus.n15 a_n2982_n1288# 0.042166f
C75 minus.n16 a_n2982_n1288# 0.042166f
C76 minus.n17 a_n2982_n1288# 0.042166f
C77 minus.n18 a_n2982_n1288# 0.127074f
C78 minus.n19 a_n2982_n1288# 0.009568f
C79 minus.t19 a_n2982_n1288# 0.182805f
C80 minus.n20 a_n2982_n1288# 0.127074f
C81 minus.n21 a_n2982_n1288# 0.042166f
C82 minus.n22 a_n2982_n1288# 0.042166f
C83 minus.n23 a_n2982_n1288# 0.042166f
C84 minus.n24 a_n2982_n1288# 0.127074f
C85 minus.n25 a_n2982_n1288# 0.009568f
C86 minus.t14 a_n2982_n1288# 0.182805f
C87 minus.n26 a_n2982_n1288# 0.127074f
C88 minus.n27 a_n2982_n1288# 0.042166f
C89 minus.n28 a_n2982_n1288# 0.042166f
C90 minus.n29 a_n2982_n1288# 0.042166f
C91 minus.n30 a_n2982_n1288# 0.127074f
C92 minus.n31 a_n2982_n1288# 0.009568f
C93 minus.t12 a_n2982_n1288# 0.182805f
C94 minus.n32 a_n2982_n1288# 0.126684f
C95 minus.n33 a_n2982_n1288# 1.29237f
C96 minus.n34 a_n2982_n1288# 0.042166f
C97 minus.n35 a_n2982_n1288# 0.009568f
C98 minus.n36 a_n2982_n1288# 0.042166f
C99 minus.n37 a_n2982_n1288# 0.009568f
C100 minus.n38 a_n2982_n1288# 0.042166f
C101 minus.n39 a_n2982_n1288# 0.009568f
C102 minus.n40 a_n2982_n1288# 0.042166f
C103 minus.n41 a_n2982_n1288# 0.009568f
C104 minus.t11 a_n2982_n1288# 0.204338f
C105 minus.t9 a_n2982_n1288# 0.182805f
C106 minus.n42 a_n2982_n1288# 0.134127f
C107 minus.n43 a_n2982_n1288# 0.108569f
C108 minus.n44 a_n2982_n1288# 0.17998f
C109 minus.n45 a_n2982_n1288# 0.042166f
C110 minus.t15 a_n2982_n1288# 0.182805f
C111 minus.n46 a_n2982_n1288# 0.127074f
C112 minus.n47 a_n2982_n1288# 0.009568f
C113 minus.t13 a_n2982_n1288# 0.182805f
C114 minus.n48 a_n2982_n1288# 0.127074f
C115 minus.n49 a_n2982_n1288# 0.042166f
C116 minus.n50 a_n2982_n1288# 0.042166f
C117 minus.n51 a_n2982_n1288# 0.042166f
C118 minus.t17 a_n2982_n1288# 0.182805f
C119 minus.n52 a_n2982_n1288# 0.127074f
C120 minus.n53 a_n2982_n1288# 0.009568f
C121 minus.t2 a_n2982_n1288# 0.182805f
C122 minus.n54 a_n2982_n1288# 0.127074f
C123 minus.n55 a_n2982_n1288# 0.042166f
C124 minus.n56 a_n2982_n1288# 0.042166f
C125 minus.n57 a_n2982_n1288# 0.042166f
C126 minus.t1 a_n2982_n1288# 0.182805f
C127 minus.n58 a_n2982_n1288# 0.127074f
C128 minus.n59 a_n2982_n1288# 0.009568f
C129 minus.t5 a_n2982_n1288# 0.182805f
C130 minus.n60 a_n2982_n1288# 0.127074f
C131 minus.n61 a_n2982_n1288# 0.042166f
C132 minus.n62 a_n2982_n1288# 0.042166f
C133 minus.n63 a_n2982_n1288# 0.042166f
C134 minus.t4 a_n2982_n1288# 0.182805f
C135 minus.n64 a_n2982_n1288# 0.127074f
C136 minus.n65 a_n2982_n1288# 0.009568f
C137 minus.t16 a_n2982_n1288# 0.182805f
C138 minus.n66 a_n2982_n1288# 0.126684f
C139 minus.n67 a_n2982_n1288# 0.292145f
C140 minus.n68 a_n2982_n1288# 1.57713f
C141 drain_left.t18 a_n2982_n1288# 0.043157f
C142 drain_left.t19 a_n2982_n1288# 0.043157f
C143 drain_left.n0 a_n2982_n1288# 0.274411f
C144 drain_left.t3 a_n2982_n1288# 0.043157f
C145 drain_left.t8 a_n2982_n1288# 0.043157f
C146 drain_left.n1 a_n2982_n1288# 0.271126f
C147 drain_left.n2 a_n2982_n1288# 0.734117f
C148 drain_left.t6 a_n2982_n1288# 0.043157f
C149 drain_left.t11 a_n2982_n1288# 0.043157f
C150 drain_left.n3 a_n2982_n1288# 0.271126f
C151 drain_left.t2 a_n2982_n1288# 0.043157f
C152 drain_left.t1 a_n2982_n1288# 0.043157f
C153 drain_left.n4 a_n2982_n1288# 0.274411f
C154 drain_left.t10 a_n2982_n1288# 0.043157f
C155 drain_left.t15 a_n2982_n1288# 0.043157f
C156 drain_left.n5 a_n2982_n1288# 0.271126f
C157 drain_left.n6 a_n2982_n1288# 0.734117f
C158 drain_left.n7 a_n2982_n1288# 1.40105f
C159 drain_left.t12 a_n2982_n1288# 0.043157f
C160 drain_left.t4 a_n2982_n1288# 0.043157f
C161 drain_left.n8 a_n2982_n1288# 0.274412f
C162 drain_left.t16 a_n2982_n1288# 0.043157f
C163 drain_left.t7 a_n2982_n1288# 0.043157f
C164 drain_left.n9 a_n2982_n1288# 0.271127f
C165 drain_left.n10 a_n2982_n1288# 0.738225f
C166 drain_left.t13 a_n2982_n1288# 0.043157f
C167 drain_left.t5 a_n2982_n1288# 0.043157f
C168 drain_left.n11 a_n2982_n1288# 0.271127f
C169 drain_left.n12 a_n2982_n1288# 0.365256f
C170 drain_left.t17 a_n2982_n1288# 0.043157f
C171 drain_left.t9 a_n2982_n1288# 0.043157f
C172 drain_left.n13 a_n2982_n1288# 0.271127f
C173 drain_left.n14 a_n2982_n1288# 0.365256f
C174 drain_left.t0 a_n2982_n1288# 0.043157f
C175 drain_left.t14 a_n2982_n1288# 0.043157f
C176 drain_left.n15 a_n2982_n1288# 0.271127f
C177 drain_left.n16 a_n2982_n1288# 0.606784f
C178 source.n0 a_n2982_n1288# 0.045747f
C179 source.n1 a_n2982_n1288# 0.10122f
C180 source.t20 a_n2982_n1288# 0.07596f
C181 source.n2 a_n2982_n1288# 0.079219f
C182 source.n3 a_n2982_n1288# 0.025537f
C183 source.n4 a_n2982_n1288# 0.016842f
C184 source.n5 a_n2982_n1288# 0.223113f
C185 source.n6 a_n2982_n1288# 0.050149f
C186 source.n7 a_n2982_n1288# 0.534925f
C187 source.t39 a_n2982_n1288# 0.049536f
C188 source.t21 a_n2982_n1288# 0.049536f
C189 source.n8 a_n2982_n1288# 0.264817f
C190 source.n9 a_n2982_n1288# 0.423024f
C191 source.t35 a_n2982_n1288# 0.049536f
C192 source.t25 a_n2982_n1288# 0.049536f
C193 source.n10 a_n2982_n1288# 0.264817f
C194 source.n11 a_n2982_n1288# 0.423024f
C195 source.t36 a_n2982_n1288# 0.049536f
C196 source.t31 a_n2982_n1288# 0.049536f
C197 source.n12 a_n2982_n1288# 0.264817f
C198 source.n13 a_n2982_n1288# 0.423024f
C199 source.t37 a_n2982_n1288# 0.049536f
C200 source.t24 a_n2982_n1288# 0.049536f
C201 source.n14 a_n2982_n1288# 0.264817f
C202 source.n15 a_n2982_n1288# 0.423024f
C203 source.n16 a_n2982_n1288# 0.045747f
C204 source.n17 a_n2982_n1288# 0.10122f
C205 source.t34 a_n2982_n1288# 0.07596f
C206 source.n18 a_n2982_n1288# 0.079219f
C207 source.n19 a_n2982_n1288# 0.025537f
C208 source.n20 a_n2982_n1288# 0.016842f
C209 source.n21 a_n2982_n1288# 0.223113f
C210 source.n22 a_n2982_n1288# 0.050149f
C211 source.n23 a_n2982_n1288# 0.162927f
C212 source.n24 a_n2982_n1288# 0.045747f
C213 source.n25 a_n2982_n1288# 0.10122f
C214 source.t15 a_n2982_n1288# 0.07596f
C215 source.n26 a_n2982_n1288# 0.079219f
C216 source.n27 a_n2982_n1288# 0.025537f
C217 source.n28 a_n2982_n1288# 0.016842f
C218 source.n29 a_n2982_n1288# 0.223113f
C219 source.n30 a_n2982_n1288# 0.050149f
C220 source.n31 a_n2982_n1288# 0.162927f
C221 source.t6 a_n2982_n1288# 0.049536f
C222 source.t2 a_n2982_n1288# 0.049536f
C223 source.n32 a_n2982_n1288# 0.264817f
C224 source.n33 a_n2982_n1288# 0.423024f
C225 source.t18 a_n2982_n1288# 0.049536f
C226 source.t8 a_n2982_n1288# 0.049536f
C227 source.n34 a_n2982_n1288# 0.264817f
C228 source.n35 a_n2982_n1288# 0.423024f
C229 source.t16 a_n2982_n1288# 0.049536f
C230 source.t11 a_n2982_n1288# 0.049536f
C231 source.n36 a_n2982_n1288# 0.264817f
C232 source.n37 a_n2982_n1288# 0.423024f
C233 source.t4 a_n2982_n1288# 0.049536f
C234 source.t19 a_n2982_n1288# 0.049536f
C235 source.n38 a_n2982_n1288# 0.264817f
C236 source.n39 a_n2982_n1288# 0.423024f
C237 source.n40 a_n2982_n1288# 0.045747f
C238 source.n41 a_n2982_n1288# 0.10122f
C239 source.t14 a_n2982_n1288# 0.07596f
C240 source.n42 a_n2982_n1288# 0.079219f
C241 source.n43 a_n2982_n1288# 0.025537f
C242 source.n44 a_n2982_n1288# 0.016842f
C243 source.n45 a_n2982_n1288# 0.223113f
C244 source.n46 a_n2982_n1288# 0.050149f
C245 source.n47 a_n2982_n1288# 0.835082f
C246 source.n48 a_n2982_n1288# 0.045747f
C247 source.n49 a_n2982_n1288# 0.10122f
C248 source.t30 a_n2982_n1288# 0.07596f
C249 source.n50 a_n2982_n1288# 0.079219f
C250 source.n51 a_n2982_n1288# 0.025537f
C251 source.n52 a_n2982_n1288# 0.016842f
C252 source.n53 a_n2982_n1288# 0.223113f
C253 source.n54 a_n2982_n1288# 0.050149f
C254 source.n55 a_n2982_n1288# 0.835082f
C255 source.t29 a_n2982_n1288# 0.049536f
C256 source.t27 a_n2982_n1288# 0.049536f
C257 source.n56 a_n2982_n1288# 0.264816f
C258 source.n57 a_n2982_n1288# 0.423026f
C259 source.t33 a_n2982_n1288# 0.049536f
C260 source.t28 a_n2982_n1288# 0.049536f
C261 source.n58 a_n2982_n1288# 0.264816f
C262 source.n59 a_n2982_n1288# 0.423026f
C263 source.t22 a_n2982_n1288# 0.049536f
C264 source.t23 a_n2982_n1288# 0.049536f
C265 source.n60 a_n2982_n1288# 0.264816f
C266 source.n61 a_n2982_n1288# 0.423026f
C267 source.t26 a_n2982_n1288# 0.049536f
C268 source.t38 a_n2982_n1288# 0.049536f
C269 source.n62 a_n2982_n1288# 0.264816f
C270 source.n63 a_n2982_n1288# 0.423026f
C271 source.n64 a_n2982_n1288# 0.045747f
C272 source.n65 a_n2982_n1288# 0.10122f
C273 source.t32 a_n2982_n1288# 0.07596f
C274 source.n66 a_n2982_n1288# 0.079219f
C275 source.n67 a_n2982_n1288# 0.025537f
C276 source.n68 a_n2982_n1288# 0.016842f
C277 source.n69 a_n2982_n1288# 0.223113f
C278 source.n70 a_n2982_n1288# 0.050149f
C279 source.n71 a_n2982_n1288# 0.162927f
C280 source.n72 a_n2982_n1288# 0.045747f
C281 source.n73 a_n2982_n1288# 0.10122f
C282 source.t3 a_n2982_n1288# 0.07596f
C283 source.n74 a_n2982_n1288# 0.079219f
C284 source.n75 a_n2982_n1288# 0.025537f
C285 source.n76 a_n2982_n1288# 0.016842f
C286 source.n77 a_n2982_n1288# 0.223113f
C287 source.n78 a_n2982_n1288# 0.050149f
C288 source.n79 a_n2982_n1288# 0.162927f
C289 source.t12 a_n2982_n1288# 0.049536f
C290 source.t10 a_n2982_n1288# 0.049536f
C291 source.n80 a_n2982_n1288# 0.264816f
C292 source.n81 a_n2982_n1288# 0.423026f
C293 source.t7 a_n2982_n1288# 0.049536f
C294 source.t17 a_n2982_n1288# 0.049536f
C295 source.n82 a_n2982_n1288# 0.264816f
C296 source.n83 a_n2982_n1288# 0.423026f
C297 source.t1 a_n2982_n1288# 0.049536f
C298 source.t0 a_n2982_n1288# 0.049536f
C299 source.n84 a_n2982_n1288# 0.264816f
C300 source.n85 a_n2982_n1288# 0.423026f
C301 source.t5 a_n2982_n1288# 0.049536f
C302 source.t9 a_n2982_n1288# 0.049536f
C303 source.n86 a_n2982_n1288# 0.264816f
C304 source.n87 a_n2982_n1288# 0.423026f
C305 source.n88 a_n2982_n1288# 0.045747f
C306 source.n89 a_n2982_n1288# 0.10122f
C307 source.t13 a_n2982_n1288# 0.07596f
C308 source.n90 a_n2982_n1288# 0.079219f
C309 source.n91 a_n2982_n1288# 0.025537f
C310 source.n92 a_n2982_n1288# 0.016842f
C311 source.n93 a_n2982_n1288# 0.223113f
C312 source.n94 a_n2982_n1288# 0.050149f
C313 source.n95 a_n2982_n1288# 0.367376f
C314 source.n96 a_n2982_n1288# 0.790157f
C315 plus.n0 a_n2982_n1288# 0.04364f
C316 plus.t5 a_n2982_n1288# 0.1892f
C317 plus.t19 a_n2982_n1288# 0.1892f
C318 plus.n1 a_n2982_n1288# 0.04364f
C319 plus.t10 a_n2982_n1288# 0.1892f
C320 plus.n2 a_n2982_n1288# 0.131519f
C321 plus.n3 a_n2982_n1288# 0.04364f
C322 plus.t2 a_n2982_n1288# 0.1892f
C323 plus.t14 a_n2982_n1288# 0.1892f
C324 plus.n4 a_n2982_n1288# 0.131519f
C325 plus.n5 a_n2982_n1288# 0.04364f
C326 plus.t6 a_n2982_n1288# 0.1892f
C327 plus.t12 a_n2982_n1288# 0.1892f
C328 plus.n6 a_n2982_n1288# 0.131519f
C329 plus.n7 a_n2982_n1288# 0.04364f
C330 plus.t3 a_n2982_n1288# 0.1892f
C331 plus.t15 a_n2982_n1288# 0.1892f
C332 plus.n8 a_n2982_n1288# 0.138818f
C333 plus.t7 a_n2982_n1288# 0.211485f
C334 plus.n9 a_n2982_n1288# 0.112367f
C335 plus.n10 a_n2982_n1288# 0.186275f
C336 plus.n11 a_n2982_n1288# 0.009903f
C337 plus.n12 a_n2982_n1288# 0.131519f
C338 plus.n13 a_n2982_n1288# 0.009903f
C339 plus.n14 a_n2982_n1288# 0.04364f
C340 plus.n15 a_n2982_n1288# 0.04364f
C341 plus.n16 a_n2982_n1288# 0.04364f
C342 plus.n17 a_n2982_n1288# 0.009903f
C343 plus.n18 a_n2982_n1288# 0.131519f
C344 plus.n19 a_n2982_n1288# 0.009903f
C345 plus.n20 a_n2982_n1288# 0.04364f
C346 plus.n21 a_n2982_n1288# 0.04364f
C347 plus.n22 a_n2982_n1288# 0.04364f
C348 plus.n23 a_n2982_n1288# 0.009903f
C349 plus.n24 a_n2982_n1288# 0.131519f
C350 plus.n25 a_n2982_n1288# 0.009903f
C351 plus.n26 a_n2982_n1288# 0.04364f
C352 plus.n27 a_n2982_n1288# 0.04364f
C353 plus.n28 a_n2982_n1288# 0.04364f
C354 plus.n29 a_n2982_n1288# 0.009903f
C355 plus.n30 a_n2982_n1288# 0.131519f
C356 plus.n31 a_n2982_n1288# 0.009903f
C357 plus.n32 a_n2982_n1288# 0.131115f
C358 plus.n33 a_n2982_n1288# 0.32997f
C359 plus.n34 a_n2982_n1288# 0.04364f
C360 plus.t1 a_n2982_n1288# 0.1892f
C361 plus.n35 a_n2982_n1288# 0.04364f
C362 plus.t0 a_n2982_n1288# 0.1892f
C363 plus.t16 a_n2982_n1288# 0.1892f
C364 plus.n36 a_n2982_n1288# 0.131519f
C365 plus.n37 a_n2982_n1288# 0.04364f
C366 plus.t11 a_n2982_n1288# 0.1892f
C367 plus.t13 a_n2982_n1288# 0.1892f
C368 plus.n38 a_n2982_n1288# 0.131519f
C369 plus.n39 a_n2982_n1288# 0.04364f
C370 plus.t8 a_n2982_n1288# 0.1892f
C371 plus.t9 a_n2982_n1288# 0.1892f
C372 plus.n40 a_n2982_n1288# 0.131519f
C373 plus.n41 a_n2982_n1288# 0.04364f
C374 plus.t4 a_n2982_n1288# 0.1892f
C375 plus.t17 a_n2982_n1288# 0.1892f
C376 plus.n42 a_n2982_n1288# 0.138818f
C377 plus.t18 a_n2982_n1288# 0.211485f
C378 plus.n43 a_n2982_n1288# 0.112367f
C379 plus.n44 a_n2982_n1288# 0.186275f
C380 plus.n45 a_n2982_n1288# 0.009903f
C381 plus.n46 a_n2982_n1288# 0.131519f
C382 plus.n47 a_n2982_n1288# 0.009903f
C383 plus.n48 a_n2982_n1288# 0.04364f
C384 plus.n49 a_n2982_n1288# 0.04364f
C385 plus.n50 a_n2982_n1288# 0.04364f
C386 plus.n51 a_n2982_n1288# 0.009903f
C387 plus.n52 a_n2982_n1288# 0.131519f
C388 plus.n53 a_n2982_n1288# 0.009903f
C389 plus.n54 a_n2982_n1288# 0.04364f
C390 plus.n55 a_n2982_n1288# 0.04364f
C391 plus.n56 a_n2982_n1288# 0.04364f
C392 plus.n57 a_n2982_n1288# 0.009903f
C393 plus.n58 a_n2982_n1288# 0.131519f
C394 plus.n59 a_n2982_n1288# 0.009903f
C395 plus.n60 a_n2982_n1288# 0.04364f
C396 plus.n61 a_n2982_n1288# 0.04364f
C397 plus.n62 a_n2982_n1288# 0.04364f
C398 plus.n63 a_n2982_n1288# 0.009903f
C399 plus.n64 a_n2982_n1288# 0.131519f
C400 plus.n65 a_n2982_n1288# 0.009903f
C401 plus.n66 a_n2982_n1288# 0.131115f
C402 plus.n67 a_n2982_n1288# 1.27156f
.ends

