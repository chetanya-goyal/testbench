* NGSPICE file created from diffpair204.ext - technology: sky130A

.subckt diffpair204 minus drain_right drain_left source plus
X0 a_n1712_n1488# a_n1712_n1488# a_n1712_n1488# a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.5
X1 drain_right.t9 minus.t0 source.t9 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X2 source.t16 minus.t1 drain_right.t8 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X3 drain_left.t9 plus.t0 source.t1 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X4 drain_left.t8 plus.t1 source.t0 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X5 drain_right.t7 minus.t2 source.t7 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X6 drain_right.t6 minus.t3 source.t14 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X7 source.t13 minus.t4 drain_right.t5 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X8 drain_left.t7 plus.t2 source.t17 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X9 drain_right.t4 minus.t5 source.t12 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X10 source.t18 plus.t3 drain_left.t6 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X11 source.t10 minus.t6 drain_right.t3 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X12 source.t19 plus.t4 drain_left.t5 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X13 a_n1712_n1488# a_n1712_n1488# a_n1712_n1488# a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X14 a_n1712_n1488# a_n1712_n1488# a_n1712_n1488# a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X15 source.t5 plus.t5 drain_left.t4 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X16 drain_right.t2 minus.t7 source.t8 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X17 source.t4 plus.t6 drain_left.t3 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X18 drain_right.t1 minus.t8 source.t11 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X19 source.t15 minus.t9 drain_right.t0 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
X20 drain_left.t2 plus.t7 source.t6 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.5
X21 drain_left.t1 plus.t8 source.t2 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.5
X22 a_n1712_n1488# a_n1712_n1488# a_n1712_n1488# a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X23 drain_left.t0 plus.t9 source.t3 a_n1712_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.5
R0 minus.n2 minus.t7 244.149
R1 minus.n14 minus.t2 244.149
R2 minus.n3 minus.t1 223.167
R3 minus.n1 minus.t5 223.167
R4 minus.n9 minus.t9 223.167
R5 minus.n10 minus.t3 223.167
R6 minus.n15 minus.t6 223.167
R7 minus.n13 minus.t0 223.167
R8 minus.n21 minus.t4 223.167
R9 minus.n22 minus.t8 223.167
R10 minus.n11 minus.n10 161.3
R11 minus.n9 minus.n0 161.3
R12 minus.n8 minus.n7 161.3
R13 minus.n6 minus.n1 161.3
R14 minus.n5 minus.n4 161.3
R15 minus.n23 minus.n22 161.3
R16 minus.n21 minus.n12 161.3
R17 minus.n20 minus.n19 161.3
R18 minus.n18 minus.n13 161.3
R19 minus.n17 minus.n16 161.3
R20 minus.n5 minus.n2 70.4033
R21 minus.n17 minus.n14 70.4033
R22 minus.n10 minus.n9 48.2005
R23 minus.n22 minus.n21 48.2005
R24 minus.n4 minus.n1 36.5157
R25 minus.n8 minus.n1 36.5157
R26 minus.n16 minus.n13 36.5157
R27 minus.n20 minus.n13 36.5157
R28 minus.n24 minus.n11 28.8509
R29 minus.n3 minus.n2 20.9576
R30 minus.n15 minus.n14 20.9576
R31 minus.n4 minus.n3 11.6853
R32 minus.n9 minus.n8 11.6853
R33 minus.n16 minus.n15 11.6853
R34 minus.n21 minus.n20 11.6853
R35 minus.n24 minus.n23 6.563
R36 minus.n11 minus.n0 0.189894
R37 minus.n7 minus.n0 0.189894
R38 minus.n7 minus.n6 0.189894
R39 minus.n6 minus.n5 0.189894
R40 minus.n18 minus.n17 0.189894
R41 minus.n19 minus.n18 0.189894
R42 minus.n19 minus.n12 0.189894
R43 minus.n23 minus.n12 0.189894
R44 minus minus.n24 0.188
R45 source.n0 source.t2 69.6943
R46 source.n5 source.t8 69.6943
R47 source.n19 source.t11 69.6942
R48 source.n14 source.t17 69.6942
R49 source.n2 source.n1 63.0943
R50 source.n4 source.n3 63.0943
R51 source.n7 source.n6 63.0943
R52 source.n9 source.n8 63.0943
R53 source.n18 source.n17 63.0942
R54 source.n16 source.n15 63.0942
R55 source.n13 source.n12 63.0942
R56 source.n11 source.n10 63.0942
R57 source.n11 source.n9 15.9006
R58 source.n20 source.n0 9.56437
R59 source.n17 source.t9 6.6005
R60 source.n17 source.t13 6.6005
R61 source.n15 source.t7 6.6005
R62 source.n15 source.t10 6.6005
R63 source.n12 source.t1 6.6005
R64 source.n12 source.t19 6.6005
R65 source.n10 source.t6 6.6005
R66 source.n10 source.t5 6.6005
R67 source.n1 source.t3 6.6005
R68 source.n1 source.t18 6.6005
R69 source.n3 source.t0 6.6005
R70 source.n3 source.t4 6.6005
R71 source.n6 source.t12 6.6005
R72 source.n6 source.t16 6.6005
R73 source.n8 source.t14 6.6005
R74 source.n8 source.t15 6.6005
R75 source.n20 source.n19 5.62119
R76 source.n5 source.n4 0.828086
R77 source.n16 source.n14 0.828086
R78 source.n9 source.n7 0.716017
R79 source.n7 source.n5 0.716017
R80 source.n4 source.n2 0.716017
R81 source.n2 source.n0 0.716017
R82 source.n13 source.n11 0.716017
R83 source.n14 source.n13 0.716017
R84 source.n18 source.n16 0.716017
R85 source.n19 source.n18 0.716017
R86 source source.n20 0.188
R87 drain_right.n1 drain_right.t7 87.0885
R88 drain_right.n7 drain_right.t6 86.3731
R89 drain_right.n6 drain_right.n4 80.4886
R90 drain_right.n3 drain_right.n2 80.2543
R91 drain_right.n6 drain_right.n5 79.7731
R92 drain_right.n1 drain_right.n0 79.773
R93 drain_right drain_right.n3 23.0366
R94 drain_right.n2 drain_right.t5 6.6005
R95 drain_right.n2 drain_right.t1 6.6005
R96 drain_right.n0 drain_right.t3 6.6005
R97 drain_right.n0 drain_right.t9 6.6005
R98 drain_right.n4 drain_right.t8 6.6005
R99 drain_right.n4 drain_right.t2 6.6005
R100 drain_right.n5 drain_right.t0 6.6005
R101 drain_right.n5 drain_right.t4 6.6005
R102 drain_right drain_right.n7 6.01097
R103 drain_right.n7 drain_right.n6 0.716017
R104 drain_right.n3 drain_right.n1 0.124033
R105 plus.n2 plus.t1 244.149
R106 plus.n14 plus.t2 244.149
R107 plus.n10 plus.t8 223.167
R108 plus.n9 plus.t3 223.167
R109 plus.n1 plus.t9 223.167
R110 plus.n3 plus.t6 223.167
R111 plus.n22 plus.t7 223.167
R112 plus.n21 plus.t5 223.167
R113 plus.n13 plus.t0 223.167
R114 plus.n15 plus.t4 223.167
R115 plus.n5 plus.n4 161.3
R116 plus.n6 plus.n1 161.3
R117 plus.n8 plus.n7 161.3
R118 plus.n9 plus.n0 161.3
R119 plus.n11 plus.n10 161.3
R120 plus.n17 plus.n16 161.3
R121 plus.n18 plus.n13 161.3
R122 plus.n20 plus.n19 161.3
R123 plus.n21 plus.n12 161.3
R124 plus.n23 plus.n22 161.3
R125 plus.n5 plus.n2 70.4033
R126 plus.n17 plus.n14 70.4033
R127 plus.n10 plus.n9 48.2005
R128 plus.n22 plus.n21 48.2005
R129 plus.n8 plus.n1 36.5157
R130 plus.n4 plus.n1 36.5157
R131 plus.n20 plus.n13 36.5157
R132 plus.n16 plus.n13 36.5157
R133 plus plus.n23 26.1411
R134 plus.n3 plus.n2 20.9576
R135 plus.n15 plus.n14 20.9576
R136 plus.n9 plus.n8 11.6853
R137 plus.n4 plus.n3 11.6853
R138 plus.n21 plus.n20 11.6853
R139 plus.n16 plus.n15 11.6853
R140 plus plus.n11 8.79785
R141 plus.n6 plus.n5 0.189894
R142 plus.n7 plus.n6 0.189894
R143 plus.n7 plus.n0 0.189894
R144 plus.n11 plus.n0 0.189894
R145 plus.n23 plus.n12 0.189894
R146 plus.n19 plus.n12 0.189894
R147 plus.n19 plus.n18 0.189894
R148 plus.n18 plus.n17 0.189894
R149 drain_left.n5 drain_left.t8 87.0886
R150 drain_left.n1 drain_left.t2 87.0885
R151 drain_left.n3 drain_left.n2 80.2543
R152 drain_left.n7 drain_left.n6 79.7731
R153 drain_left.n5 drain_left.n4 79.7731
R154 drain_left.n1 drain_left.n0 79.773
R155 drain_left drain_left.n3 23.5898
R156 drain_left.n2 drain_left.t5 6.6005
R157 drain_left.n2 drain_left.t7 6.6005
R158 drain_left.n0 drain_left.t4 6.6005
R159 drain_left.n0 drain_left.t9 6.6005
R160 drain_left.n6 drain_left.t6 6.6005
R161 drain_left.n6 drain_left.t1 6.6005
R162 drain_left.n4 drain_left.t3 6.6005
R163 drain_left.n4 drain_left.t0 6.6005
R164 drain_left drain_left.n7 6.36873
R165 drain_left.n7 drain_left.n5 0.716017
R166 drain_left.n3 drain_left.n1 0.124033
C0 plus drain_left 1.86202f
C1 minus source 1.87353f
C2 plus source 1.88767f
C3 drain_left source 5.93325f
C4 drain_right minus 1.6974f
C5 plus drain_right 0.326279f
C6 drain_right drain_left 0.843971f
C7 drain_right source 5.93099f
C8 plus minus 3.62235f
C9 minus drain_left 0.176946f
C10 drain_right a_n1712_n1488# 3.8739f
C11 drain_left a_n1712_n1488# 4.1077f
C12 source a_n1712_n1488# 2.919983f
C13 minus a_n1712_n1488# 5.931834f
C14 plus a_n1712_n1488# 6.476689f
C15 drain_left.t2 a_n1712_n1488# 0.431603f
C16 drain_left.t4 a_n1712_n1488# 0.046415f
C17 drain_left.t9 a_n1712_n1488# 0.046415f
C18 drain_left.n0 a_n1712_n1488# 0.334738f
C19 drain_left.n1 a_n1712_n1488# 0.452799f
C20 drain_left.t5 a_n1712_n1488# 0.046415f
C21 drain_left.t7 a_n1712_n1488# 0.046415f
C22 drain_left.n2 a_n1712_n1488# 0.336184f
C23 drain_left.n3 a_n1712_n1488# 0.813848f
C24 drain_left.t8 a_n1712_n1488# 0.431604f
C25 drain_left.t3 a_n1712_n1488# 0.046415f
C26 drain_left.t0 a_n1712_n1488# 0.046415f
C27 drain_left.n4 a_n1712_n1488# 0.33474f
C28 drain_left.n5 a_n1712_n1488# 0.486468f
C29 drain_left.t6 a_n1712_n1488# 0.046415f
C30 drain_left.t1 a_n1712_n1488# 0.046415f
C31 drain_left.n6 a_n1712_n1488# 0.33474f
C32 drain_left.n7 a_n1712_n1488# 0.415208f
C33 plus.n0 a_n1712_n1488# 0.024757f
C34 plus.t8 a_n1712_n1488# 0.111358f
C35 plus.t3 a_n1712_n1488# 0.111358f
C36 plus.t9 a_n1712_n1488# 0.111358f
C37 plus.n1 a_n1712_n1488# 0.069385f
C38 plus.t1 a_n1712_n1488# 0.117101f
C39 plus.n2 a_n1712_n1488# 0.061228f
C40 plus.t6 a_n1712_n1488# 0.111358f
C41 plus.n3 a_n1712_n1488# 0.068011f
C42 plus.n4 a_n1712_n1488# 0.005618f
C43 plus.n5 a_n1712_n1488# 0.078976f
C44 plus.n6 a_n1712_n1488# 0.024757f
C45 plus.n7 a_n1712_n1488# 0.024757f
C46 plus.n8 a_n1712_n1488# 0.005618f
C47 plus.n9 a_n1712_n1488# 0.068011f
C48 plus.n10 a_n1712_n1488# 0.06679f
C49 plus.n11 a_n1712_n1488# 0.188793f
C50 plus.n12 a_n1712_n1488# 0.024757f
C51 plus.t7 a_n1712_n1488# 0.111358f
C52 plus.t5 a_n1712_n1488# 0.111358f
C53 plus.t0 a_n1712_n1488# 0.111358f
C54 plus.n13 a_n1712_n1488# 0.069385f
C55 plus.t2 a_n1712_n1488# 0.117101f
C56 plus.n14 a_n1712_n1488# 0.061228f
C57 plus.t4 a_n1712_n1488# 0.111358f
C58 plus.n15 a_n1712_n1488# 0.068011f
C59 plus.n16 a_n1712_n1488# 0.005618f
C60 plus.n17 a_n1712_n1488# 0.078976f
C61 plus.n18 a_n1712_n1488# 0.024757f
C62 plus.n19 a_n1712_n1488# 0.024757f
C63 plus.n20 a_n1712_n1488# 0.005618f
C64 plus.n21 a_n1712_n1488# 0.068011f
C65 plus.n22 a_n1712_n1488# 0.06679f
C66 plus.n23 a_n1712_n1488# 0.568459f
C67 drain_right.t7 a_n1712_n1488# 0.437279f
C68 drain_right.t3 a_n1712_n1488# 0.047025f
C69 drain_right.t9 a_n1712_n1488# 0.047025f
C70 drain_right.n0 a_n1712_n1488# 0.33914f
C71 drain_right.n1 a_n1712_n1488# 0.458755f
C72 drain_right.t5 a_n1712_n1488# 0.047025f
C73 drain_right.t1 a_n1712_n1488# 0.047025f
C74 drain_right.n2 a_n1712_n1488# 0.340605f
C75 drain_right.n3 a_n1712_n1488# 0.785178f
C76 drain_right.t8 a_n1712_n1488# 0.047025f
C77 drain_right.t2 a_n1712_n1488# 0.047025f
C78 drain_right.n4 a_n1712_n1488# 0.341438f
C79 drain_right.t0 a_n1712_n1488# 0.047025f
C80 drain_right.t4 a_n1712_n1488# 0.047025f
C81 drain_right.n5 a_n1712_n1488# 0.339142f
C82 drain_right.n6 a_n1712_n1488# 0.506192f
C83 drain_right.t6 a_n1712_n1488# 0.435271f
C84 drain_right.n7 a_n1712_n1488# 0.418562f
C85 source.t2 a_n1712_n1488# 0.459505f
C86 source.n0 a_n1712_n1488# 0.649728f
C87 source.t3 a_n1712_n1488# 0.055337f
C88 source.t18 a_n1712_n1488# 0.055337f
C89 source.n1 a_n1712_n1488# 0.350866f
C90 source.n2 a_n1712_n1488# 0.310971f
C91 source.t0 a_n1712_n1488# 0.055337f
C92 source.t4 a_n1712_n1488# 0.055337f
C93 source.n3 a_n1712_n1488# 0.350866f
C94 source.n4 a_n1712_n1488# 0.3194f
C95 source.t8 a_n1712_n1488# 0.459505f
C96 source.n5 a_n1712_n1488# 0.361679f
C97 source.t12 a_n1712_n1488# 0.055337f
C98 source.t16 a_n1712_n1488# 0.055337f
C99 source.n6 a_n1712_n1488# 0.350866f
C100 source.n7 a_n1712_n1488# 0.310971f
C101 source.t14 a_n1712_n1488# 0.055337f
C102 source.t15 a_n1712_n1488# 0.055337f
C103 source.n8 a_n1712_n1488# 0.350866f
C104 source.n9 a_n1712_n1488# 0.907701f
C105 source.t6 a_n1712_n1488# 0.055337f
C106 source.t5 a_n1712_n1488# 0.055337f
C107 source.n10 a_n1712_n1488# 0.350863f
C108 source.n11 a_n1712_n1488# 0.907703f
C109 source.t1 a_n1712_n1488# 0.055337f
C110 source.t19 a_n1712_n1488# 0.055337f
C111 source.n12 a_n1712_n1488# 0.350863f
C112 source.n13 a_n1712_n1488# 0.310974f
C113 source.t17 a_n1712_n1488# 0.459503f
C114 source.n14 a_n1712_n1488# 0.361681f
C115 source.t7 a_n1712_n1488# 0.055337f
C116 source.t10 a_n1712_n1488# 0.055337f
C117 source.n15 a_n1712_n1488# 0.350863f
C118 source.n16 a_n1712_n1488# 0.319403f
C119 source.t9 a_n1712_n1488# 0.055337f
C120 source.t13 a_n1712_n1488# 0.055337f
C121 source.n17 a_n1712_n1488# 0.350863f
C122 source.n18 a_n1712_n1488# 0.310974f
C123 source.t11 a_n1712_n1488# 0.459503f
C124 source.n19 a_n1712_n1488# 0.476844f
C125 source.n20 a_n1712_n1488# 0.68236f
C126 minus.n0 a_n1712_n1488# 0.024418f
C127 minus.t5 a_n1712_n1488# 0.109831f
C128 minus.n1 a_n1712_n1488# 0.068433f
C129 minus.t7 a_n1712_n1488# 0.115495f
C130 minus.n2 a_n1712_n1488# 0.060388f
C131 minus.t1 a_n1712_n1488# 0.109831f
C132 minus.n3 a_n1712_n1488# 0.067078f
C133 minus.n4 a_n1712_n1488# 0.005541f
C134 minus.n5 a_n1712_n1488# 0.077893f
C135 minus.n6 a_n1712_n1488# 0.024418f
C136 minus.n7 a_n1712_n1488# 0.024418f
C137 minus.n8 a_n1712_n1488# 0.005541f
C138 minus.t9 a_n1712_n1488# 0.109831f
C139 minus.n9 a_n1712_n1488# 0.067078f
C140 minus.t3 a_n1712_n1488# 0.109831f
C141 minus.n10 a_n1712_n1488# 0.065874f
C142 minus.n11 a_n1712_n1488# 0.595319f
C143 minus.n12 a_n1712_n1488# 0.024418f
C144 minus.t0 a_n1712_n1488# 0.109831f
C145 minus.n13 a_n1712_n1488# 0.068433f
C146 minus.t2 a_n1712_n1488# 0.115495f
C147 minus.n14 a_n1712_n1488# 0.060388f
C148 minus.t6 a_n1712_n1488# 0.109831f
C149 minus.n15 a_n1712_n1488# 0.067078f
C150 minus.n16 a_n1712_n1488# 0.005541f
C151 minus.n17 a_n1712_n1488# 0.077893f
C152 minus.n18 a_n1712_n1488# 0.024418f
C153 minus.n19 a_n1712_n1488# 0.024418f
C154 minus.n20 a_n1712_n1488# 0.005541f
C155 minus.t4 a_n1712_n1488# 0.109831f
C156 minus.n21 a_n1712_n1488# 0.067078f
C157 minus.t8 a_n1712_n1488# 0.109831f
C158 minus.n22 a_n1712_n1488# 0.065874f
C159 minus.n23 a_n1712_n1488# 0.163252f
C160 minus.n24 a_n1712_n1488# 0.733597f
.ends

