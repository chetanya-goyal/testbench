* NGSPICE file created from diffpair115.ext - technology: sky130A

.subckt diffpair115 minus drain_right drain_left source plus
X0 source.t22 minus.t0 drain_right.t9 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X1 source.t1 plus.t0 drain_left.t11 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X2 source.t21 minus.t1 drain_right.t3 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X3 drain_right.t10 minus.t2 source.t20 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X4 drain_right.t0 minus.t3 source.t19 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X5 a_n1598_n1288# a_n1598_n1288# a_n1598_n1288# a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.3
X6 source.t0 plus.t1 drain_left.t10 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X7 a_n1598_n1288# a_n1598_n1288# a_n1598_n1288# a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X8 a_n1598_n1288# a_n1598_n1288# a_n1598_n1288# a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X9 drain_left.t9 plus.t2 source.t3 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X10 source.t7 plus.t3 drain_left.t8 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X11 drain_left.t7 plus.t4 source.t9 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X12 source.t18 minus.t4 drain_right.t4 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X13 source.t8 plus.t5 drain_left.t6 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X14 source.t17 minus.t5 drain_right.t5 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X15 source.t2 plus.t6 drain_left.t5 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X16 drain_right.t7 minus.t6 source.t16 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X17 drain_left.t4 plus.t7 source.t5 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X18 drain_right.t8 minus.t7 source.t15 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X19 drain_right.t1 minus.t8 source.t14 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X20 drain_left.t3 plus.t8 source.t6 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X21 source.t10 plus.t9 drain_left.t2 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X22 a_n1598_n1288# a_n1598_n1288# a_n1598_n1288# a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X23 source.t13 minus.t9 drain_right.t6 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X24 drain_right.t11 minus.t10 source.t12 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X25 source.t11 minus.t11 drain_right.t2 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X26 drain_left.t1 plus.t10 source.t4 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X27 drain_left.t0 plus.t11 source.t23 a_n1598_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
R0 minus.n13 minus.t1 312.57
R1 minus.n2 minus.t6 312.57
R2 minus.n28 minus.t7 312.57
R3 minus.n17 minus.t0 312.57
R4 minus.n12 minus.t10 265.101
R5 minus.n10 minus.t5 265.101
R6 minus.n3 minus.t2 265.101
R7 minus.n4 minus.t11 265.101
R8 minus.n27 minus.t9 265.101
R9 minus.n25 minus.t3 265.101
R10 minus.n19 minus.t4 265.101
R11 minus.n18 minus.t8 265.101
R12 minus.n6 minus.n2 161.489
R13 minus.n21 minus.n17 161.489
R14 minus.n14 minus.n13 161.3
R15 minus.n11 minus.n0 161.3
R16 minus.n9 minus.n8 161.3
R17 minus.n7 minus.n1 161.3
R18 minus.n6 minus.n5 161.3
R19 minus.n29 minus.n28 161.3
R20 minus.n26 minus.n15 161.3
R21 minus.n24 minus.n23 161.3
R22 minus.n22 minus.n16 161.3
R23 minus.n21 minus.n20 161.3
R24 minus.n9 minus.n1 73.0308
R25 minus.n24 minus.n16 73.0308
R26 minus.n11 minus.n10 63.5369
R27 minus.n5 minus.n3 63.5369
R28 minus.n20 minus.n19 63.5369
R29 minus.n26 minus.n25 63.5369
R30 minus.n13 minus.n12 44.549
R31 minus.n4 minus.n2 44.549
R32 minus.n18 minus.n17 44.549
R33 minus.n28 minus.n27 44.549
R34 minus.n12 minus.n11 28.4823
R35 minus.n5 minus.n4 28.4823
R36 minus.n20 minus.n18 28.4823
R37 minus.n27 minus.n26 28.4823
R38 minus.n30 minus.n14 27.6103
R39 minus.n10 minus.n9 9.49444
R40 minus.n3 minus.n1 9.49444
R41 minus.n19 minus.n16 9.49444
R42 minus.n25 minus.n24 9.49444
R43 minus.n30 minus.n29 6.51186
R44 minus.n14 minus.n0 0.189894
R45 minus.n8 minus.n0 0.189894
R46 minus.n8 minus.n7 0.189894
R47 minus.n7 minus.n6 0.189894
R48 minus.n22 minus.n21 0.189894
R49 minus.n23 minus.n22 0.189894
R50 minus.n23 minus.n15 0.189894
R51 minus.n29 minus.n15 0.189894
R52 minus minus.n30 0.188
R53 drain_right.n6 drain_right.n4 101.338
R54 drain_right.n3 drain_right.n2 101.284
R55 drain_right.n3 drain_right.n0 101.284
R56 drain_right.n6 drain_right.n5 100.796
R57 drain_right.n8 drain_right.n7 100.796
R58 drain_right.n3 drain_right.n1 100.796
R59 drain_right drain_right.n3 21.9536
R60 drain_right.n1 drain_right.t4 9.9005
R61 drain_right.n1 drain_right.t0 9.9005
R62 drain_right.n2 drain_right.t6 9.9005
R63 drain_right.n2 drain_right.t8 9.9005
R64 drain_right.n0 drain_right.t9 9.9005
R65 drain_right.n0 drain_right.t1 9.9005
R66 drain_right.n4 drain_right.t2 9.9005
R67 drain_right.n4 drain_right.t7 9.9005
R68 drain_right.n5 drain_right.t5 9.9005
R69 drain_right.n5 drain_right.t10 9.9005
R70 drain_right.n7 drain_right.t3 9.9005
R71 drain_right.n7 drain_right.t11 9.9005
R72 drain_right drain_right.n8 6.19632
R73 drain_right.n8 drain_right.n6 0.543603
R74 source.n74 source.n72 289.615
R75 source.n62 source.n60 289.615
R76 source.n54 source.n52 289.615
R77 source.n42 source.n40 289.615
R78 source.n2 source.n0 289.615
R79 source.n14 source.n12 289.615
R80 source.n22 source.n20 289.615
R81 source.n34 source.n32 289.615
R82 source.n75 source.n74 185
R83 source.n63 source.n62 185
R84 source.n55 source.n54 185
R85 source.n43 source.n42 185
R86 source.n3 source.n2 185
R87 source.n15 source.n14 185
R88 source.n23 source.n22 185
R89 source.n35 source.n34 185
R90 source.t15 source.n73 167.117
R91 source.t22 source.n61 167.117
R92 source.t4 source.n53 167.117
R93 source.t2 source.n41 167.117
R94 source.t5 source.n1 167.117
R95 source.t0 source.n13 167.117
R96 source.t16 source.n21 167.117
R97 source.t21 source.n33 167.117
R98 source.n9 source.n8 84.1169
R99 source.n11 source.n10 84.1169
R100 source.n29 source.n28 84.1169
R101 source.n31 source.n30 84.1169
R102 source.n71 source.n70 84.1168
R103 source.n69 source.n68 84.1168
R104 source.n51 source.n50 84.1168
R105 source.n49 source.n48 84.1168
R106 source.n74 source.t15 52.3082
R107 source.n62 source.t22 52.3082
R108 source.n54 source.t4 52.3082
R109 source.n42 source.t2 52.3082
R110 source.n2 source.t5 52.3082
R111 source.n14 source.t0 52.3082
R112 source.n22 source.t16 52.3082
R113 source.n34 source.t21 52.3082
R114 source.n79 source.n78 31.4096
R115 source.n67 source.n66 31.4096
R116 source.n59 source.n58 31.4096
R117 source.n47 source.n46 31.4096
R118 source.n7 source.n6 31.4096
R119 source.n19 source.n18 31.4096
R120 source.n27 source.n26 31.4096
R121 source.n39 source.n38 31.4096
R122 source.n47 source.n39 14.2551
R123 source.n70 source.t19 9.9005
R124 source.n70 source.t13 9.9005
R125 source.n68 source.t14 9.9005
R126 source.n68 source.t18 9.9005
R127 source.n50 source.t3 9.9005
R128 source.n50 source.t8 9.9005
R129 source.n48 source.t6 9.9005
R130 source.n48 source.t1 9.9005
R131 source.n8 source.t23 9.9005
R132 source.n8 source.t7 9.9005
R133 source.n10 source.t9 9.9005
R134 source.n10 source.t10 9.9005
R135 source.n28 source.t20 9.9005
R136 source.n28 source.t11 9.9005
R137 source.n30 source.t12 9.9005
R138 source.n30 source.t17 9.9005
R139 source.n75 source.n73 9.71174
R140 source.n63 source.n61 9.71174
R141 source.n55 source.n53 9.71174
R142 source.n43 source.n41 9.71174
R143 source.n3 source.n1 9.71174
R144 source.n15 source.n13 9.71174
R145 source.n23 source.n21 9.71174
R146 source.n35 source.n33 9.71174
R147 source.n78 source.n77 9.45567
R148 source.n66 source.n65 9.45567
R149 source.n58 source.n57 9.45567
R150 source.n46 source.n45 9.45567
R151 source.n6 source.n5 9.45567
R152 source.n18 source.n17 9.45567
R153 source.n26 source.n25 9.45567
R154 source.n38 source.n37 9.45567
R155 source.n77 source.n76 9.3005
R156 source.n65 source.n64 9.3005
R157 source.n57 source.n56 9.3005
R158 source.n45 source.n44 9.3005
R159 source.n5 source.n4 9.3005
R160 source.n17 source.n16 9.3005
R161 source.n25 source.n24 9.3005
R162 source.n37 source.n36 9.3005
R163 source.n80 source.n7 8.72059
R164 source.n78 source.n72 8.14595
R165 source.n66 source.n60 8.14595
R166 source.n58 source.n52 8.14595
R167 source.n46 source.n40 8.14595
R168 source.n6 source.n0 8.14595
R169 source.n18 source.n12 8.14595
R170 source.n26 source.n20 8.14595
R171 source.n38 source.n32 8.14595
R172 source.n76 source.n75 7.3702
R173 source.n64 source.n63 7.3702
R174 source.n56 source.n55 7.3702
R175 source.n44 source.n43 7.3702
R176 source.n4 source.n3 7.3702
R177 source.n16 source.n15 7.3702
R178 source.n24 source.n23 7.3702
R179 source.n36 source.n35 7.3702
R180 source.n76 source.n72 5.81868
R181 source.n64 source.n60 5.81868
R182 source.n56 source.n52 5.81868
R183 source.n44 source.n40 5.81868
R184 source.n4 source.n0 5.81868
R185 source.n16 source.n12 5.81868
R186 source.n24 source.n20 5.81868
R187 source.n36 source.n32 5.81868
R188 source.n80 source.n79 5.53498
R189 source.n77 source.n73 3.44771
R190 source.n65 source.n61 3.44771
R191 source.n57 source.n53 3.44771
R192 source.n45 source.n41 3.44771
R193 source.n5 source.n1 3.44771
R194 source.n17 source.n13 3.44771
R195 source.n25 source.n21 3.44771
R196 source.n37 source.n33 3.44771
R197 source.n39 source.n31 0.543603
R198 source.n31 source.n29 0.543603
R199 source.n29 source.n27 0.543603
R200 source.n19 source.n11 0.543603
R201 source.n11 source.n9 0.543603
R202 source.n9 source.n7 0.543603
R203 source.n49 source.n47 0.543603
R204 source.n51 source.n49 0.543603
R205 source.n59 source.n51 0.543603
R206 source.n69 source.n67 0.543603
R207 source.n71 source.n69 0.543603
R208 source.n79 source.n71 0.543603
R209 source.n27 source.n19 0.470328
R210 source.n67 source.n59 0.470328
R211 source source.n80 0.188
R212 plus.n2 plus.t1 312.57
R213 plus.n13 plus.t7 312.57
R214 plus.n17 plus.t10 312.57
R215 plus.n28 plus.t6 312.57
R216 plus.n3 plus.t4 265.101
R217 plus.n4 plus.t9 265.101
R218 plus.n10 plus.t11 265.101
R219 plus.n12 plus.t3 265.101
R220 plus.n19 plus.t5 265.101
R221 plus.n18 plus.t2 265.101
R222 plus.n25 plus.t0 265.101
R223 plus.n27 plus.t8 265.101
R224 plus.n6 plus.n2 161.489
R225 plus.n21 plus.n17 161.489
R226 plus.n6 plus.n5 161.3
R227 plus.n7 plus.n1 161.3
R228 plus.n9 plus.n8 161.3
R229 plus.n11 plus.n0 161.3
R230 plus.n14 plus.n13 161.3
R231 plus.n21 plus.n20 161.3
R232 plus.n22 plus.n16 161.3
R233 plus.n24 plus.n23 161.3
R234 plus.n26 plus.n15 161.3
R235 plus.n29 plus.n28 161.3
R236 plus.n9 plus.n1 73.0308
R237 plus.n24 plus.n16 73.0308
R238 plus.n5 plus.n4 63.5369
R239 plus.n11 plus.n10 63.5369
R240 plus.n26 plus.n25 63.5369
R241 plus.n20 plus.n18 63.5369
R242 plus.n3 plus.n2 44.549
R243 plus.n13 plus.n12 44.549
R244 plus.n28 plus.n27 44.549
R245 plus.n19 plus.n17 44.549
R246 plus.n5 plus.n3 28.4823
R247 plus.n12 plus.n11 28.4823
R248 plus.n27 plus.n26 28.4823
R249 plus.n20 plus.n19 28.4823
R250 plus plus.n29 25.2793
R251 plus.n4 plus.n1 9.49444
R252 plus.n10 plus.n9 9.49444
R253 plus.n25 plus.n24 9.49444
R254 plus.n18 plus.n16 9.49444
R255 plus plus.n14 8.36792
R256 plus.n7 plus.n6 0.189894
R257 plus.n8 plus.n7 0.189894
R258 plus.n8 plus.n0 0.189894
R259 plus.n14 plus.n0 0.189894
R260 plus.n29 plus.n15 0.189894
R261 plus.n23 plus.n15 0.189894
R262 plus.n23 plus.n22 0.189894
R263 plus.n22 plus.n21 0.189894
R264 drain_left.n6 drain_left.n4 101.338
R265 drain_left.n3 drain_left.n2 101.284
R266 drain_left.n3 drain_left.n0 101.284
R267 drain_left.n8 drain_left.n7 100.796
R268 drain_left.n6 drain_left.n5 100.796
R269 drain_left.n3 drain_left.n1 100.796
R270 drain_left drain_left.n3 22.5068
R271 drain_left.n1 drain_left.t11 9.9005
R272 drain_left.n1 drain_left.t9 9.9005
R273 drain_left.n2 drain_left.t6 9.9005
R274 drain_left.n2 drain_left.t1 9.9005
R275 drain_left.n0 drain_left.t5 9.9005
R276 drain_left.n0 drain_left.t3 9.9005
R277 drain_left.n7 drain_left.t8 9.9005
R278 drain_left.n7 drain_left.t4 9.9005
R279 drain_left.n5 drain_left.t2 9.9005
R280 drain_left.n5 drain_left.t0 9.9005
R281 drain_left.n4 drain_left.t10 9.9005
R282 drain_left.n4 drain_left.t7 9.9005
R283 drain_left drain_left.n8 6.19632
R284 drain_left.n8 drain_left.n6 0.543603
C0 drain_right plus 0.313762f
C1 source minus 1.28014f
C2 source drain_left 5.84919f
C3 minus drain_left 0.176707f
C4 source plus 1.29411f
C5 minus plus 3.29942f
C6 drain_left plus 1.29432f
C7 drain_right source 5.84895f
C8 drain_right minus 1.14089f
C9 drain_right drain_left 0.786036f
C10 drain_right a_n1598_n1288# 3.50777f
C11 drain_left a_n1598_n1288# 3.72367f
C12 source a_n1598_n1288# 2.999241f
C13 minus a_n1598_n1288# 5.398246f
C14 plus a_n1598_n1288# 6.036979f
C15 drain_left.t5 a_n1598_n1288# 0.039465f
C16 drain_left.t3 a_n1598_n1288# 0.039465f
C17 drain_left.n0 a_n1598_n1288# 0.249305f
C18 drain_left.t11 a_n1598_n1288# 0.039465f
C19 drain_left.t9 a_n1598_n1288# 0.039465f
C20 drain_left.n1 a_n1598_n1288# 0.247931f
C21 drain_left.t6 a_n1598_n1288# 0.039465f
C22 drain_left.t1 a_n1598_n1288# 0.039465f
C23 drain_left.n2 a_n1598_n1288# 0.249305f
C24 drain_left.n3 a_n1598_n1288# 1.45738f
C25 drain_left.t10 a_n1598_n1288# 0.039465f
C26 drain_left.t7 a_n1598_n1288# 0.039465f
C27 drain_left.n4 a_n1598_n1288# 0.249478f
C28 drain_left.t2 a_n1598_n1288# 0.039465f
C29 drain_left.t0 a_n1598_n1288# 0.039465f
C30 drain_left.n5 a_n1598_n1288# 0.247932f
C31 drain_left.n6 a_n1598_n1288# 0.565547f
C32 drain_left.t8 a_n1598_n1288# 0.039465f
C33 drain_left.t4 a_n1598_n1288# 0.039465f
C34 drain_left.n7 a_n1598_n1288# 0.247932f
C35 drain_left.n8 a_n1598_n1288# 0.486363f
C36 plus.n0 a_n1598_n1288# 0.030793f
C37 plus.t3 a_n1598_n1288# 0.054366f
C38 plus.t11 a_n1598_n1288# 0.054366f
C39 plus.n1 a_n1598_n1288# 0.011449f
C40 plus.t1 a_n1598_n1288# 0.060493f
C41 plus.n2 a_n1598_n1288# 0.046945f
C42 plus.t4 a_n1598_n1288# 0.054366f
C43 plus.n3 a_n1598_n1288# 0.03797f
C44 plus.t9 a_n1598_n1288# 0.054366f
C45 plus.n4 a_n1598_n1288# 0.03797f
C46 plus.n5 a_n1598_n1288# 0.012683f
C47 plus.n6 a_n1598_n1288# 0.070082f
C48 plus.n7 a_n1598_n1288# 0.030793f
C49 plus.n8 a_n1598_n1288# 0.030793f
C50 plus.n9 a_n1598_n1288# 0.011449f
C51 plus.n10 a_n1598_n1288# 0.03797f
C52 plus.n11 a_n1598_n1288# 0.012683f
C53 plus.n12 a_n1598_n1288# 0.03797f
C54 plus.t7 a_n1598_n1288# 0.060493f
C55 plus.n13 a_n1598_n1288# 0.046899f
C56 plus.n14 a_n1598_n1288# 0.221041f
C57 plus.n15 a_n1598_n1288# 0.030793f
C58 plus.t6 a_n1598_n1288# 0.060493f
C59 plus.t8 a_n1598_n1288# 0.054366f
C60 plus.t0 a_n1598_n1288# 0.054366f
C61 plus.n16 a_n1598_n1288# 0.011449f
C62 plus.t10 a_n1598_n1288# 0.060493f
C63 plus.n17 a_n1598_n1288# 0.046945f
C64 plus.t2 a_n1598_n1288# 0.054366f
C65 plus.n18 a_n1598_n1288# 0.03797f
C66 plus.t5 a_n1598_n1288# 0.054366f
C67 plus.n19 a_n1598_n1288# 0.03797f
C68 plus.n20 a_n1598_n1288# 0.012683f
C69 plus.n21 a_n1598_n1288# 0.070082f
C70 plus.n22 a_n1598_n1288# 0.030793f
C71 plus.n23 a_n1598_n1288# 0.030793f
C72 plus.n24 a_n1598_n1288# 0.011449f
C73 plus.n25 a_n1598_n1288# 0.03797f
C74 plus.n26 a_n1598_n1288# 0.012683f
C75 plus.n27 a_n1598_n1288# 0.03797f
C76 plus.n28 a_n1598_n1288# 0.046899f
C77 plus.n29 a_n1598_n1288# 0.66368f
C78 source.n0 a_n1598_n1288# 0.037033f
C79 source.n1 a_n1598_n1288# 0.081939f
C80 source.t5 a_n1598_n1288# 0.061491f
C81 source.n2 a_n1598_n1288# 0.064129f
C82 source.n3 a_n1598_n1288# 0.020673f
C83 source.n4 a_n1598_n1288# 0.013634f
C84 source.n5 a_n1598_n1288# 0.180613f
C85 source.n6 a_n1598_n1288# 0.040596f
C86 source.n7 a_n1598_n1288# 0.383081f
C87 source.t23 a_n1598_n1288# 0.0401f
C88 source.t7 a_n1598_n1288# 0.0401f
C89 source.n8 a_n1598_n1288# 0.214373f
C90 source.n9 a_n1598_n1288# 0.286061f
C91 source.t9 a_n1598_n1288# 0.0401f
C92 source.t10 a_n1598_n1288# 0.0401f
C93 source.n10 a_n1598_n1288# 0.214373f
C94 source.n11 a_n1598_n1288# 0.286061f
C95 source.n12 a_n1598_n1288# 0.037033f
C96 source.n13 a_n1598_n1288# 0.081939f
C97 source.t0 a_n1598_n1288# 0.061491f
C98 source.n14 a_n1598_n1288# 0.064129f
C99 source.n15 a_n1598_n1288# 0.020673f
C100 source.n16 a_n1598_n1288# 0.013634f
C101 source.n17 a_n1598_n1288# 0.180613f
C102 source.n18 a_n1598_n1288# 0.040596f
C103 source.n19 a_n1598_n1288# 0.1037f
C104 source.n20 a_n1598_n1288# 0.037033f
C105 source.n21 a_n1598_n1288# 0.081939f
C106 source.t16 a_n1598_n1288# 0.061491f
C107 source.n22 a_n1598_n1288# 0.064129f
C108 source.n23 a_n1598_n1288# 0.020673f
C109 source.n24 a_n1598_n1288# 0.013634f
C110 source.n25 a_n1598_n1288# 0.180613f
C111 source.n26 a_n1598_n1288# 0.040596f
C112 source.n27 a_n1598_n1288# 0.1037f
C113 source.t20 a_n1598_n1288# 0.0401f
C114 source.t11 a_n1598_n1288# 0.0401f
C115 source.n28 a_n1598_n1288# 0.214373f
C116 source.n29 a_n1598_n1288# 0.286061f
C117 source.t12 a_n1598_n1288# 0.0401f
C118 source.t17 a_n1598_n1288# 0.0401f
C119 source.n30 a_n1598_n1288# 0.214373f
C120 source.n31 a_n1598_n1288# 0.286061f
C121 source.n32 a_n1598_n1288# 0.037033f
C122 source.n33 a_n1598_n1288# 0.081939f
C123 source.t21 a_n1598_n1288# 0.061491f
C124 source.n34 a_n1598_n1288# 0.064129f
C125 source.n35 a_n1598_n1288# 0.020673f
C126 source.n36 a_n1598_n1288# 0.013634f
C127 source.n37 a_n1598_n1288# 0.180613f
C128 source.n38 a_n1598_n1288# 0.040596f
C129 source.n39 a_n1598_n1288# 0.619628f
C130 source.n40 a_n1598_n1288# 0.037033f
C131 source.n41 a_n1598_n1288# 0.081939f
C132 source.t2 a_n1598_n1288# 0.061491f
C133 source.n42 a_n1598_n1288# 0.064129f
C134 source.n43 a_n1598_n1288# 0.020673f
C135 source.n44 a_n1598_n1288# 0.013634f
C136 source.n45 a_n1598_n1288# 0.180613f
C137 source.n46 a_n1598_n1288# 0.040596f
C138 source.n47 a_n1598_n1288# 0.619628f
C139 source.t6 a_n1598_n1288# 0.0401f
C140 source.t1 a_n1598_n1288# 0.0401f
C141 source.n48 a_n1598_n1288# 0.214372f
C142 source.n49 a_n1598_n1288# 0.286063f
C143 source.t3 a_n1598_n1288# 0.0401f
C144 source.t8 a_n1598_n1288# 0.0401f
C145 source.n50 a_n1598_n1288# 0.214372f
C146 source.n51 a_n1598_n1288# 0.286063f
C147 source.n52 a_n1598_n1288# 0.037033f
C148 source.n53 a_n1598_n1288# 0.081939f
C149 source.t4 a_n1598_n1288# 0.061491f
C150 source.n54 a_n1598_n1288# 0.064129f
C151 source.n55 a_n1598_n1288# 0.020673f
C152 source.n56 a_n1598_n1288# 0.013634f
C153 source.n57 a_n1598_n1288# 0.180613f
C154 source.n58 a_n1598_n1288# 0.040596f
C155 source.n59 a_n1598_n1288# 0.1037f
C156 source.n60 a_n1598_n1288# 0.037033f
C157 source.n61 a_n1598_n1288# 0.081939f
C158 source.t22 a_n1598_n1288# 0.061491f
C159 source.n62 a_n1598_n1288# 0.064129f
C160 source.n63 a_n1598_n1288# 0.020673f
C161 source.n64 a_n1598_n1288# 0.013634f
C162 source.n65 a_n1598_n1288# 0.180613f
C163 source.n66 a_n1598_n1288# 0.040596f
C164 source.n67 a_n1598_n1288# 0.1037f
C165 source.t14 a_n1598_n1288# 0.0401f
C166 source.t18 a_n1598_n1288# 0.0401f
C167 source.n68 a_n1598_n1288# 0.214372f
C168 source.n69 a_n1598_n1288# 0.286063f
C169 source.t19 a_n1598_n1288# 0.0401f
C170 source.t13 a_n1598_n1288# 0.0401f
C171 source.n70 a_n1598_n1288# 0.214372f
C172 source.n71 a_n1598_n1288# 0.286063f
C173 source.n72 a_n1598_n1288# 0.037033f
C174 source.n73 a_n1598_n1288# 0.081939f
C175 source.t15 a_n1598_n1288# 0.061491f
C176 source.n74 a_n1598_n1288# 0.064129f
C177 source.n75 a_n1598_n1288# 0.020673f
C178 source.n76 a_n1598_n1288# 0.013634f
C179 source.n77 a_n1598_n1288# 0.180613f
C180 source.n78 a_n1598_n1288# 0.040596f
C181 source.n79 a_n1598_n1288# 0.246926f
C182 source.n80 a_n1598_n1288# 0.627295f
C183 drain_right.t9 a_n1598_n1288# 0.040141f
C184 drain_right.t1 a_n1598_n1288# 0.040141f
C185 drain_right.n0 a_n1598_n1288# 0.253575f
C186 drain_right.t4 a_n1598_n1288# 0.040141f
C187 drain_right.t0 a_n1598_n1288# 0.040141f
C188 drain_right.n1 a_n1598_n1288# 0.252178f
C189 drain_right.t6 a_n1598_n1288# 0.040141f
C190 drain_right.t8 a_n1598_n1288# 0.040141f
C191 drain_right.n2 a_n1598_n1288# 0.253575f
C192 drain_right.n3 a_n1598_n1288# 1.43246f
C193 drain_right.t2 a_n1598_n1288# 0.040141f
C194 drain_right.t7 a_n1598_n1288# 0.040141f
C195 drain_right.n4 a_n1598_n1288# 0.253752f
C196 drain_right.t5 a_n1598_n1288# 0.040141f
C197 drain_right.t10 a_n1598_n1288# 0.040141f
C198 drain_right.n5 a_n1598_n1288# 0.252179f
C199 drain_right.n6 a_n1598_n1288# 0.575235f
C200 drain_right.t3 a_n1598_n1288# 0.040141f
C201 drain_right.t11 a_n1598_n1288# 0.040141f
C202 drain_right.n7 a_n1598_n1288# 0.252179f
C203 drain_right.n8 a_n1598_n1288# 0.494694f
C204 minus.n0 a_n1598_n1288# 0.030222f
C205 minus.t1 a_n1598_n1288# 0.059373f
C206 minus.t10 a_n1598_n1288# 0.053359f
C207 minus.t5 a_n1598_n1288# 0.053359f
C208 minus.n1 a_n1598_n1288# 0.011237f
C209 minus.t6 a_n1598_n1288# 0.059373f
C210 minus.n2 a_n1598_n1288# 0.046076f
C211 minus.t2 a_n1598_n1288# 0.053359f
C212 minus.n3 a_n1598_n1288# 0.037267f
C213 minus.t11 a_n1598_n1288# 0.053359f
C214 minus.n4 a_n1598_n1288# 0.037267f
C215 minus.n5 a_n1598_n1288# 0.012448f
C216 minus.n6 a_n1598_n1288# 0.068785f
C217 minus.n7 a_n1598_n1288# 0.030222f
C218 minus.n8 a_n1598_n1288# 0.030222f
C219 minus.n9 a_n1598_n1288# 0.011237f
C220 minus.n10 a_n1598_n1288# 0.037267f
C221 minus.n11 a_n1598_n1288# 0.012448f
C222 minus.n12 a_n1598_n1288# 0.037267f
C223 minus.n13 a_n1598_n1288# 0.046031f
C224 minus.n14 a_n1598_n1288# 0.680557f
C225 minus.n15 a_n1598_n1288# 0.030222f
C226 minus.t9 a_n1598_n1288# 0.053359f
C227 minus.t3 a_n1598_n1288# 0.053359f
C228 minus.n16 a_n1598_n1288# 0.011237f
C229 minus.t0 a_n1598_n1288# 0.059373f
C230 minus.n17 a_n1598_n1288# 0.046076f
C231 minus.t8 a_n1598_n1288# 0.053359f
C232 minus.n18 a_n1598_n1288# 0.037267f
C233 minus.t4 a_n1598_n1288# 0.053359f
C234 minus.n19 a_n1598_n1288# 0.037267f
C235 minus.n20 a_n1598_n1288# 0.012448f
C236 minus.n21 a_n1598_n1288# 0.068785f
C237 minus.n22 a_n1598_n1288# 0.030222f
C238 minus.n23 a_n1598_n1288# 0.030222f
C239 minus.n24 a_n1598_n1288# 0.011237f
C240 minus.n25 a_n1598_n1288# 0.037267f
C241 minus.n26 a_n1598_n1288# 0.012448f
C242 minus.n27 a_n1598_n1288# 0.037267f
C243 minus.t7 a_n1598_n1288# 0.059373f
C244 minus.n28 a_n1598_n1288# 0.046031f
C245 minus.n29 a_n1598_n1288# 0.198431f
C246 minus.n30 a_n1598_n1288# 0.840809f
.ends

