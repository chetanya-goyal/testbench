* NGSPICE file created from diffpair111.ext - technology: sky130A

.subckt diffpair111 minus drain_right drain_left source plus
X0 a_n1094_n1292# a_n1094_n1292# a_n1094_n1292# a_n1094_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.3
X1 drain_right.t3 minus.t0 source.t6 a_n1094_n1292# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X2 drain_right.t2 minus.t1 source.t4 a_n1094_n1292# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X3 source.t5 minus.t2 drain_right.t1 a_n1094_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X4 a_n1094_n1292# a_n1094_n1292# a_n1094_n1292# a_n1094_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X5 drain_left.t3 plus.t0 source.t3 a_n1094_n1292# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X6 a_n1094_n1292# a_n1094_n1292# a_n1094_n1292# a_n1094_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X7 source.t7 minus.t3 drain_right.t0 a_n1094_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X8 a_n1094_n1292# a_n1094_n1292# a_n1094_n1292# a_n1094_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X9 source.t0 plus.t1 drain_left.t2 a_n1094_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X10 drain_left.t1 plus.t2 source.t1 a_n1094_n1292# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X11 source.t2 plus.t3 drain_left.t0 a_n1094_n1292# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
R0 minus.n0 minus.t2 311.11
R1 minus.n0 minus.t0 311.11
R2 minus.n1 minus.t1 311.11
R3 minus.n1 minus.t3 311.11
R4 minus.n2 minus.n0 187.012
R5 minus.n2 minus.n1 167.809
R6 minus minus.n2 0.188
R7 source.n58 source.n56 289.615
R8 source.n50 source.n48 289.615
R9 source.n42 source.n40 289.615
R10 source.n34 source.n32 289.615
R11 source.n2 source.n0 289.615
R12 source.n10 source.n8 289.615
R13 source.n18 source.n16 289.615
R14 source.n26 source.n24 289.615
R15 source.n59 source.n58 185
R16 source.n51 source.n50 185
R17 source.n43 source.n42 185
R18 source.n35 source.n34 185
R19 source.n3 source.n2 185
R20 source.n11 source.n10 185
R21 source.n19 source.n18 185
R22 source.n27 source.n26 185
R23 source.t4 source.n57 167.117
R24 source.t7 source.n49 167.117
R25 source.t3 source.n41 167.117
R26 source.t2 source.n33 167.117
R27 source.t1 source.n1 167.117
R28 source.t0 source.n9 167.117
R29 source.t6 source.n17 167.117
R30 source.t5 source.n25 167.117
R31 source.n58 source.t4 52.3082
R32 source.n50 source.t7 52.3082
R33 source.n42 source.t3 52.3082
R34 source.n34 source.t2 52.3082
R35 source.n2 source.t1 52.3082
R36 source.n10 source.t0 52.3082
R37 source.n18 source.t6 52.3082
R38 source.n26 source.t5 52.3082
R39 source.n63 source.n62 31.4096
R40 source.n55 source.n54 31.4096
R41 source.n47 source.n46 31.4096
R42 source.n39 source.n38 31.4096
R43 source.n7 source.n6 31.4096
R44 source.n15 source.n14 31.4096
R45 source.n23 source.n22 31.4096
R46 source.n31 source.n30 31.4096
R47 source.n39 source.n31 14.2702
R48 source.n59 source.n57 9.71174
R49 source.n51 source.n49 9.71174
R50 source.n43 source.n41 9.71174
R51 source.n35 source.n33 9.71174
R52 source.n3 source.n1 9.71174
R53 source.n11 source.n9 9.71174
R54 source.n19 source.n17 9.71174
R55 source.n27 source.n25 9.71174
R56 source.n62 source.n61 9.45567
R57 source.n54 source.n53 9.45567
R58 source.n46 source.n45 9.45567
R59 source.n38 source.n37 9.45567
R60 source.n6 source.n5 9.45567
R61 source.n14 source.n13 9.45567
R62 source.n22 source.n21 9.45567
R63 source.n30 source.n29 9.45567
R64 source.n61 source.n60 9.3005
R65 source.n53 source.n52 9.3005
R66 source.n45 source.n44 9.3005
R67 source.n37 source.n36 9.3005
R68 source.n5 source.n4 9.3005
R69 source.n13 source.n12 9.3005
R70 source.n21 source.n20 9.3005
R71 source.n29 source.n28 9.3005
R72 source.n64 source.n7 8.73574
R73 source.n62 source.n56 8.14595
R74 source.n54 source.n48 8.14595
R75 source.n46 source.n40 8.14595
R76 source.n38 source.n32 8.14595
R77 source.n6 source.n0 8.14595
R78 source.n14 source.n8 8.14595
R79 source.n22 source.n16 8.14595
R80 source.n30 source.n24 8.14595
R81 source.n60 source.n59 7.3702
R82 source.n52 source.n51 7.3702
R83 source.n44 source.n43 7.3702
R84 source.n36 source.n35 7.3702
R85 source.n4 source.n3 7.3702
R86 source.n12 source.n11 7.3702
R87 source.n20 source.n19 7.3702
R88 source.n28 source.n27 7.3702
R89 source.n60 source.n56 5.81868
R90 source.n52 source.n48 5.81868
R91 source.n44 source.n40 5.81868
R92 source.n36 source.n32 5.81868
R93 source.n4 source.n0 5.81868
R94 source.n12 source.n8 5.81868
R95 source.n20 source.n16 5.81868
R96 source.n28 source.n24 5.81868
R97 source.n64 source.n63 5.53498
R98 source.n61 source.n57 3.44771
R99 source.n53 source.n49 3.44771
R100 source.n45 source.n41 3.44771
R101 source.n37 source.n33 3.44771
R102 source.n5 source.n1 3.44771
R103 source.n13 source.n9 3.44771
R104 source.n21 source.n17 3.44771
R105 source.n29 source.n25 3.44771
R106 source.n31 source.n23 0.543603
R107 source.n15 source.n7 0.543603
R108 source.n47 source.n39 0.543603
R109 source.n63 source.n55 0.543603
R110 source.n23 source.n15 0.470328
R111 source.n55 source.n47 0.470328
R112 source source.n64 0.188
R113 drain_right drain_right.n0 121.135
R114 drain_right drain_right.n1 106.992
R115 drain_right.n0 drain_right.t0 9.9005
R116 drain_right.n0 drain_right.t2 9.9005
R117 drain_right.n1 drain_right.t1 9.9005
R118 drain_right.n1 drain_right.t3 9.9005
R119 plus.n0 plus.t1 311.11
R120 plus.n0 plus.t2 311.11
R121 plus.n1 plus.t0 311.11
R122 plus.n1 plus.t3 311.11
R123 plus plus.n1 184.681
R124 plus plus.n0 169.665
R125 drain_left drain_left.n0 121.688
R126 drain_left drain_left.n1 106.992
R127 drain_left.n0 drain_left.t0 9.9005
R128 drain_left.n0 drain_left.t3 9.9005
R129 drain_left.n1 drain_left.t2 9.9005
R130 drain_left.n1 drain_left.t1 9.9005
C0 source plus 0.592995f
C1 minus drain_left 0.177036f
C2 drain_right drain_left 0.477659f
C3 minus source 0.579032f
C4 drain_right source 2.69753f
C5 minus plus 2.66409f
C6 drain_right plus 0.261383f
C7 drain_left source 2.69899f
C8 drain_right minus 0.581551f
C9 drain_left plus 0.68253f
C10 drain_right a_n1094_n1292# 3.58534f
C11 drain_left a_n1094_n1292# 3.70846f
C12 source a_n1094_n1292# 2.796051f
C13 minus a_n1094_n1292# 3.373366f
C14 plus a_n1094_n1292# 5.21293f
C15 drain_left.t0 a_n1094_n1292# 0.035949f
C16 drain_left.t3 a_n1094_n1292# 0.035949f
C17 drain_left.n0 a_n1094_n1292# 0.323735f
C18 drain_left.t2 a_n1094_n1292# 0.035949f
C19 drain_left.t1 a_n1094_n1292# 0.035949f
C20 drain_left.n1 a_n1094_n1292# 0.252029f
C21 plus.t1 a_n1094_n1292# 0.083956f
C22 plus.t2 a_n1094_n1292# 0.083956f
C23 plus.n0 a_n1094_n1292# 0.128637f
C24 plus.t3 a_n1094_n1292# 0.083956f
C25 plus.t0 a_n1094_n1292# 0.083956f
C26 plus.n1 a_n1094_n1292# 0.217966f
C27 drain_right.t0 a_n1094_n1292# 0.037174f
C28 drain_right.t2 a_n1094_n1292# 0.037174f
C29 drain_right.n0 a_n1094_n1292# 0.324737f
C30 drain_right.t1 a_n1094_n1292# 0.037174f
C31 drain_right.t3 a_n1094_n1292# 0.037174f
C32 drain_right.n1 a_n1094_n1292# 0.260618f
C33 source.n0 a_n1094_n1292# 0.028727f
C34 source.n1 a_n1094_n1292# 0.063561f
C35 source.t1 a_n1094_n1292# 0.047699f
C36 source.n2 a_n1094_n1292# 0.049745f
C37 source.n3 a_n1094_n1292# 0.016036f
C38 source.n4 a_n1094_n1292# 0.010576f
C39 source.n5 a_n1094_n1292# 0.140104f
C40 source.n6 a_n1094_n1292# 0.031491f
C41 source.n7 a_n1094_n1292# 0.297935f
C42 source.n8 a_n1094_n1292# 0.028727f
C43 source.n9 a_n1094_n1292# 0.063561f
C44 source.t0 a_n1094_n1292# 0.047699f
C45 source.n10 a_n1094_n1292# 0.049745f
C46 source.n11 a_n1094_n1292# 0.016036f
C47 source.n12 a_n1094_n1292# 0.010576f
C48 source.n13 a_n1094_n1292# 0.140104f
C49 source.n14 a_n1094_n1292# 0.031491f
C50 source.n15 a_n1094_n1292# 0.080441f
C51 source.n16 a_n1094_n1292# 0.028727f
C52 source.n17 a_n1094_n1292# 0.063561f
C53 source.t6 a_n1094_n1292# 0.047699f
C54 source.n18 a_n1094_n1292# 0.049745f
C55 source.n19 a_n1094_n1292# 0.016036f
C56 source.n20 a_n1094_n1292# 0.010576f
C57 source.n21 a_n1094_n1292# 0.140104f
C58 source.n22 a_n1094_n1292# 0.031491f
C59 source.n23 a_n1094_n1292# 0.080441f
C60 source.n24 a_n1094_n1292# 0.028727f
C61 source.n25 a_n1094_n1292# 0.063561f
C62 source.t5 a_n1094_n1292# 0.047699f
C63 source.n26 a_n1094_n1292# 0.049745f
C64 source.n27 a_n1094_n1292# 0.016036f
C65 source.n28 a_n1094_n1292# 0.010576f
C66 source.n29 a_n1094_n1292# 0.140104f
C67 source.n30 a_n1094_n1292# 0.031491f
C68 source.n31 a_n1094_n1292# 0.481897f
C69 source.n32 a_n1094_n1292# 0.028727f
C70 source.n33 a_n1094_n1292# 0.063561f
C71 source.t2 a_n1094_n1292# 0.047699f
C72 source.n34 a_n1094_n1292# 0.049745f
C73 source.n35 a_n1094_n1292# 0.016036f
C74 source.n36 a_n1094_n1292# 0.010576f
C75 source.n37 a_n1094_n1292# 0.140104f
C76 source.n38 a_n1094_n1292# 0.031491f
C77 source.n39 a_n1094_n1292# 0.481897f
C78 source.n40 a_n1094_n1292# 0.028727f
C79 source.n41 a_n1094_n1292# 0.063561f
C80 source.t3 a_n1094_n1292# 0.047699f
C81 source.n42 a_n1094_n1292# 0.049745f
C82 source.n43 a_n1094_n1292# 0.016036f
C83 source.n44 a_n1094_n1292# 0.010576f
C84 source.n45 a_n1094_n1292# 0.140104f
C85 source.n46 a_n1094_n1292# 0.031491f
C86 source.n47 a_n1094_n1292# 0.080441f
C87 source.n48 a_n1094_n1292# 0.028727f
C88 source.n49 a_n1094_n1292# 0.063561f
C89 source.t7 a_n1094_n1292# 0.047699f
C90 source.n50 a_n1094_n1292# 0.049745f
C91 source.n51 a_n1094_n1292# 0.016036f
C92 source.n52 a_n1094_n1292# 0.010576f
C93 source.n53 a_n1094_n1292# 0.140104f
C94 source.n54 a_n1094_n1292# 0.031491f
C95 source.n55 a_n1094_n1292# 0.080441f
C96 source.n56 a_n1094_n1292# 0.028727f
C97 source.n57 a_n1094_n1292# 0.063561f
C98 source.t4 a_n1094_n1292# 0.047699f
C99 source.n58 a_n1094_n1292# 0.049745f
C100 source.n59 a_n1094_n1292# 0.016036f
C101 source.n60 a_n1094_n1292# 0.010576f
C102 source.n61 a_n1094_n1292# 0.140104f
C103 source.n62 a_n1094_n1292# 0.031491f
C104 source.n63 a_n1094_n1292# 0.191544f
C105 source.n64 a_n1094_n1292# 0.488315f
C106 minus.t2 a_n1094_n1292# 0.081345f
C107 minus.t0 a_n1094_n1292# 0.081345f
C108 minus.n0 a_n1094_n1292# 0.223839f
C109 minus.t3 a_n1094_n1292# 0.081345f
C110 minus.t1 a_n1094_n1292# 0.081345f
C111 minus.n1 a_n1094_n1292# 0.120402f
C112 minus.n2 a_n1094_n1292# 2.0031f
.ends

