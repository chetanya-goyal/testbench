* NGSPICE file created from diffpair530.ext - technology: sky130A

.subckt diffpair530 minus drain_right drain_left source plus
X0 drain_right minus source a_n1088_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=5.85 ps=30.78 w=15 l=0.6
X1 drain_left plus source a_n1088_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=5.85 ps=30.78 w=15 l=0.6
X2 drain_right minus source a_n1088_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=5.85 ps=30.78 w=15 l=0.6
X3 drain_left plus source a_n1088_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=5.85 ps=30.78 w=15 l=0.6
X4 a_n1088_n3892# a_n1088_n3892# a_n1088_n3892# a_n1088_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.6
X5 a_n1088_n3892# a_n1088_n3892# a_n1088_n3892# a_n1088_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.6
X6 a_n1088_n3892# a_n1088_n3892# a_n1088_n3892# a_n1088_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.6
X7 a_n1088_n3892# a_n1088_n3892# a_n1088_n3892# a_n1088_n3892# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.6
.ends

