* NGSPICE file created from diffpair29.ext - technology: sky130A

.subckt diffpair29 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t47 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X1 drain_left.t22 plus.t1 source.t45 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X2 source.t5 minus.t0 drain_right.t23 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X3 drain_left.t21 plus.t2 source.t42 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X4 drain_left.t20 plus.t3 source.t34 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X5 source.t16 minus.t1 drain_right.t22 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X6 drain_left.t19 plus.t4 source.t24 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X7 source.t20 minus.t2 drain_right.t21 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X8 drain_right.t20 minus.t3 source.t18 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X9 source.t4 minus.t4 drain_right.t19 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X10 source.t15 minus.t5 drain_right.t18 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X11 source.t19 minus.t6 drain_right.t17 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X12 source.t26 plus.t5 drain_left.t18 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X13 drain_right.t16 minus.t7 source.t17 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X14 source.t14 minus.t8 drain_right.t15 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X15 source.t13 minus.t9 drain_right.t14 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X16 a_n2224_n1088# a_n2224_n1088# a_n2224_n1088# a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.25
X17 source.t12 minus.t10 drain_right.t13 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X18 drain_right.t12 minus.t11 source.t11 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X19 drain_right.t11 minus.t12 source.t21 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X20 a_n2224_n1088# a_n2224_n1088# a_n2224_n1088# a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X21 source.t23 minus.t13 drain_right.t10 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X22 drain_right.t9 minus.t14 source.t22 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X23 source.t29 plus.t6 drain_left.t17 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X24 source.t30 plus.t7 drain_left.t16 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X25 source.t40 plus.t8 drain_left.t15 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X26 source.t32 plus.t9 drain_left.t14 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X27 drain_left.t13 plus.t10 source.t37 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X28 source.t10 minus.t15 drain_right.t8 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X29 drain_left.t12 plus.t11 source.t41 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X30 source.t28 plus.t12 drain_left.t11 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X31 drain_right.t7 minus.t16 source.t9 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X32 drain_left.t10 plus.t13 source.t33 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X33 source.t25 plus.t14 drain_left.t9 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X34 drain_right.t6 minus.t17 source.t3 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.25
X35 drain_left.t8 plus.t15 source.t27 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X36 source.t8 minus.t18 drain_right.t5 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X37 a_n2224_n1088# a_n2224_n1088# a_n2224_n1088# a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X38 source.t39 plus.t16 drain_left.t7 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X39 source.t46 plus.t17 drain_left.t6 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.25
X40 source.t44 plus.t18 drain_left.t5 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X41 drain_left.t4 plus.t19 source.t38 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X42 a_n2224_n1088# a_n2224_n1088# a_n2224_n1088# a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.25
X43 source.t43 plus.t20 drain_left.t3 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X44 drain_right.t4 minus.t19 source.t1 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X45 drain_right.t3 minus.t20 source.t2 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X46 source.t36 plus.t21 drain_left.t2 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X47 drain_right.t2 minus.t21 source.t6 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X48 drain_right.t1 minus.t22 source.t7 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X49 drain_left.t1 plus.t22 source.t35 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X50 drain_left.t0 plus.t23 source.t31 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
X51 drain_right.t0 minus.t23 source.t0 a_n2224_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.25
R0 plus.n6 plus.t5 249.472
R1 plus.n33 plus.t2 249.472
R2 plus.n42 plus.t11 249.472
R3 plus.n68 plus.t17 249.472
R4 plus.n7 plus.t1 221.72
R5 plus.n8 plus.t9 221.72
R6 plus.n14 plus.t0 221.72
R7 plus.n16 plus.t8 221.72
R8 plus.n3 plus.t22 221.72
R9 plus.n21 plus.t7 221.72
R10 plus.n23 plus.t4 221.72
R11 plus.n24 plus.t14 221.72
R12 plus.n30 plus.t3 221.72
R13 plus.n32 plus.t12 221.72
R14 plus.n44 plus.t6 221.72
R15 plus.n43 plus.t15 221.72
R16 plus.n50 plus.t20 221.72
R17 plus.n52 plus.t10 221.72
R18 plus.n39 plus.t16 221.72
R19 plus.n57 plus.t13 221.72
R20 plus.n59 plus.t18 221.72
R21 plus.n38 plus.t23 221.72
R22 plus.n65 plus.t21 221.72
R23 plus.n67 plus.t19 221.72
R24 plus.n10 plus.n6 161.489
R25 plus.n46 plus.n42 161.489
R26 plus.n10 plus.n9 161.3
R27 plus.n11 plus.n5 161.3
R28 plus.n13 plus.n12 161.3
R29 plus.n15 plus.n4 161.3
R30 plus.n18 plus.n17 161.3
R31 plus.n20 plus.n19 161.3
R32 plus.n22 plus.n2 161.3
R33 plus.n26 plus.n25 161.3
R34 plus.n27 plus.n1 161.3
R35 plus.n29 plus.n28 161.3
R36 plus.n31 plus.n0 161.3
R37 plus.n34 plus.n33 161.3
R38 plus.n46 plus.n45 161.3
R39 plus.n47 plus.n41 161.3
R40 plus.n49 plus.n48 161.3
R41 plus.n51 plus.n40 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n56 plus.n55 161.3
R44 plus.n58 plus.n37 161.3
R45 plus.n61 plus.n60 161.3
R46 plus.n62 plus.n36 161.3
R47 plus.n64 plus.n63 161.3
R48 plus.n66 plus.n35 161.3
R49 plus.n69 plus.n68 161.3
R50 plus.n13 plus.n5 73.0308
R51 plus.n29 plus.n1 73.0308
R52 plus.n64 plus.n36 73.0308
R53 plus.n49 plus.n41 73.0308
R54 plus.n9 plus.n8 68.649
R55 plus.n31 plus.n30 68.649
R56 plus.n66 plus.n65 68.649
R57 plus.n45 plus.n43 68.649
R58 plus.n15 plus.n14 65.7278
R59 plus.n25 plus.n24 65.7278
R60 plus.n60 plus.n38 65.7278
R61 plus.n51 plus.n50 65.7278
R62 plus.n7 plus.n6 56.9641
R63 plus.n33 plus.n32 56.9641
R64 plus.n68 plus.n67 56.9641
R65 plus.n44 plus.n42 56.9641
R66 plus.n17 plus.n16 54.0429
R67 plus.n23 plus.n22 54.0429
R68 plus.n59 plus.n58 54.0429
R69 plus.n53 plus.n52 54.0429
R70 plus.n20 plus.n3 42.3581
R71 plus.n21 plus.n20 42.3581
R72 plus.n57 plus.n56 42.3581
R73 plus.n56 plus.n39 42.3581
R74 plus.n17 plus.n3 30.6732
R75 plus.n22 plus.n21 30.6732
R76 plus.n58 plus.n57 30.6732
R77 plus.n53 plus.n39 30.6732
R78 plus plus.n69 27.1922
R79 plus.n16 plus.n15 18.9884
R80 plus.n25 plus.n23 18.9884
R81 plus.n60 plus.n59 18.9884
R82 plus.n52 plus.n51 18.9884
R83 plus.n9 plus.n7 16.0672
R84 plus.n32 plus.n31 16.0672
R85 plus.n67 plus.n66 16.0672
R86 plus.n45 plus.n44 16.0672
R87 plus plus.n34 7.90959
R88 plus.n14 plus.n13 7.30353
R89 plus.n24 plus.n1 7.30353
R90 plus.n38 plus.n36 7.30353
R91 plus.n50 plus.n49 7.30353
R92 plus.n8 plus.n5 4.38232
R93 plus.n30 plus.n29 4.38232
R94 plus.n65 plus.n64 4.38232
R95 plus.n43 plus.n41 4.38232
R96 plus.n11 plus.n10 0.189894
R97 plus.n12 plus.n11 0.189894
R98 plus.n12 plus.n4 0.189894
R99 plus.n18 plus.n4 0.189894
R100 plus.n19 plus.n18 0.189894
R101 plus.n19 plus.n2 0.189894
R102 plus.n26 plus.n2 0.189894
R103 plus.n27 plus.n26 0.189894
R104 plus.n28 plus.n27 0.189894
R105 plus.n28 plus.n0 0.189894
R106 plus.n34 plus.n0 0.189894
R107 plus.n69 plus.n35 0.189894
R108 plus.n63 plus.n35 0.189894
R109 plus.n63 plus.n62 0.189894
R110 plus.n62 plus.n61 0.189894
R111 plus.n61 plus.n37 0.189894
R112 plus.n55 plus.n37 0.189894
R113 plus.n55 plus.n54 0.189894
R114 plus.n54 plus.n40 0.189894
R115 plus.n48 plus.n40 0.189894
R116 plus.n48 plus.n47 0.189894
R117 plus.n47 plus.n46 0.189894
R118 source.n0 source.t42 243.255
R119 source.n11 source.t26 243.255
R120 source.n12 source.t3 243.255
R121 source.n23 source.t8 243.255
R122 source.n47 source.t22 243.254
R123 source.n36 source.t19 243.254
R124 source.n35 source.t41 243.254
R125 source.n24 source.t46 243.254
R126 source.n2 source.n1 223.454
R127 source.n4 source.n3 223.454
R128 source.n6 source.n5 223.454
R129 source.n8 source.n7 223.454
R130 source.n10 source.n9 223.454
R131 source.n14 source.n13 223.454
R132 source.n16 source.n15 223.454
R133 source.n18 source.n17 223.454
R134 source.n20 source.n19 223.454
R135 source.n22 source.n21 223.454
R136 source.n46 source.n45 223.453
R137 source.n44 source.n43 223.453
R138 source.n42 source.n41 223.453
R139 source.n40 source.n39 223.453
R140 source.n38 source.n37 223.453
R141 source.n34 source.n33 223.453
R142 source.n32 source.n31 223.453
R143 source.n30 source.n29 223.453
R144 source.n28 source.n27 223.453
R145 source.n26 source.n25 223.453
R146 source.n45 source.t11 19.8005
R147 source.n45 source.t10 19.8005
R148 source.n43 source.t17 19.8005
R149 source.n43 source.t4 19.8005
R150 source.n41 source.t21 19.8005
R151 source.n41 source.t14 19.8005
R152 source.n39 source.t0 19.8005
R153 source.n39 source.t15 19.8005
R154 source.n37 source.t7 19.8005
R155 source.n37 source.t5 19.8005
R156 source.n33 source.t27 19.8005
R157 source.n33 source.t29 19.8005
R158 source.n31 source.t37 19.8005
R159 source.n31 source.t43 19.8005
R160 source.n29 source.t33 19.8005
R161 source.n29 source.t39 19.8005
R162 source.n27 source.t31 19.8005
R163 source.n27 source.t44 19.8005
R164 source.n25 source.t38 19.8005
R165 source.n25 source.t36 19.8005
R166 source.n1 source.t34 19.8005
R167 source.n1 source.t28 19.8005
R168 source.n3 source.t24 19.8005
R169 source.n3 source.t25 19.8005
R170 source.n5 source.t35 19.8005
R171 source.n5 source.t30 19.8005
R172 source.n7 source.t47 19.8005
R173 source.n7 source.t40 19.8005
R174 source.n9 source.t45 19.8005
R175 source.n9 source.t32 19.8005
R176 source.n13 source.t9 19.8005
R177 source.n13 source.t20 19.8005
R178 source.n15 source.t1 19.8005
R179 source.n15 source.t16 19.8005
R180 source.n17 source.t2 19.8005
R181 source.n17 source.t12 19.8005
R182 source.n19 source.t6 19.8005
R183 source.n19 source.t13 19.8005
R184 source.n21 source.t18 19.8005
R185 source.n21 source.t23 19.8005
R186 source.n24 source.n23 13.4544
R187 source.n48 source.n0 7.94146
R188 source.n48 source.n47 5.51343
R189 source.n23 source.n22 0.5005
R190 source.n22 source.n20 0.5005
R191 source.n20 source.n18 0.5005
R192 source.n18 source.n16 0.5005
R193 source.n16 source.n14 0.5005
R194 source.n14 source.n12 0.5005
R195 source.n11 source.n10 0.5005
R196 source.n10 source.n8 0.5005
R197 source.n8 source.n6 0.5005
R198 source.n6 source.n4 0.5005
R199 source.n4 source.n2 0.5005
R200 source.n2 source.n0 0.5005
R201 source.n26 source.n24 0.5005
R202 source.n28 source.n26 0.5005
R203 source.n30 source.n28 0.5005
R204 source.n32 source.n30 0.5005
R205 source.n34 source.n32 0.5005
R206 source.n35 source.n34 0.5005
R207 source.n38 source.n36 0.5005
R208 source.n40 source.n38 0.5005
R209 source.n42 source.n40 0.5005
R210 source.n44 source.n42 0.5005
R211 source.n46 source.n44 0.5005
R212 source.n47 source.n46 0.5005
R213 source.n12 source.n11 0.470328
R214 source.n36 source.n35 0.470328
R215 source source.n48 0.188
R216 drain_left.n13 drain_left.n11 240.632
R217 drain_left.n7 drain_left.n5 240.631
R218 drain_left.n2 drain_left.n0 240.631
R219 drain_left.n21 drain_left.n20 240.132
R220 drain_left.n19 drain_left.n18 240.132
R221 drain_left.n17 drain_left.n16 240.132
R222 drain_left.n15 drain_left.n14 240.132
R223 drain_left.n13 drain_left.n12 240.132
R224 drain_left.n7 drain_left.n6 240.131
R225 drain_left.n9 drain_left.n8 240.131
R226 drain_left.n4 drain_left.n3 240.131
R227 drain_left.n2 drain_left.n1 240.131
R228 drain_left drain_left.n10 23.7837
R229 drain_left.n5 drain_left.t17 19.8005
R230 drain_left.n5 drain_left.t12 19.8005
R231 drain_left.n6 drain_left.t3 19.8005
R232 drain_left.n6 drain_left.t8 19.8005
R233 drain_left.n8 drain_left.t7 19.8005
R234 drain_left.n8 drain_left.t13 19.8005
R235 drain_left.n3 drain_left.t5 19.8005
R236 drain_left.n3 drain_left.t10 19.8005
R237 drain_left.n1 drain_left.t2 19.8005
R238 drain_left.n1 drain_left.t0 19.8005
R239 drain_left.n0 drain_left.t6 19.8005
R240 drain_left.n0 drain_left.t4 19.8005
R241 drain_left.n20 drain_left.t11 19.8005
R242 drain_left.n20 drain_left.t21 19.8005
R243 drain_left.n18 drain_left.t9 19.8005
R244 drain_left.n18 drain_left.t20 19.8005
R245 drain_left.n16 drain_left.t16 19.8005
R246 drain_left.n16 drain_left.t19 19.8005
R247 drain_left.n14 drain_left.t15 19.8005
R248 drain_left.n14 drain_left.t1 19.8005
R249 drain_left.n12 drain_left.t14 19.8005
R250 drain_left.n12 drain_left.t23 19.8005
R251 drain_left.n11 drain_left.t18 19.8005
R252 drain_left.n11 drain_left.t22 19.8005
R253 drain_left drain_left.n21 6.15322
R254 drain_left.n9 drain_left.n7 0.5005
R255 drain_left.n4 drain_left.n2 0.5005
R256 drain_left.n15 drain_left.n13 0.5005
R257 drain_left.n17 drain_left.n15 0.5005
R258 drain_left.n19 drain_left.n17 0.5005
R259 drain_left.n21 drain_left.n19 0.5005
R260 drain_left.n10 drain_left.n9 0.195154
R261 drain_left.n10 drain_left.n4 0.195154
R262 minus.n33 minus.t18 249.472
R263 minus.n7 minus.t17 249.472
R264 minus.n68 minus.t14 249.472
R265 minus.n41 minus.t6 249.472
R266 minus.n32 minus.t3 221.72
R267 minus.n30 minus.t13 221.72
R268 minus.n3 minus.t21 221.72
R269 minus.n24 minus.t9 221.72
R270 minus.n22 minus.t20 221.72
R271 minus.n4 minus.t10 221.72
R272 minus.n17 minus.t19 221.72
R273 minus.n15 minus.t1 221.72
R274 minus.n8 minus.t16 221.72
R275 minus.n9 minus.t2 221.72
R276 minus.n67 minus.t15 221.72
R277 minus.n65 minus.t11 221.72
R278 minus.n59 minus.t4 221.72
R279 minus.n58 minus.t7 221.72
R280 minus.n56 minus.t8 221.72
R281 minus.n38 minus.t12 221.72
R282 minus.n51 minus.t5 221.72
R283 minus.n49 minus.t23 221.72
R284 minus.n43 minus.t0 221.72
R285 minus.n42 minus.t22 221.72
R286 minus.n11 minus.n7 161.489
R287 minus.n45 minus.n41 161.489
R288 minus.n34 minus.n33 161.3
R289 minus.n31 minus.n0 161.3
R290 minus.n29 minus.n28 161.3
R291 minus.n27 minus.n1 161.3
R292 minus.n26 minus.n25 161.3
R293 minus.n23 minus.n2 161.3
R294 minus.n21 minus.n20 161.3
R295 minus.n19 minus.n18 161.3
R296 minus.n16 minus.n5 161.3
R297 minus.n14 minus.n13 161.3
R298 minus.n12 minus.n6 161.3
R299 minus.n11 minus.n10 161.3
R300 minus.n69 minus.n68 161.3
R301 minus.n66 minus.n35 161.3
R302 minus.n64 minus.n63 161.3
R303 minus.n62 minus.n36 161.3
R304 minus.n61 minus.n60 161.3
R305 minus.n57 minus.n37 161.3
R306 minus.n55 minus.n54 161.3
R307 minus.n53 minus.n52 161.3
R308 minus.n50 minus.n39 161.3
R309 minus.n48 minus.n47 161.3
R310 minus.n46 minus.n40 161.3
R311 minus.n45 minus.n44 161.3
R312 minus.n29 minus.n1 73.0308
R313 minus.n14 minus.n6 73.0308
R314 minus.n48 minus.n40 73.0308
R315 minus.n64 minus.n36 73.0308
R316 minus.n31 minus.n30 68.649
R317 minus.n10 minus.n8 68.649
R318 minus.n44 minus.n43 68.649
R319 minus.n66 minus.n65 68.649
R320 minus.n25 minus.n3 65.7278
R321 minus.n16 minus.n15 65.7278
R322 minus.n50 minus.n49 65.7278
R323 minus.n60 minus.n59 65.7278
R324 minus.n33 minus.n32 56.9641
R325 minus.n9 minus.n7 56.9641
R326 minus.n42 minus.n41 56.9641
R327 minus.n68 minus.n67 56.9641
R328 minus.n24 minus.n23 54.0429
R329 minus.n18 minus.n17 54.0429
R330 minus.n52 minus.n51 54.0429
R331 minus.n58 minus.n57 54.0429
R332 minus.n22 minus.n21 42.3581
R333 minus.n21 minus.n4 42.3581
R334 minus.n55 minus.n38 42.3581
R335 minus.n56 minus.n55 42.3581
R336 minus.n23 minus.n22 30.6732
R337 minus.n18 minus.n4 30.6732
R338 minus.n52 minus.n38 30.6732
R339 minus.n57 minus.n56 30.6732
R340 minus.n70 minus.n34 29.1444
R341 minus.n25 minus.n24 18.9884
R342 minus.n17 minus.n16 18.9884
R343 minus.n51 minus.n50 18.9884
R344 minus.n60 minus.n58 18.9884
R345 minus.n32 minus.n31 16.0672
R346 minus.n10 minus.n9 16.0672
R347 minus.n44 minus.n42 16.0672
R348 minus.n67 minus.n66 16.0672
R349 minus.n3 minus.n1 7.30353
R350 minus.n15 minus.n14 7.30353
R351 minus.n49 minus.n48 7.30353
R352 minus.n59 minus.n36 7.30353
R353 minus.n70 minus.n69 6.43232
R354 minus.n30 minus.n29 4.38232
R355 minus.n8 minus.n6 4.38232
R356 minus.n43 minus.n40 4.38232
R357 minus.n65 minus.n64 4.38232
R358 minus.n34 minus.n0 0.189894
R359 minus.n28 minus.n0 0.189894
R360 minus.n28 minus.n27 0.189894
R361 minus.n27 minus.n26 0.189894
R362 minus.n26 minus.n2 0.189894
R363 minus.n20 minus.n2 0.189894
R364 minus.n20 minus.n19 0.189894
R365 minus.n19 minus.n5 0.189894
R366 minus.n13 minus.n5 0.189894
R367 minus.n13 minus.n12 0.189894
R368 minus.n12 minus.n11 0.189894
R369 minus.n46 minus.n45 0.189894
R370 minus.n47 minus.n46 0.189894
R371 minus.n47 minus.n39 0.189894
R372 minus.n53 minus.n39 0.189894
R373 minus.n54 minus.n53 0.189894
R374 minus.n54 minus.n37 0.189894
R375 minus.n61 minus.n37 0.189894
R376 minus.n62 minus.n61 0.189894
R377 minus.n63 minus.n62 0.189894
R378 minus.n63 minus.n35 0.189894
R379 minus.n69 minus.n35 0.189894
R380 minus minus.n70 0.188
R381 drain_right.n13 drain_right.n11 240.632
R382 drain_right.n7 drain_right.n5 240.631
R383 drain_right.n2 drain_right.n0 240.631
R384 drain_right.n13 drain_right.n12 240.132
R385 drain_right.n15 drain_right.n14 240.132
R386 drain_right.n17 drain_right.n16 240.132
R387 drain_right.n19 drain_right.n18 240.132
R388 drain_right.n21 drain_right.n20 240.132
R389 drain_right.n7 drain_right.n6 240.131
R390 drain_right.n9 drain_right.n8 240.131
R391 drain_right.n4 drain_right.n3 240.131
R392 drain_right.n2 drain_right.n1 240.131
R393 drain_right drain_right.n10 23.2305
R394 drain_right.n5 drain_right.t8 19.8005
R395 drain_right.n5 drain_right.t9 19.8005
R396 drain_right.n6 drain_right.t19 19.8005
R397 drain_right.n6 drain_right.t12 19.8005
R398 drain_right.n8 drain_right.t15 19.8005
R399 drain_right.n8 drain_right.t16 19.8005
R400 drain_right.n3 drain_right.t18 19.8005
R401 drain_right.n3 drain_right.t11 19.8005
R402 drain_right.n1 drain_right.t23 19.8005
R403 drain_right.n1 drain_right.t0 19.8005
R404 drain_right.n0 drain_right.t17 19.8005
R405 drain_right.n0 drain_right.t1 19.8005
R406 drain_right.n11 drain_right.t21 19.8005
R407 drain_right.n11 drain_right.t6 19.8005
R408 drain_right.n12 drain_right.t22 19.8005
R409 drain_right.n12 drain_right.t7 19.8005
R410 drain_right.n14 drain_right.t13 19.8005
R411 drain_right.n14 drain_right.t4 19.8005
R412 drain_right.n16 drain_right.t14 19.8005
R413 drain_right.n16 drain_right.t3 19.8005
R414 drain_right.n18 drain_right.t10 19.8005
R415 drain_right.n18 drain_right.t2 19.8005
R416 drain_right.n20 drain_right.t5 19.8005
R417 drain_right.n20 drain_right.t20 19.8005
R418 drain_right drain_right.n21 6.15322
R419 drain_right.n9 drain_right.n7 0.5005
R420 drain_right.n4 drain_right.n2 0.5005
R421 drain_right.n21 drain_right.n19 0.5005
R422 drain_right.n19 drain_right.n17 0.5005
R423 drain_right.n17 drain_right.n15 0.5005
R424 drain_right.n15 drain_right.n13 0.5005
R425 drain_right.n10 drain_right.n9 0.195154
R426 drain_right.n10 drain_right.n4 0.195154
C0 drain_right plus 0.382759f
C1 drain_right source 7.459009f
C2 drain_left plus 1.43512f
C3 drain_left source 7.45859f
C4 drain_right minus 1.21656f
C5 source plus 1.59819f
C6 drain_left minus 0.179776f
C7 minus plus 3.90714f
C8 drain_right drain_left 1.19776f
C9 source minus 1.58432f
C10 drain_right a_n2224_n1088# 4.3878f
C11 drain_left a_n2224_n1088# 4.68942f
C12 source a_n2224_n1088# 2.738475f
C13 minus a_n2224_n1088# 7.823098f
C14 plus a_n2224_n1088# 8.493916f
C15 drain_right.t17 a_n2224_n1088# 0.022119f
C16 drain_right.t1 a_n2224_n1088# 0.022119f
C17 drain_right.n0 a_n2224_n1088# 0.086566f
C18 drain_right.t23 a_n2224_n1088# 0.022119f
C19 drain_right.t0 a_n2224_n1088# 0.022119f
C20 drain_right.n1 a_n2224_n1088# 0.085948f
C21 drain_right.n2 a_n2224_n1088# 0.582524f
C22 drain_right.t18 a_n2224_n1088# 0.022119f
C23 drain_right.t11 a_n2224_n1088# 0.022119f
C24 drain_right.n3 a_n2224_n1088# 0.085948f
C25 drain_right.n4 a_n2224_n1088# 0.261728f
C26 drain_right.t8 a_n2224_n1088# 0.022119f
C27 drain_right.t9 a_n2224_n1088# 0.022119f
C28 drain_right.n5 a_n2224_n1088# 0.086566f
C29 drain_right.t19 a_n2224_n1088# 0.022119f
C30 drain_right.t12 a_n2224_n1088# 0.022119f
C31 drain_right.n6 a_n2224_n1088# 0.085948f
C32 drain_right.n7 a_n2224_n1088# 0.582524f
C33 drain_right.t15 a_n2224_n1088# 0.022119f
C34 drain_right.t16 a_n2224_n1088# 0.022119f
C35 drain_right.n8 a_n2224_n1088# 0.085948f
C36 drain_right.n9 a_n2224_n1088# 0.261728f
C37 drain_right.n10 a_n2224_n1088# 0.798316f
C38 drain_right.t21 a_n2224_n1088# 0.022119f
C39 drain_right.t6 a_n2224_n1088# 0.022119f
C40 drain_right.n11 a_n2224_n1088# 0.086566f
C41 drain_right.t22 a_n2224_n1088# 0.022119f
C42 drain_right.t7 a_n2224_n1088# 0.022119f
C43 drain_right.n12 a_n2224_n1088# 0.085948f
C44 drain_right.n13 a_n2224_n1088# 0.582524f
C45 drain_right.t13 a_n2224_n1088# 0.022119f
C46 drain_right.t4 a_n2224_n1088# 0.022119f
C47 drain_right.n14 a_n2224_n1088# 0.085948f
C48 drain_right.n15 a_n2224_n1088# 0.285934f
C49 drain_right.t14 a_n2224_n1088# 0.022119f
C50 drain_right.t3 a_n2224_n1088# 0.022119f
C51 drain_right.n16 a_n2224_n1088# 0.085948f
C52 drain_right.n17 a_n2224_n1088# 0.285934f
C53 drain_right.t10 a_n2224_n1088# 0.022119f
C54 drain_right.t2 a_n2224_n1088# 0.022119f
C55 drain_right.n18 a_n2224_n1088# 0.085948f
C56 drain_right.n19 a_n2224_n1088# 0.285934f
C57 drain_right.t5 a_n2224_n1088# 0.022119f
C58 drain_right.t20 a_n2224_n1088# 0.022119f
C59 drain_right.n20 a_n2224_n1088# 0.085948f
C60 drain_right.n21 a_n2224_n1088# 0.516978f
C61 minus.n0 a_n2224_n1088# 0.028931f
C62 minus.t18 a_n2224_n1088# 0.024898f
C63 minus.t3 a_n2224_n1088# 0.022296f
C64 minus.t13 a_n2224_n1088# 0.022296f
C65 minus.n1 a_n2224_n1088# 0.010489f
C66 minus.n2 a_n2224_n1088# 0.028931f
C67 minus.t21 a_n2224_n1088# 0.022296f
C68 minus.n3 a_n2224_n1088# 0.024458f
C69 minus.t9 a_n2224_n1088# 0.022296f
C70 minus.t20 a_n2224_n1088# 0.022296f
C71 minus.t10 a_n2224_n1088# 0.022296f
C72 minus.n4 a_n2224_n1088# 0.024458f
C73 minus.n5 a_n2224_n1088# 0.028931f
C74 minus.t19 a_n2224_n1088# 0.022296f
C75 minus.t1 a_n2224_n1088# 0.022296f
C76 minus.n6 a_n2224_n1088# 0.010132f
C77 minus.t17 a_n2224_n1088# 0.024898f
C78 minus.n7 a_n2224_n1088# 0.031847f
C79 minus.t16 a_n2224_n1088# 0.022296f
C80 minus.n8 a_n2224_n1088# 0.024458f
C81 minus.t2 a_n2224_n1088# 0.022296f
C82 minus.n9 a_n2224_n1088# 0.024458f
C83 minus.n10 a_n2224_n1088# 0.011024f
C84 minus.n11 a_n2224_n1088# 0.060144f
C85 minus.n12 a_n2224_n1088# 0.028931f
C86 minus.n13 a_n2224_n1088# 0.028931f
C87 minus.n14 a_n2224_n1088# 0.010489f
C88 minus.n15 a_n2224_n1088# 0.024458f
C89 minus.n16 a_n2224_n1088# 0.011024f
C90 minus.n17 a_n2224_n1088# 0.024458f
C91 minus.n18 a_n2224_n1088# 0.011024f
C92 minus.n19 a_n2224_n1088# 0.028931f
C93 minus.n20 a_n2224_n1088# 0.028931f
C94 minus.n21 a_n2224_n1088# 0.011024f
C95 minus.n22 a_n2224_n1088# 0.024458f
C96 minus.n23 a_n2224_n1088# 0.011024f
C97 minus.n24 a_n2224_n1088# 0.024458f
C98 minus.n25 a_n2224_n1088# 0.011024f
C99 minus.n26 a_n2224_n1088# 0.028931f
C100 minus.n27 a_n2224_n1088# 0.028931f
C101 minus.n28 a_n2224_n1088# 0.028931f
C102 minus.n29 a_n2224_n1088# 0.010132f
C103 minus.n30 a_n2224_n1088# 0.024458f
C104 minus.n31 a_n2224_n1088# 0.011024f
C105 minus.n32 a_n2224_n1088# 0.024458f
C106 minus.n33 a_n2224_n1088# 0.031811f
C107 minus.n34 a_n2224_n1088# 0.71419f
C108 minus.n35 a_n2224_n1088# 0.028931f
C109 minus.t15 a_n2224_n1088# 0.022296f
C110 minus.t11 a_n2224_n1088# 0.022296f
C111 minus.n36 a_n2224_n1088# 0.010489f
C112 minus.n37 a_n2224_n1088# 0.028931f
C113 minus.t7 a_n2224_n1088# 0.022296f
C114 minus.t8 a_n2224_n1088# 0.022296f
C115 minus.t12 a_n2224_n1088# 0.022296f
C116 minus.n38 a_n2224_n1088# 0.024458f
C117 minus.n39 a_n2224_n1088# 0.028931f
C118 minus.t5 a_n2224_n1088# 0.022296f
C119 minus.t23 a_n2224_n1088# 0.022296f
C120 minus.n40 a_n2224_n1088# 0.010132f
C121 minus.t6 a_n2224_n1088# 0.024898f
C122 minus.n41 a_n2224_n1088# 0.031847f
C123 minus.t22 a_n2224_n1088# 0.022296f
C124 minus.n42 a_n2224_n1088# 0.024458f
C125 minus.t0 a_n2224_n1088# 0.022296f
C126 minus.n43 a_n2224_n1088# 0.024458f
C127 minus.n44 a_n2224_n1088# 0.011024f
C128 minus.n45 a_n2224_n1088# 0.060144f
C129 minus.n46 a_n2224_n1088# 0.028931f
C130 minus.n47 a_n2224_n1088# 0.028931f
C131 minus.n48 a_n2224_n1088# 0.010489f
C132 minus.n49 a_n2224_n1088# 0.024458f
C133 minus.n50 a_n2224_n1088# 0.011024f
C134 minus.n51 a_n2224_n1088# 0.024458f
C135 minus.n52 a_n2224_n1088# 0.011024f
C136 minus.n53 a_n2224_n1088# 0.028931f
C137 minus.n54 a_n2224_n1088# 0.028931f
C138 minus.n55 a_n2224_n1088# 0.011024f
C139 minus.n56 a_n2224_n1088# 0.024458f
C140 minus.n57 a_n2224_n1088# 0.011024f
C141 minus.n58 a_n2224_n1088# 0.024458f
C142 minus.t4 a_n2224_n1088# 0.022296f
C143 minus.n59 a_n2224_n1088# 0.024458f
C144 minus.n60 a_n2224_n1088# 0.011024f
C145 minus.n61 a_n2224_n1088# 0.028931f
C146 minus.n62 a_n2224_n1088# 0.028931f
C147 minus.n63 a_n2224_n1088# 0.028931f
C148 minus.n64 a_n2224_n1088# 0.010132f
C149 minus.n65 a_n2224_n1088# 0.024458f
C150 minus.n66 a_n2224_n1088# 0.011024f
C151 minus.n67 a_n2224_n1088# 0.024458f
C152 minus.t14 a_n2224_n1088# 0.024898f
C153 minus.n68 a_n2224_n1088# 0.031811f
C154 minus.n69 a_n2224_n1088# 0.184513f
C155 minus.n70 a_n2224_n1088# 0.884575f
C156 drain_left.t6 a_n2224_n1088# 0.021801f
C157 drain_left.t4 a_n2224_n1088# 0.021801f
C158 drain_left.n0 a_n2224_n1088# 0.08532f
C159 drain_left.t2 a_n2224_n1088# 0.021801f
C160 drain_left.t0 a_n2224_n1088# 0.021801f
C161 drain_left.n1 a_n2224_n1088# 0.084711f
C162 drain_left.n2 a_n2224_n1088# 0.574142f
C163 drain_left.t5 a_n2224_n1088# 0.021801f
C164 drain_left.t10 a_n2224_n1088# 0.021801f
C165 drain_left.n3 a_n2224_n1088# 0.084711f
C166 drain_left.n4 a_n2224_n1088# 0.257962f
C167 drain_left.t17 a_n2224_n1088# 0.021801f
C168 drain_left.t12 a_n2224_n1088# 0.021801f
C169 drain_left.n5 a_n2224_n1088# 0.08532f
C170 drain_left.t3 a_n2224_n1088# 0.021801f
C171 drain_left.t8 a_n2224_n1088# 0.021801f
C172 drain_left.n6 a_n2224_n1088# 0.084711f
C173 drain_left.n7 a_n2224_n1088# 0.574142f
C174 drain_left.t7 a_n2224_n1088# 0.021801f
C175 drain_left.t13 a_n2224_n1088# 0.021801f
C176 drain_left.n8 a_n2224_n1088# 0.084711f
C177 drain_left.n9 a_n2224_n1088# 0.257962f
C178 drain_left.n10 a_n2224_n1088# 0.840007f
C179 drain_left.t18 a_n2224_n1088# 0.021801f
C180 drain_left.t22 a_n2224_n1088# 0.021801f
C181 drain_left.n11 a_n2224_n1088# 0.08532f
C182 drain_left.t14 a_n2224_n1088# 0.021801f
C183 drain_left.t23 a_n2224_n1088# 0.021801f
C184 drain_left.n12 a_n2224_n1088# 0.084711f
C185 drain_left.n13 a_n2224_n1088# 0.574142f
C186 drain_left.t15 a_n2224_n1088# 0.021801f
C187 drain_left.t1 a_n2224_n1088# 0.021801f
C188 drain_left.n14 a_n2224_n1088# 0.084711f
C189 drain_left.n15 a_n2224_n1088# 0.281819f
C190 drain_left.t16 a_n2224_n1088# 0.021801f
C191 drain_left.t19 a_n2224_n1088# 0.021801f
C192 drain_left.n16 a_n2224_n1088# 0.084711f
C193 drain_left.n17 a_n2224_n1088# 0.281819f
C194 drain_left.t9 a_n2224_n1088# 0.021801f
C195 drain_left.t20 a_n2224_n1088# 0.021801f
C196 drain_left.n18 a_n2224_n1088# 0.084711f
C197 drain_left.n19 a_n2224_n1088# 0.281819f
C198 drain_left.t11 a_n2224_n1088# 0.021801f
C199 drain_left.t21 a_n2224_n1088# 0.021801f
C200 drain_left.n20 a_n2224_n1088# 0.084711f
C201 drain_left.n21 a_n2224_n1088# 0.509539f
C202 source.t42 a_n2224_n1088# 0.145783f
C203 source.n0 a_n2224_n1088# 0.617716f
C204 source.t34 a_n2224_n1088# 0.026192f
C205 source.t28 a_n2224_n1088# 0.026192f
C206 source.n1 a_n2224_n1088# 0.084946f
C207 source.n2 a_n2224_n1088# 0.310368f
C208 source.t24 a_n2224_n1088# 0.026192f
C209 source.t25 a_n2224_n1088# 0.026192f
C210 source.n3 a_n2224_n1088# 0.084946f
C211 source.n4 a_n2224_n1088# 0.310368f
C212 source.t35 a_n2224_n1088# 0.026192f
C213 source.t30 a_n2224_n1088# 0.026192f
C214 source.n5 a_n2224_n1088# 0.084946f
C215 source.n6 a_n2224_n1088# 0.310368f
C216 source.t47 a_n2224_n1088# 0.026192f
C217 source.t40 a_n2224_n1088# 0.026192f
C218 source.n7 a_n2224_n1088# 0.084946f
C219 source.n8 a_n2224_n1088# 0.310368f
C220 source.t45 a_n2224_n1088# 0.026192f
C221 source.t32 a_n2224_n1088# 0.026192f
C222 source.n9 a_n2224_n1088# 0.084946f
C223 source.n10 a_n2224_n1088# 0.310368f
C224 source.t26 a_n2224_n1088# 0.145783f
C225 source.n11 a_n2224_n1088# 0.317743f
C226 source.t3 a_n2224_n1088# 0.145783f
C227 source.n12 a_n2224_n1088# 0.317743f
C228 source.t9 a_n2224_n1088# 0.026192f
C229 source.t20 a_n2224_n1088# 0.026192f
C230 source.n13 a_n2224_n1088# 0.084946f
C231 source.n14 a_n2224_n1088# 0.310368f
C232 source.t1 a_n2224_n1088# 0.026192f
C233 source.t16 a_n2224_n1088# 0.026192f
C234 source.n15 a_n2224_n1088# 0.084946f
C235 source.n16 a_n2224_n1088# 0.310368f
C236 source.t2 a_n2224_n1088# 0.026192f
C237 source.t12 a_n2224_n1088# 0.026192f
C238 source.n17 a_n2224_n1088# 0.084946f
C239 source.n18 a_n2224_n1088# 0.310368f
C240 source.t6 a_n2224_n1088# 0.026192f
C241 source.t13 a_n2224_n1088# 0.026192f
C242 source.n19 a_n2224_n1088# 0.084946f
C243 source.n20 a_n2224_n1088# 0.310368f
C244 source.t18 a_n2224_n1088# 0.026192f
C245 source.t23 a_n2224_n1088# 0.026192f
C246 source.n21 a_n2224_n1088# 0.084946f
C247 source.n22 a_n2224_n1088# 0.310368f
C248 source.t8 a_n2224_n1088# 0.145783f
C249 source.n23 a_n2224_n1088# 0.882355f
C250 source.t46 a_n2224_n1088# 0.145783f
C251 source.n24 a_n2224_n1088# 0.882355f
C252 source.t38 a_n2224_n1088# 0.026192f
C253 source.t36 a_n2224_n1088# 0.026192f
C254 source.n25 a_n2224_n1088# 0.084946f
C255 source.n26 a_n2224_n1088# 0.310368f
C256 source.t31 a_n2224_n1088# 0.026192f
C257 source.t44 a_n2224_n1088# 0.026192f
C258 source.n27 a_n2224_n1088# 0.084946f
C259 source.n28 a_n2224_n1088# 0.310368f
C260 source.t33 a_n2224_n1088# 0.026192f
C261 source.t39 a_n2224_n1088# 0.026192f
C262 source.n29 a_n2224_n1088# 0.084946f
C263 source.n30 a_n2224_n1088# 0.310368f
C264 source.t37 a_n2224_n1088# 0.026192f
C265 source.t43 a_n2224_n1088# 0.026192f
C266 source.n31 a_n2224_n1088# 0.084946f
C267 source.n32 a_n2224_n1088# 0.310368f
C268 source.t27 a_n2224_n1088# 0.026192f
C269 source.t29 a_n2224_n1088# 0.026192f
C270 source.n33 a_n2224_n1088# 0.084946f
C271 source.n34 a_n2224_n1088# 0.310368f
C272 source.t41 a_n2224_n1088# 0.145783f
C273 source.n35 a_n2224_n1088# 0.317743f
C274 source.t19 a_n2224_n1088# 0.145783f
C275 source.n36 a_n2224_n1088# 0.317743f
C276 source.t7 a_n2224_n1088# 0.026192f
C277 source.t5 a_n2224_n1088# 0.026192f
C278 source.n37 a_n2224_n1088# 0.084946f
C279 source.n38 a_n2224_n1088# 0.310368f
C280 source.t0 a_n2224_n1088# 0.026192f
C281 source.t15 a_n2224_n1088# 0.026192f
C282 source.n39 a_n2224_n1088# 0.084946f
C283 source.n40 a_n2224_n1088# 0.310368f
C284 source.t21 a_n2224_n1088# 0.026192f
C285 source.t14 a_n2224_n1088# 0.026192f
C286 source.n41 a_n2224_n1088# 0.084946f
C287 source.n42 a_n2224_n1088# 0.310368f
C288 source.t17 a_n2224_n1088# 0.026192f
C289 source.t4 a_n2224_n1088# 0.026192f
C290 source.n43 a_n2224_n1088# 0.084946f
C291 source.n44 a_n2224_n1088# 0.310368f
C292 source.t11 a_n2224_n1088# 0.026192f
C293 source.t10 a_n2224_n1088# 0.026192f
C294 source.n45 a_n2224_n1088# 0.084946f
C295 source.n46 a_n2224_n1088# 0.310368f
C296 source.t22 a_n2224_n1088# 0.145783f
C297 source.n47 a_n2224_n1088# 0.501162f
C298 source.n48 a_n2224_n1088# 0.669407f
C299 plus.n0 a_n2224_n1088# 0.029371f
C300 plus.t12 a_n2224_n1088# 0.022636f
C301 plus.t3 a_n2224_n1088# 0.022636f
C302 plus.n1 a_n2224_n1088# 0.010649f
C303 plus.n2 a_n2224_n1088# 0.029371f
C304 plus.t4 a_n2224_n1088# 0.022636f
C305 plus.t7 a_n2224_n1088# 0.022636f
C306 plus.t22 a_n2224_n1088# 0.022636f
C307 plus.n3 a_n2224_n1088# 0.024831f
C308 plus.n4 a_n2224_n1088# 0.029371f
C309 plus.t8 a_n2224_n1088# 0.022636f
C310 plus.t0 a_n2224_n1088# 0.022636f
C311 plus.n5 a_n2224_n1088# 0.010287f
C312 plus.t5 a_n2224_n1088# 0.025277f
C313 plus.n6 a_n2224_n1088# 0.032332f
C314 plus.t1 a_n2224_n1088# 0.022636f
C315 plus.n7 a_n2224_n1088# 0.024831f
C316 plus.t9 a_n2224_n1088# 0.022636f
C317 plus.n8 a_n2224_n1088# 0.024831f
C318 plus.n9 a_n2224_n1088# 0.011192f
C319 plus.n10 a_n2224_n1088# 0.06106f
C320 plus.n11 a_n2224_n1088# 0.029371f
C321 plus.n12 a_n2224_n1088# 0.029371f
C322 plus.n13 a_n2224_n1088# 0.010649f
C323 plus.n14 a_n2224_n1088# 0.024831f
C324 plus.n15 a_n2224_n1088# 0.011192f
C325 plus.n16 a_n2224_n1088# 0.024831f
C326 plus.n17 a_n2224_n1088# 0.011192f
C327 plus.n18 a_n2224_n1088# 0.029371f
C328 plus.n19 a_n2224_n1088# 0.029371f
C329 plus.n20 a_n2224_n1088# 0.011192f
C330 plus.n21 a_n2224_n1088# 0.024831f
C331 plus.n22 a_n2224_n1088# 0.011192f
C332 plus.n23 a_n2224_n1088# 0.024831f
C333 plus.t14 a_n2224_n1088# 0.022636f
C334 plus.n24 a_n2224_n1088# 0.024831f
C335 plus.n25 a_n2224_n1088# 0.011192f
C336 plus.n26 a_n2224_n1088# 0.029371f
C337 plus.n27 a_n2224_n1088# 0.029371f
C338 plus.n28 a_n2224_n1088# 0.029371f
C339 plus.n29 a_n2224_n1088# 0.010287f
C340 plus.n30 a_n2224_n1088# 0.024831f
C341 plus.n31 a_n2224_n1088# 0.011192f
C342 plus.n32 a_n2224_n1088# 0.024831f
C343 plus.t2 a_n2224_n1088# 0.025277f
C344 plus.n33 a_n2224_n1088# 0.032295f
C345 plus.n34 a_n2224_n1088# 0.19642f
C346 plus.n35 a_n2224_n1088# 0.029371f
C347 plus.t17 a_n2224_n1088# 0.025277f
C348 plus.t19 a_n2224_n1088# 0.022636f
C349 plus.t21 a_n2224_n1088# 0.022636f
C350 plus.n36 a_n2224_n1088# 0.010649f
C351 plus.n37 a_n2224_n1088# 0.029371f
C352 plus.t23 a_n2224_n1088# 0.022636f
C353 plus.n38 a_n2224_n1088# 0.024831f
C354 plus.t18 a_n2224_n1088# 0.022636f
C355 plus.t13 a_n2224_n1088# 0.022636f
C356 plus.t16 a_n2224_n1088# 0.022636f
C357 plus.n39 a_n2224_n1088# 0.024831f
C358 plus.n40 a_n2224_n1088# 0.029371f
C359 plus.t10 a_n2224_n1088# 0.022636f
C360 plus.t20 a_n2224_n1088# 0.022636f
C361 plus.n41 a_n2224_n1088# 0.010287f
C362 plus.t11 a_n2224_n1088# 0.025277f
C363 plus.n42 a_n2224_n1088# 0.032332f
C364 plus.t15 a_n2224_n1088# 0.022636f
C365 plus.n43 a_n2224_n1088# 0.024831f
C366 plus.t6 a_n2224_n1088# 0.022636f
C367 plus.n44 a_n2224_n1088# 0.024831f
C368 plus.n45 a_n2224_n1088# 0.011192f
C369 plus.n46 a_n2224_n1088# 0.06106f
C370 plus.n47 a_n2224_n1088# 0.029371f
C371 plus.n48 a_n2224_n1088# 0.029371f
C372 plus.n49 a_n2224_n1088# 0.010649f
C373 plus.n50 a_n2224_n1088# 0.024831f
C374 plus.n51 a_n2224_n1088# 0.011192f
C375 plus.n52 a_n2224_n1088# 0.024831f
C376 plus.n53 a_n2224_n1088# 0.011192f
C377 plus.n54 a_n2224_n1088# 0.029371f
C378 plus.n55 a_n2224_n1088# 0.029371f
C379 plus.n56 a_n2224_n1088# 0.011192f
C380 plus.n57 a_n2224_n1088# 0.024831f
C381 plus.n58 a_n2224_n1088# 0.011192f
C382 plus.n59 a_n2224_n1088# 0.024831f
C383 plus.n60 a_n2224_n1088# 0.011192f
C384 plus.n61 a_n2224_n1088# 0.029371f
C385 plus.n62 a_n2224_n1088# 0.029371f
C386 plus.n63 a_n2224_n1088# 0.029371f
C387 plus.n64 a_n2224_n1088# 0.010287f
C388 plus.n65 a_n2224_n1088# 0.024831f
C389 plus.n66 a_n2224_n1088# 0.011192f
C390 plus.n67 a_n2224_n1088# 0.024831f
C391 plus.n68 a_n2224_n1088# 0.032295f
C392 plus.n69 a_n2224_n1088# 0.700613f
.ends

