* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_right.t9 minus.t0 source.t16 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X1 source.t5 plus.t0 drain_left.t9 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X2 drain_right.t8 minus.t1 source.t13 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X3 a_n1472_n1288# a_n1472_n1288# a_n1472_n1288# a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.3
X4 source.t10 minus.t2 drain_right.t7 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X5 drain_left.t8 plus.t1 source.t7 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X6 drain_left.t7 plus.t2 source.t6 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X7 drain_left.t6 plus.t3 source.t0 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X8 source.t4 plus.t4 drain_left.t5 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X9 drain_right.t6 minus.t3 source.t15 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X10 source.t1 plus.t5 drain_left.t4 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X11 source.t17 minus.t4 drain_right.t5 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X12 a_n1472_n1288# a_n1472_n1288# a_n1472_n1288# a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X13 drain_right.t4 minus.t5 source.t14 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X14 source.t12 minus.t6 drain_right.t3 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X15 drain_left.t3 plus.t6 source.t3 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X16 drain_left.t2 plus.t7 source.t2 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X17 drain_right.t2 minus.t7 source.t11 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X18 drain_right.t1 minus.t8 source.t9 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X19 source.t8 minus.t9 drain_right.t0 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X20 a_n1472_n1288# a_n1472_n1288# a_n1472_n1288# a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X21 drain_left.t1 plus.t8 source.t18 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X22 source.t19 plus.t9 drain_left.t0 a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X23 a_n1472_n1288# a_n1472_n1288# a_n1472_n1288# a_n1472_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
R0 minus.n9 minus.t8 303.077
R1 minus.n3 minus.t5 303.077
R2 minus.n20 minus.t7 303.077
R3 minus.n14 minus.t0 303.077
R4 minus.n6 minus.t1 265.101
R5 minus.n8 minus.t4 265.101
R6 minus.n2 minus.t9 265.101
R7 minus.n17 minus.t3 265.101
R8 minus.n19 minus.t2 265.101
R9 minus.n13 minus.t6 265.101
R10 minus.n4 minus.n3 161.489
R11 minus.n15 minus.n14 161.489
R12 minus.n10 minus.n9 161.3
R13 minus.n7 minus.n0 161.3
R14 minus.n6 minus.n5 161.3
R15 minus.n4 minus.n1 161.3
R16 minus.n21 minus.n20 161.3
R17 minus.n18 minus.n11 161.3
R18 minus.n17 minus.n16 161.3
R19 minus.n15 minus.n12 161.3
R20 minus.n7 minus.n6 73.0308
R21 minus.n6 minus.n1 73.0308
R22 minus.n17 minus.n12 73.0308
R23 minus.n18 minus.n17 73.0308
R24 minus.n9 minus.n8 54.0429
R25 minus.n3 minus.n2 54.0429
R26 minus.n14 minus.n13 54.0429
R27 minus.n20 minus.n19 54.0429
R28 minus.n22 minus.n10 27.1085
R29 minus.n8 minus.n7 18.9884
R30 minus.n2 minus.n1 18.9884
R31 minus.n13 minus.n12 18.9884
R32 minus.n19 minus.n18 18.9884
R33 minus.n22 minus.n21 6.48724
R34 minus.n10 minus.n0 0.189894
R35 minus.n5 minus.n0 0.189894
R36 minus.n5 minus.n4 0.189894
R37 minus.n16 minus.n15 0.189894
R38 minus.n16 minus.n11 0.189894
R39 minus.n21 minus.n11 0.189894
R40 minus minus.n22 0.188
R41 source.n42 source.n40 289.615
R42 source.n30 source.n28 289.615
R43 source.n2 source.n0 289.615
R44 source.n14 source.n12 289.615
R45 source.n43 source.n42 185
R46 source.n31 source.n30 185
R47 source.n3 source.n2 185
R48 source.n15 source.n14 185
R49 source.t11 source.n41 167.117
R50 source.t18 source.n29 167.117
R51 source.t0 source.n1 167.117
R52 source.t14 source.n13 167.117
R53 source.n9 source.n8 84.1169
R54 source.n11 source.n10 84.1169
R55 source.n21 source.n20 84.1169
R56 source.n23 source.n22 84.1169
R57 source.n39 source.n38 84.1168
R58 source.n37 source.n36 84.1168
R59 source.n27 source.n26 84.1168
R60 source.n25 source.n24 84.1168
R61 source.n42 source.t11 52.3082
R62 source.n30 source.t18 52.3082
R63 source.n2 source.t0 52.3082
R64 source.n14 source.t14 52.3082
R65 source.n47 source.n46 31.4096
R66 source.n35 source.n34 31.4096
R67 source.n7 source.n6 31.4096
R68 source.n19 source.n18 31.4096
R69 source.n25 source.n23 14.7982
R70 source.n38 source.t15 9.9005
R71 source.n38 source.t10 9.9005
R72 source.n36 source.t16 9.9005
R73 source.n36 source.t12 9.9005
R74 source.n26 source.t6 9.9005
R75 source.n26 source.t1 9.9005
R76 source.n24 source.t3 9.9005
R77 source.n24 source.t5 9.9005
R78 source.n8 source.t2 9.9005
R79 source.n8 source.t19 9.9005
R80 source.n10 source.t7 9.9005
R81 source.n10 source.t4 9.9005
R82 source.n20 source.t13 9.9005
R83 source.n20 source.t8 9.9005
R84 source.n22 source.t9 9.9005
R85 source.n22 source.t17 9.9005
R86 source.n43 source.n41 9.71174
R87 source.n31 source.n29 9.71174
R88 source.n3 source.n1 9.71174
R89 source.n15 source.n13 9.71174
R90 source.n46 source.n45 9.45567
R91 source.n34 source.n33 9.45567
R92 source.n6 source.n5 9.45567
R93 source.n18 source.n17 9.45567
R94 source.n45 source.n44 9.3005
R95 source.n33 source.n32 9.3005
R96 source.n5 source.n4 9.3005
R97 source.n17 source.n16 9.3005
R98 source.n48 source.n7 8.72059
R99 source.n46 source.n40 8.14595
R100 source.n34 source.n28 8.14595
R101 source.n6 source.n0 8.14595
R102 source.n18 source.n12 8.14595
R103 source.n44 source.n43 7.3702
R104 source.n32 source.n31 7.3702
R105 source.n4 source.n3 7.3702
R106 source.n16 source.n15 7.3702
R107 source.n44 source.n40 5.81868
R108 source.n32 source.n28 5.81868
R109 source.n4 source.n0 5.81868
R110 source.n16 source.n12 5.81868
R111 source.n48 source.n47 5.53498
R112 source.n45 source.n41 3.44771
R113 source.n33 source.n29 3.44771
R114 source.n5 source.n1 3.44771
R115 source.n17 source.n13 3.44771
R116 source.n19 source.n11 0.741879
R117 source.n37 source.n35 0.741879
R118 source.n23 source.n21 0.543603
R119 source.n21 source.n19 0.543603
R120 source.n11 source.n9 0.543603
R121 source.n9 source.n7 0.543603
R122 source.n27 source.n25 0.543603
R123 source.n35 source.n27 0.543603
R124 source.n39 source.n37 0.543603
R125 source.n47 source.n39 0.543603
R126 source source.n48 0.188
R127 drain_right.n2 drain_right.n0 289.615
R128 drain_right.n16 drain_right.n14 289.615
R129 drain_right.n3 drain_right.n2 185
R130 drain_right.n17 drain_right.n16 185
R131 drain_right.t9 drain_right.n1 167.117
R132 drain_right.t1 drain_right.n15 167.117
R133 drain_right.n13 drain_right.n11 101.338
R134 drain_right.n10 drain_right.n9 101.147
R135 drain_right.n13 drain_right.n12 100.796
R136 drain_right.n8 drain_right.n7 100.796
R137 drain_right.n2 drain_right.t9 52.3082
R138 drain_right.n16 drain_right.t1 52.3082
R139 drain_right.n8 drain_right.n6 48.6315
R140 drain_right.n21 drain_right.n20 48.0884
R141 drain_right drain_right.n10 21.5463
R142 drain_right.n9 drain_right.t7 9.9005
R143 drain_right.n9 drain_right.t2 9.9005
R144 drain_right.n7 drain_right.t3 9.9005
R145 drain_right.n7 drain_right.t6 9.9005
R146 drain_right.n11 drain_right.t0 9.9005
R147 drain_right.n11 drain_right.t4 9.9005
R148 drain_right.n12 drain_right.t5 9.9005
R149 drain_right.n12 drain_right.t8 9.9005
R150 drain_right.n3 drain_right.n1 9.71174
R151 drain_right.n17 drain_right.n15 9.71174
R152 drain_right.n6 drain_right.n5 9.45567
R153 drain_right.n20 drain_right.n19 9.45567
R154 drain_right.n5 drain_right.n4 9.3005
R155 drain_right.n19 drain_right.n18 9.3005
R156 drain_right.n6 drain_right.n0 8.14595
R157 drain_right.n20 drain_right.n14 8.14595
R158 drain_right.n4 drain_right.n3 7.3702
R159 drain_right.n18 drain_right.n17 7.3702
R160 drain_right drain_right.n21 5.92477
R161 drain_right.n4 drain_right.n0 5.81868
R162 drain_right.n18 drain_right.n14 5.81868
R163 drain_right.n5 drain_right.n1 3.44771
R164 drain_right.n19 drain_right.n15 3.44771
R165 drain_right.n21 drain_right.n13 0.543603
R166 drain_right.n10 drain_right.n8 0.0809298
R167 plus.n3 plus.t1 303.077
R168 plus.n9 plus.t3 303.077
R169 plus.n14 plus.t8 303.077
R170 plus.n20 plus.t6 303.077
R171 plus.n6 plus.t7 265.101
R172 plus.n2 plus.t4 265.101
R173 plus.n8 plus.t9 265.101
R174 plus.n17 plus.t2 265.101
R175 plus.n13 plus.t5 265.101
R176 plus.n19 plus.t0 265.101
R177 plus.n4 plus.n3 161.489
R178 plus.n15 plus.n14 161.489
R179 plus.n4 plus.n1 161.3
R180 plus.n6 plus.n5 161.3
R181 plus.n7 plus.n0 161.3
R182 plus.n10 plus.n9 161.3
R183 plus.n15 plus.n12 161.3
R184 plus.n17 plus.n16 161.3
R185 plus.n18 plus.n11 161.3
R186 plus.n21 plus.n20 161.3
R187 plus.n6 plus.n1 73.0308
R188 plus.n7 plus.n6 73.0308
R189 plus.n18 plus.n17 73.0308
R190 plus.n17 plus.n12 73.0308
R191 plus.n3 plus.n2 54.0429
R192 plus.n9 plus.n8 54.0429
R193 plus.n20 plus.n19 54.0429
R194 plus.n14 plus.n13 54.0429
R195 plus plus.n21 24.7774
R196 plus.n2 plus.n1 18.9884
R197 plus.n8 plus.n7 18.9884
R198 plus.n19 plus.n18 18.9884
R199 plus.n13 plus.n12 18.9884
R200 plus plus.n10 8.3433
R201 plus.n5 plus.n4 0.189894
R202 plus.n5 plus.n0 0.189894
R203 plus.n10 plus.n0 0.189894
R204 plus.n21 plus.n11 0.189894
R205 plus.n16 plus.n11 0.189894
R206 plus.n16 plus.n15 0.189894
R207 drain_left.n2 drain_left.n0 289.615
R208 drain_left.n13 drain_left.n11 289.615
R209 drain_left.n3 drain_left.n2 185
R210 drain_left.n14 drain_left.n13 185
R211 drain_left.t3 drain_left.n1 167.117
R212 drain_left.t8 drain_left.n12 167.117
R213 drain_left.n10 drain_left.n9 101.147
R214 drain_left.n21 drain_left.n20 100.796
R215 drain_left.n19 drain_left.n18 100.796
R216 drain_left.n8 drain_left.n7 100.796
R217 drain_left.n2 drain_left.t3 52.3082
R218 drain_left.n13 drain_left.t8 52.3082
R219 drain_left.n8 drain_left.n6 48.6315
R220 drain_left.n19 drain_left.n17 48.6315
R221 drain_left drain_left.n10 22.0995
R222 drain_left.n9 drain_left.t4 9.9005
R223 drain_left.n9 drain_left.t1 9.9005
R224 drain_left.n7 drain_left.t9 9.9005
R225 drain_left.n7 drain_left.t7 9.9005
R226 drain_left.n20 drain_left.t0 9.9005
R227 drain_left.n20 drain_left.t6 9.9005
R228 drain_left.n18 drain_left.t5 9.9005
R229 drain_left.n18 drain_left.t2 9.9005
R230 drain_left.n3 drain_left.n1 9.71174
R231 drain_left.n14 drain_left.n12 9.71174
R232 drain_left.n6 drain_left.n5 9.45567
R233 drain_left.n17 drain_left.n16 9.45567
R234 drain_left.n5 drain_left.n4 9.3005
R235 drain_left.n16 drain_left.n15 9.3005
R236 drain_left.n6 drain_left.n0 8.14595
R237 drain_left.n17 drain_left.n11 8.14595
R238 drain_left.n4 drain_left.n3 7.3702
R239 drain_left.n15 drain_left.n14 7.3702
R240 drain_left drain_left.n21 6.19632
R241 drain_left.n4 drain_left.n0 5.81868
R242 drain_left.n15 drain_left.n11 5.81868
R243 drain_left.n5 drain_left.n1 3.44771
R244 drain_left.n16 drain_left.n12 3.44771
R245 drain_left.n21 drain_left.n19 0.543603
R246 drain_left.n10 drain_left.n8 0.0809298
C0 drain_left drain_right 0.72073f
C1 drain_left plus 1.13324f
C2 drain_left minus 0.177605f
C3 drain_right source 5.29465f
C4 plus source 1.12913f
C5 minus source 1.11506f
C6 drain_right plus 0.30186f
C7 drain_right minus 0.99334f
C8 plus minus 3.14368f
C9 drain_left source 5.29756f
C10 drain_right a_n1472_n1288# 3.51251f
C11 drain_left a_n1472_n1288# 3.72178f
C12 source a_n1472_n1288# 2.43248f
C13 minus a_n1472_n1288# 4.896002f
C14 plus a_n1472_n1288# 5.544253f
C15 drain_left.n0 a_n1472_n1288# 0.033862f
C16 drain_left.n1 a_n1472_n1288# 0.074924f
C17 drain_left.t3 a_n1472_n1288# 0.056226f
C18 drain_left.n2 a_n1472_n1288# 0.058638f
C19 drain_left.n3 a_n1472_n1288# 0.018903f
C20 drain_left.n4 a_n1472_n1288# 0.012467f
C21 drain_left.n5 a_n1472_n1288# 0.16515f
C22 drain_left.n6 a_n1472_n1288# 0.054094f
C23 drain_left.t9 a_n1472_n1288# 0.036667f
C24 drain_left.t7 a_n1472_n1288# 0.036667f
C25 drain_left.n7 a_n1472_n1288# 0.230352f
C26 drain_left.n8 a_n1472_n1288# 0.314475f
C27 drain_left.t4 a_n1472_n1288# 0.036667f
C28 drain_left.t1 a_n1472_n1288# 0.036667f
C29 drain_left.n9 a_n1472_n1288# 0.23124f
C30 drain_left.n10 a_n1472_n1288# 0.828149f
C31 drain_left.n11 a_n1472_n1288# 0.033862f
C32 drain_left.n12 a_n1472_n1288# 0.074924f
C33 drain_left.t8 a_n1472_n1288# 0.056226f
C34 drain_left.n13 a_n1472_n1288# 0.058638f
C35 drain_left.n14 a_n1472_n1288# 0.018903f
C36 drain_left.n15 a_n1472_n1288# 0.012467f
C37 drain_left.n16 a_n1472_n1288# 0.16515f
C38 drain_left.n17 a_n1472_n1288# 0.054094f
C39 drain_left.t5 a_n1472_n1288# 0.036667f
C40 drain_left.t2 a_n1472_n1288# 0.036667f
C41 drain_left.n18 a_n1472_n1288# 0.230353f
C42 drain_left.n19 a_n1472_n1288# 0.342374f
C43 drain_left.t0 a_n1472_n1288# 0.036667f
C44 drain_left.t6 a_n1472_n1288# 0.036667f
C45 drain_left.n20 a_n1472_n1288# 0.230353f
C46 drain_left.n21 a_n1472_n1288# 0.451878f
C47 plus.n0 a_n1472_n1288# 0.032187f
C48 plus.t9 a_n1472_n1288# 0.056828f
C49 plus.t7 a_n1472_n1288# 0.056828f
C50 plus.n1 a_n1472_n1288# 0.013257f
C51 plus.t1 a_n1472_n1288# 0.06195f
C52 plus.t4 a_n1472_n1288# 0.056828f
C53 plus.n2 a_n1472_n1288# 0.039689f
C54 plus.n3 a_n1472_n1288# 0.04906f
C55 plus.n4 a_n1472_n1288# 0.070679f
C56 plus.n5 a_n1472_n1288# 0.032187f
C57 plus.n6 a_n1472_n1288# 0.050367f
C58 plus.n7 a_n1472_n1288# 0.013257f
C59 plus.n8 a_n1472_n1288# 0.039689f
C60 plus.t3 a_n1472_n1288# 0.06195f
C61 plus.n9 a_n1472_n1288# 0.049015f
C62 plus.n10 a_n1472_n1288# 0.229081f
C63 plus.n11 a_n1472_n1288# 0.032187f
C64 plus.t6 a_n1472_n1288# 0.06195f
C65 plus.t0 a_n1472_n1288# 0.056828f
C66 plus.t2 a_n1472_n1288# 0.056828f
C67 plus.n12 a_n1472_n1288# 0.013257f
C68 plus.t5 a_n1472_n1288# 0.056828f
C69 plus.n13 a_n1472_n1288# 0.039689f
C70 plus.t8 a_n1472_n1288# 0.06195f
C71 plus.n14 a_n1472_n1288# 0.04906f
C72 plus.n15 a_n1472_n1288# 0.070679f
C73 plus.n16 a_n1472_n1288# 0.032187f
C74 plus.n17 a_n1472_n1288# 0.050367f
C75 plus.n18 a_n1472_n1288# 0.013257f
C76 plus.n19 a_n1472_n1288# 0.039689f
C77 plus.n20 a_n1472_n1288# 0.049015f
C78 plus.n21 a_n1472_n1288# 0.671517f
C79 drain_right.n0 a_n1472_n1288# 0.034452f
C80 drain_right.n1 a_n1472_n1288# 0.076229f
C81 drain_right.t9 a_n1472_n1288# 0.057206f
C82 drain_right.n2 a_n1472_n1288# 0.05966f
C83 drain_right.n3 a_n1472_n1288# 0.019232f
C84 drain_right.n4 a_n1472_n1288# 0.012684f
C85 drain_right.n5 a_n1472_n1288# 0.168027f
C86 drain_right.n6 a_n1472_n1288# 0.055037f
C87 drain_right.t3 a_n1472_n1288# 0.037306f
C88 drain_right.t6 a_n1472_n1288# 0.037306f
C89 drain_right.n7 a_n1472_n1288# 0.234365f
C90 drain_right.n8 a_n1472_n1288# 0.319954f
C91 drain_right.t7 a_n1472_n1288# 0.037306f
C92 drain_right.t2 a_n1472_n1288# 0.037306f
C93 drain_right.n9 a_n1472_n1288# 0.235269f
C94 drain_right.n10 a_n1472_n1288# 0.79616f
C95 drain_right.t0 a_n1472_n1288# 0.037306f
C96 drain_right.t4 a_n1472_n1288# 0.037306f
C97 drain_right.n11 a_n1472_n1288# 0.235828f
C98 drain_right.t5 a_n1472_n1288# 0.037306f
C99 drain_right.t8 a_n1472_n1288# 0.037306f
C100 drain_right.n12 a_n1472_n1288# 0.234366f
C101 drain_right.n13 a_n1472_n1288# 0.534603f
C102 drain_right.n14 a_n1472_n1288# 0.034452f
C103 drain_right.n15 a_n1472_n1288# 0.076229f
C104 drain_right.t1 a_n1472_n1288# 0.057206f
C105 drain_right.n16 a_n1472_n1288# 0.05966f
C106 drain_right.n17 a_n1472_n1288# 0.019232f
C107 drain_right.n18 a_n1472_n1288# 0.012684f
C108 drain_right.n19 a_n1472_n1288# 0.168027f
C109 drain_right.n20 a_n1472_n1288# 0.054076f
C110 drain_right.n21 a_n1472_n1288# 0.282939f
C111 source.n0 a_n1472_n1288# 0.042035f
C112 source.n1 a_n1472_n1288# 0.093008f
C113 source.t0 a_n1472_n1288# 0.069798f
C114 source.n2 a_n1472_n1288# 0.072792f
C115 source.n3 a_n1472_n1288# 0.023465f
C116 source.n4 a_n1472_n1288# 0.015476f
C117 source.n5 a_n1472_n1288# 0.205014f
C118 source.n6 a_n1472_n1288# 0.046081f
C119 source.n7 a_n1472_n1288# 0.434834f
C120 source.t2 a_n1472_n1288# 0.045517f
C121 source.t19 a_n1472_n1288# 0.045517f
C122 source.n8 a_n1472_n1288# 0.243334f
C123 source.n9 a_n1472_n1288# 0.324707f
C124 source.t7 a_n1472_n1288# 0.045517f
C125 source.t4 a_n1472_n1288# 0.045517f
C126 source.n10 a_n1472_n1288# 0.243334f
C127 source.n11 a_n1472_n1288# 0.343107f
C128 source.n12 a_n1472_n1288# 0.042035f
C129 source.n13 a_n1472_n1288# 0.093008f
C130 source.t14 a_n1472_n1288# 0.069798f
C131 source.n14 a_n1472_n1288# 0.072792f
C132 source.n15 a_n1472_n1288# 0.023465f
C133 source.n16 a_n1472_n1288# 0.015476f
C134 source.n17 a_n1472_n1288# 0.205014f
C135 source.n18 a_n1472_n1288# 0.046081f
C136 source.n19 a_n1472_n1288# 0.14291f
C137 source.t13 a_n1472_n1288# 0.045517f
C138 source.t8 a_n1472_n1288# 0.045517f
C139 source.n20 a_n1472_n1288# 0.243334f
C140 source.n21 a_n1472_n1288# 0.324707f
C141 source.t9 a_n1472_n1288# 0.045517f
C142 source.t17 a_n1472_n1288# 0.045517f
C143 source.n22 a_n1472_n1288# 0.243334f
C144 source.n23 a_n1472_n1288# 0.953935f
C145 source.t3 a_n1472_n1288# 0.045517f
C146 source.t5 a_n1472_n1288# 0.045517f
C147 source.n24 a_n1472_n1288# 0.243333f
C148 source.n25 a_n1472_n1288# 0.953936f
C149 source.t6 a_n1472_n1288# 0.045517f
C150 source.t1 a_n1472_n1288# 0.045517f
C151 source.n26 a_n1472_n1288# 0.243333f
C152 source.n27 a_n1472_n1288# 0.324709f
C153 source.n28 a_n1472_n1288# 0.042035f
C154 source.n29 a_n1472_n1288# 0.093008f
C155 source.t18 a_n1472_n1288# 0.069798f
C156 source.n30 a_n1472_n1288# 0.072792f
C157 source.n31 a_n1472_n1288# 0.023465f
C158 source.n32 a_n1472_n1288# 0.015476f
C159 source.n33 a_n1472_n1288# 0.205014f
C160 source.n34 a_n1472_n1288# 0.046081f
C161 source.n35 a_n1472_n1288# 0.14291f
C162 source.t16 a_n1472_n1288# 0.045517f
C163 source.t12 a_n1472_n1288# 0.045517f
C164 source.n36 a_n1472_n1288# 0.243333f
C165 source.n37 a_n1472_n1288# 0.343109f
C166 source.t15 a_n1472_n1288# 0.045517f
C167 source.t10 a_n1472_n1288# 0.045517f
C168 source.n38 a_n1472_n1288# 0.243333f
C169 source.n39 a_n1472_n1288# 0.324709f
C170 source.n40 a_n1472_n1288# 0.042035f
C171 source.n41 a_n1472_n1288# 0.093008f
C172 source.t11 a_n1472_n1288# 0.069798f
C173 source.n42 a_n1472_n1288# 0.072792f
C174 source.n43 a_n1472_n1288# 0.023465f
C175 source.n44 a_n1472_n1288# 0.015476f
C176 source.n45 a_n1472_n1288# 0.205014f
C177 source.n46 a_n1472_n1288# 0.046081f
C178 source.n47 a_n1472_n1288# 0.280285f
C179 source.n48 a_n1472_n1288# 0.71204f
C180 minus.n0 a_n1472_n1288# 0.031525f
C181 minus.t8 a_n1472_n1288# 0.060676f
C182 minus.t4 a_n1472_n1288# 0.055659f
C183 minus.t1 a_n1472_n1288# 0.055659f
C184 minus.n1 a_n1472_n1288# 0.012985f
C185 minus.t9 a_n1472_n1288# 0.055659f
C186 minus.n2 a_n1472_n1288# 0.038873f
C187 minus.t5 a_n1472_n1288# 0.060676f
C188 minus.n3 a_n1472_n1288# 0.048051f
C189 minus.n4 a_n1472_n1288# 0.069225f
C190 minus.n5 a_n1472_n1288# 0.031525f
C191 minus.n6 a_n1472_n1288# 0.049331f
C192 minus.n7 a_n1472_n1288# 0.012985f
C193 minus.n8 a_n1472_n1288# 0.038873f
C194 minus.n9 a_n1472_n1288# 0.048007f
C195 minus.n10 a_n1472_n1288# 0.686138f
C196 minus.n11 a_n1472_n1288# 0.031525f
C197 minus.t2 a_n1472_n1288# 0.055659f
C198 minus.t3 a_n1472_n1288# 0.055659f
C199 minus.n12 a_n1472_n1288# 0.012985f
C200 minus.t0 a_n1472_n1288# 0.060676f
C201 minus.t6 a_n1472_n1288# 0.055659f
C202 minus.n13 a_n1472_n1288# 0.038873f
C203 minus.n14 a_n1472_n1288# 0.048051f
C204 minus.n15 a_n1472_n1288# 0.069225f
C205 minus.n16 a_n1472_n1288# 0.031525f
C206 minus.n17 a_n1472_n1288# 0.049331f
C207 minus.n18 a_n1472_n1288# 0.012985f
C208 minus.n19 a_n1472_n1288# 0.038873f
C209 minus.t7 a_n1472_n1288# 0.060676f
C210 minus.n20 a_n1472_n1288# 0.048007f
C211 minus.n21 a_n1472_n1288# 0.205154f
C212 minus.n22 a_n1472_n1288# 0.848591f
.ends

