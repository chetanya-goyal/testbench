* NGSPICE file created from diffpair671.ext - technology: sky130A

.subckt diffpair671 minus drain_right drain_left source plus
X0 drain_right minus source a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X1 source plus drain_left a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X2 drain_right minus source a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X3 source minus drain_right a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X4 a_n1094_n5892# a_n1094_n5892# a_n1094_n5892# a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.3
X5 drain_left plus source a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X6 a_n1094_n5892# a_n1094_n5892# a_n1094_n5892# a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X7 source minus drain_right a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X8 a_n1094_n5892# a_n1094_n5892# a_n1094_n5892# a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X9 source plus drain_left a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X10 a_n1094_n5892# a_n1094_n5892# a_n1094_n5892# a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X11 drain_left plus source a_n1094_n5892# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
.ends

