* NGSPICE file created from diffpair643.ext - technology: sky130A

.subckt diffpair643 minus drain_right drain_left source plus
X0 drain_right.t7 minus.t0 source.t13 a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X1 a_n1366_n5888# a_n1366_n5888# a_n1366_n5888# a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=95 ps=407.6 w=25 l=0.15
X2 source.t10 minus.t1 drain_right.t6 a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X3 drain_left.t7 plus.t0 source.t14 a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X4 a_n1366_n5888# a_n1366_n5888# a_n1366_n5888# a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X5 source.t12 minus.t2 drain_right.t5 a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X6 a_n1366_n5888# a_n1366_n5888# a_n1366_n5888# a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X7 source.t15 plus.t1 drain_left.t6 a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X8 drain_right.t4 minus.t3 source.t9 a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X9 drain_left.t5 plus.t2 source.t1 a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X10 a_n1366_n5888# a_n1366_n5888# a_n1366_n5888# a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=0 ps=0 w=25 l=0.15
X11 source.t8 minus.t4 drain_right.t3 a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X12 source.t0 plus.t3 drain_left.t4 a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=11.875 pd=50.95 as=6.25 ps=25.5 w=25 l=0.15
X13 drain_right.t2 minus.t5 source.t7 a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X14 drain_right.t1 minus.t6 source.t11 a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X15 drain_left.t3 plus.t4 source.t4 a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=11.875 ps=50.95 w=25 l=0.15
X16 source.t2 plus.t5 drain_left.t2 a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X17 source.t5 plus.t6 drain_left.t1 a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X18 drain_left.t0 plus.t7 source.t3 a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
X19 source.t6 minus.t7 drain_right.t0 a_n1366_n5888# sky130_fd_pr__nfet_01v8 ad=6.25 pd=25.5 as=6.25 ps=25.5 w=25 l=0.15
R0 minus.n5 minus.t4 4294.91
R1 minus.n1 minus.t3 4294.91
R2 minus.n12 minus.t0 4294.91
R3 minus.n8 minus.t1 4294.91
R4 minus.n4 minus.t5 4225.53
R5 minus.n2 minus.t2 4225.53
R6 minus.n11 minus.t7 4225.53
R7 minus.n9 minus.t6 4225.53
R8 minus.n1 minus.n0 161.489
R9 minus.n8 minus.n7 161.489
R10 minus.n6 minus.n5 161.3
R11 minus.n3 minus.n0 161.3
R12 minus.n13 minus.n12 161.3
R13 minus.n10 minus.n7 161.3
R14 minus.n4 minus.n3 47.4702
R15 minus.n3 minus.n2 47.4702
R16 minus.n10 minus.n9 47.4702
R17 minus.n11 minus.n10 47.4702
R18 minus.n14 minus.n6 44.224
R19 minus.n5 minus.n4 25.5611
R20 minus.n2 minus.n1 25.5611
R21 minus.n9 minus.n8 25.5611
R22 minus.n12 minus.n11 25.5611
R23 minus.n14 minus.n13 6.58005
R24 minus.n6 minus.n0 0.189894
R25 minus.n13 minus.n7 0.189894
R26 minus minus.n14 0.188
R27 source.n3 source.t0 43.2366
R28 source.n4 source.t9 43.2366
R29 source.n7 source.t8 43.2366
R30 source.n15 source.t13 43.2365
R31 source.n12 source.t10 43.2365
R32 source.n11 source.t1 43.2365
R33 source.n8 source.t15 43.2365
R34 source.n0 source.t4 43.2365
R35 source.n14 source.n13 42.0366
R36 source.n10 source.n9 42.0366
R37 source.n2 source.n1 42.0366
R38 source.n6 source.n5 42.0366
R39 source.n8 source.n7 31.6966
R40 source.n16 source.n0 26.1535
R41 source.n16 source.n15 5.5436
R42 source.n13 source.t11 1.2005
R43 source.n13 source.t6 1.2005
R44 source.n9 source.t14 1.2005
R45 source.n9 source.t2 1.2005
R46 source.n1 source.t3 1.2005
R47 source.n1 source.t5 1.2005
R48 source.n5 source.t7 1.2005
R49 source.n5 source.t12 1.2005
R50 source.n7 source.n6 0.560845
R51 source.n6 source.n4 0.560845
R52 source.n3 source.n2 0.560845
R53 source.n2 source.n0 0.560845
R54 source.n10 source.n8 0.560845
R55 source.n11 source.n10 0.560845
R56 source.n14 source.n12 0.560845
R57 source.n15 source.n14 0.560845
R58 source.n4 source.n3 0.470328
R59 source.n12 source.n11 0.470328
R60 source source.n16 0.188
R61 drain_right.n5 drain_right.n3 59.2756
R62 drain_right.n2 drain_right.n1 58.9403
R63 drain_right.n2 drain_right.n0 58.9403
R64 drain_right.n5 drain_right.n4 58.7154
R65 drain_right drain_right.n2 38.6235
R66 drain_right drain_right.n5 6.21356
R67 drain_right.n1 drain_right.t0 1.2005
R68 drain_right.n1 drain_right.t7 1.2005
R69 drain_right.n0 drain_right.t6 1.2005
R70 drain_right.n0 drain_right.t1 1.2005
R71 drain_right.n3 drain_right.t5 1.2005
R72 drain_right.n3 drain_right.t4 1.2005
R73 drain_right.n4 drain_right.t3 1.2005
R74 drain_right.n4 drain_right.t2 1.2005
R75 plus.n1 plus.t3 4294.91
R76 plus.n5 plus.t4 4294.91
R77 plus.n8 plus.t2 4294.91
R78 plus.n12 plus.t1 4294.91
R79 plus.n2 plus.t7 4225.53
R80 plus.n4 plus.t6 4225.53
R81 plus.n9 plus.t5 4225.53
R82 plus.n11 plus.t0 4225.53
R83 plus.n1 plus.n0 161.489
R84 plus.n8 plus.n7 161.489
R85 plus.n3 plus.n0 161.3
R86 plus.n6 plus.n5 161.3
R87 plus.n10 plus.n7 161.3
R88 plus.n13 plus.n12 161.3
R89 plus.n3 plus.n2 47.4702
R90 plus.n4 plus.n3 47.4702
R91 plus.n11 plus.n10 47.4702
R92 plus.n10 plus.n9 47.4702
R93 plus plus.n13 33.1808
R94 plus.n2 plus.n1 25.5611
R95 plus.n5 plus.n4 25.5611
R96 plus.n12 plus.n11 25.5611
R97 plus.n9 plus.n8 25.5611
R98 plus plus.n6 17.1482
R99 plus.n6 plus.n0 0.189894
R100 plus.n13 plus.n7 0.189894
R101 drain_left.n5 drain_left.n3 59.2758
R102 drain_left.n2 drain_left.n1 58.9403
R103 drain_left.n2 drain_left.n0 58.9403
R104 drain_left.n5 drain_left.n4 58.7153
R105 drain_left drain_left.n2 39.1768
R106 drain_left drain_left.n5 6.21356
R107 drain_left.n1 drain_left.t2 1.2005
R108 drain_left.n1 drain_left.t5 1.2005
R109 drain_left.n0 drain_left.t6 1.2005
R110 drain_left.n0 drain_left.t7 1.2005
R111 drain_left.n4 drain_left.t1 1.2005
R112 drain_left.n4 drain_left.t3 1.2005
R113 drain_left.n3 drain_left.t4 1.2005
R114 drain_left.n3 drain_left.t0 1.2005
C0 drain_right source 33.196102f
C1 drain_right plus 0.282599f
C2 drain_right minus 4.15789f
C3 source drain_left 33.1968f
C4 drain_left plus 4.28729f
C5 drain_left minus 0.170499f
C6 source plus 2.99088f
C7 source minus 2.97684f
C8 minus plus 7.24248f
C9 drain_right drain_left 0.640281f
C10 drain_right a_n1366_n5888# 7.77925f
C11 drain_left a_n1366_n5888# 7.97342f
C12 source a_n1366_n5888# 15.66515f
C13 minus a_n1366_n5888# 5.87051f
C14 plus a_n1366_n5888# 9.13688f
C15 drain_left.t6 a_n1366_n5888# 0.847269f
C16 drain_left.t7 a_n1366_n5888# 0.847269f
C17 drain_left.n0 a_n1366_n5888# 5.73099f
C18 drain_left.t2 a_n1366_n5888# 0.847269f
C19 drain_left.t5 a_n1366_n5888# 0.847269f
C20 drain_left.n1 a_n1366_n5888# 5.73099f
C21 drain_left.n2 a_n1366_n5888# 2.82352f
C22 drain_left.t4 a_n1366_n5888# 0.847269f
C23 drain_left.t0 a_n1366_n5888# 0.847269f
C24 drain_left.n3 a_n1366_n5888# 5.73309f
C25 drain_left.t1 a_n1366_n5888# 0.847269f
C26 drain_left.t3 a_n1366_n5888# 0.847269f
C27 drain_left.n4 a_n1366_n5888# 5.729741f
C28 drain_left.n5 a_n1366_n5888# 0.927414f
C29 plus.n0 a_n1366_n5888# 0.146883f
C30 plus.t6 a_n1366_n5888# 0.65439f
C31 plus.t7 a_n1366_n5888# 0.65439f
C32 plus.t3 a_n1366_n5888# 0.658468f
C33 plus.n1 a_n1366_n5888# 0.274788f
C34 plus.n2 a_n1366_n5888# 0.247677f
C35 plus.n3 a_n1366_n5888# 0.02631f
C36 plus.n4 a_n1366_n5888# 0.247677f
C37 plus.t4 a_n1366_n5888# 0.658468f
C38 plus.n5 a_n1366_n5888# 0.274689f
C39 plus.n6 a_n1366_n5888# 1.11825f
C40 plus.n7 a_n1366_n5888# 0.146883f
C41 plus.t1 a_n1366_n5888# 0.658468f
C42 plus.t0 a_n1366_n5888# 0.65439f
C43 plus.t5 a_n1366_n5888# 0.65439f
C44 plus.t2 a_n1366_n5888# 0.658468f
C45 plus.n8 a_n1366_n5888# 0.274788f
C46 plus.n9 a_n1366_n5888# 0.247677f
C47 plus.n10 a_n1366_n5888# 0.02631f
C48 plus.n11 a_n1366_n5888# 0.247677f
C49 plus.n12 a_n1366_n5888# 0.274689f
C50 plus.n13 a_n1366_n5888# 2.2525f
C51 drain_right.t6 a_n1366_n5888# 0.847512f
C52 drain_right.t1 a_n1366_n5888# 0.847512f
C53 drain_right.n0 a_n1366_n5888# 5.73264f
C54 drain_right.t0 a_n1366_n5888# 0.847512f
C55 drain_right.t7 a_n1366_n5888# 0.847512f
C56 drain_right.n1 a_n1366_n5888# 5.73264f
C57 drain_right.n2 a_n1366_n5888# 2.76525f
C58 drain_right.t5 a_n1366_n5888# 0.847512f
C59 drain_right.t4 a_n1366_n5888# 0.847512f
C60 drain_right.n3 a_n1366_n5888# 5.73472f
C61 drain_right.t3 a_n1366_n5888# 0.847512f
C62 drain_right.t2 a_n1366_n5888# 0.847512f
C63 drain_right.n4 a_n1366_n5888# 5.7314f
C64 drain_right.n5 a_n1366_n5888# 0.92768f
C65 source.t4 a_n1366_n5888# 4.96343f
C66 source.n0 a_n1366_n5888# 1.89925f
C67 source.t3 a_n1366_n5888# 0.601905f
C68 source.t5 a_n1366_n5888# 0.601905f
C69 source.n1 a_n1366_n5888# 4.00453f
C70 source.n2 a_n1366_n5888# 0.281178f
C71 source.t0 a_n1366_n5888# 4.96345f
C72 source.n3 a_n1366_n5888# 0.399821f
C73 source.t9 a_n1366_n5888# 4.96345f
C74 source.n4 a_n1366_n5888# 0.399821f
C75 source.t7 a_n1366_n5888# 0.601905f
C76 source.t12 a_n1366_n5888# 0.601905f
C77 source.n5 a_n1366_n5888# 4.00453f
C78 source.n6 a_n1366_n5888# 0.281178f
C79 source.t8 a_n1366_n5888# 4.96345f
C80 source.n7 a_n1366_n5888# 2.27173f
C81 source.t15 a_n1366_n5888# 4.96343f
C82 source.n8 a_n1366_n5888# 2.27175f
C83 source.t14 a_n1366_n5888# 0.601905f
C84 source.t2 a_n1366_n5888# 0.601905f
C85 source.n9 a_n1366_n5888# 4.00453f
C86 source.n10 a_n1366_n5888# 0.281179f
C87 source.t1 a_n1366_n5888# 4.96343f
C88 source.n11 a_n1366_n5888# 0.399834f
C89 source.t10 a_n1366_n5888# 4.96343f
C90 source.n12 a_n1366_n5888# 0.399834f
C91 source.t11 a_n1366_n5888# 0.601905f
C92 source.t6 a_n1366_n5888# 0.601905f
C93 source.n13 a_n1366_n5888# 4.00453f
C94 source.n14 a_n1366_n5888# 0.281179f
C95 source.t13 a_n1366_n5888# 4.96343f
C96 source.n15 a_n1366_n5888# 0.514239f
C97 source.n16 a_n1366_n5888# 2.14432f
C98 minus.n0 a_n1366_n5888# 0.144619f
C99 minus.t4 a_n1366_n5888# 0.648319f
C100 minus.t5 a_n1366_n5888# 0.644304f
C101 minus.t2 a_n1366_n5888# 0.644304f
C102 minus.t3 a_n1366_n5888# 0.648319f
C103 minus.n1 a_n1366_n5888# 0.270553f
C104 minus.n2 a_n1366_n5888# 0.24386f
C105 minus.n3 a_n1366_n5888# 0.025904f
C106 minus.n4 a_n1366_n5888# 0.24386f
C107 minus.n5 a_n1366_n5888# 0.270455f
C108 minus.n6 a_n1366_n5888# 2.91877f
C109 minus.n7 a_n1366_n5888# 0.144619f
C110 minus.t7 a_n1366_n5888# 0.644304f
C111 minus.t6 a_n1366_n5888# 0.644304f
C112 minus.t1 a_n1366_n5888# 0.648319f
C113 minus.n8 a_n1366_n5888# 0.270553f
C114 minus.n9 a_n1366_n5888# 0.24386f
C115 minus.n10 a_n1366_n5888# 0.025904f
C116 minus.n11 a_n1366_n5888# 0.24386f
C117 minus.t0 a_n1366_n5888# 0.648319f
C118 minus.n12 a_n1366_n5888# 0.270455f
C119 minus.n13 a_n1366_n5888# 0.410692f
C120 minus.n14 a_n1366_n5888# 3.46145f
.ends

