* NGSPICE file created from diffpair504.ext - technology: sky130A

.subckt diffpair504 minus drain_right drain_left source plus
X0 source.t15 plus.t0 drain_left.t9 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X1 source.t14 plus.t1 drain_left.t3 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X2 drain_left.t2 plus.t2 source.t13 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X3 source.t0 minus.t0 drain_right.t9 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X4 source.t4 minus.t1 drain_right.t8 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X5 drain_right.t7 minus.t2 source.t17 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X6 source.t12 plus.t3 drain_left.t5 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X7 drain_left.t1 plus.t4 source.t11 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X8 a_n1412_n3888# a_n1412_n3888# a_n1412_n3888# a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.25
X9 source.t18 minus.t3 drain_right.t6 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X10 drain_left.t4 plus.t5 source.t10 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X11 drain_right.t5 minus.t4 source.t19 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X12 drain_left.t6 plus.t6 source.t9 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X13 drain_left.t7 plus.t7 source.t8 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X14 a_n1412_n3888# a_n1412_n3888# a_n1412_n3888# a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X15 drain_left.t8 plus.t8 source.t7 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X16 drain_right.t4 minus.t5 source.t3 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X17 drain_right.t3 minus.t6 source.t2 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.25
X18 source.t5 minus.t7 drain_right.t2 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X19 drain_right.t1 minus.t8 source.t1 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.25
X20 a_n1412_n3888# a_n1412_n3888# a_n1412_n3888# a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X21 source.t6 plus.t9 drain_left.t0 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
X22 a_n1412_n3888# a_n1412_n3888# a_n1412_n3888# a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.25
X23 drain_right.t0 minus.t9 source.t16 a_n1412_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.25
R0 plus.n2 plus.t4 1631.2
R1 plus.n8 plus.t6 1631.2
R2 plus.n12 plus.t2 1631.2
R3 plus.n18 plus.t5 1631.2
R4 plus.n1 plus.t1 1571.32
R5 plus.n5 plus.t7 1571.32
R6 plus.n7 plus.t0 1571.32
R7 plus.n11 plus.t9 1571.32
R8 plus.n15 plus.t8 1571.32
R9 plus.n17 plus.t3 1571.32
R10 plus.n3 plus.n2 161.489
R11 plus.n13 plus.n12 161.489
R12 plus.n4 plus.n3 161.3
R13 plus.n6 plus.n0 161.3
R14 plus.n9 plus.n8 161.3
R15 plus.n14 plus.n13 161.3
R16 plus.n16 plus.n10 161.3
R17 plus.n19 plus.n18 161.3
R18 plus.n4 plus.n1 48.2005
R19 plus.n7 plus.n6 48.2005
R20 plus.n17 plus.n16 48.2005
R21 plus.n14 plus.n11 48.2005
R22 plus.n5 plus.n4 36.5157
R23 plus.n6 plus.n5 36.5157
R24 plus.n16 plus.n15 36.5157
R25 plus.n15 plus.n14 36.5157
R26 plus plus.n19 29.5028
R27 plus.n2 plus.n1 24.8308
R28 plus.n8 plus.n7 24.8308
R29 plus.n18 plus.n17 24.8308
R30 plus.n12 plus.n11 24.8308
R31 plus plus.n9 13.296
R32 plus.n3 plus.n0 0.189894
R33 plus.n9 plus.n0 0.189894
R34 plus.n19 plus.n10 0.189894
R35 plus.n13 plus.n10 0.189894
R36 drain_left.n5 drain_left.t1 62.6998
R37 drain_left.n1 drain_left.t4 62.6996
R38 drain_left.n3 drain_left.n2 61.1992
R39 drain_left.n5 drain_left.n4 60.8798
R40 drain_left.n7 drain_left.n6 60.8796
R41 drain_left.n1 drain_left.n0 60.8796
R42 drain_left drain_left.n3 31.7648
R43 drain_left drain_left.n7 6.15322
R44 drain_left.n2 drain_left.t0 1.3205
R45 drain_left.n2 drain_left.t2 1.3205
R46 drain_left.n0 drain_left.t5 1.3205
R47 drain_left.n0 drain_left.t8 1.3205
R48 drain_left.n6 drain_left.t9 1.3205
R49 drain_left.n6 drain_left.t6 1.3205
R50 drain_left.n4 drain_left.t3 1.3205
R51 drain_left.n4 drain_left.t7 1.3205
R52 drain_left.n7 drain_left.n5 0.5005
R53 drain_left.n3 drain_left.n1 0.070154
R54 source.n5 source.t2 45.521
R55 source.n19 source.t19 45.5208
R56 source.n14 source.t13 45.5208
R57 source.n0 source.t9 45.5208
R58 source.n2 source.n1 44.201
R59 source.n4 source.n3 44.201
R60 source.n7 source.n6 44.201
R61 source.n9 source.n8 44.201
R62 source.n18 source.n17 44.2008
R63 source.n16 source.n15 44.2008
R64 source.n13 source.n12 44.2008
R65 source.n11 source.n10 44.2008
R66 source.n11 source.n9 24.5605
R67 source.n20 source.n0 18.5475
R68 source.n20 source.n19 5.51343
R69 source.n17 source.t16 1.3205
R70 source.n17 source.t5 1.3205
R71 source.n15 source.t17 1.3205
R72 source.n15 source.t18 1.3205
R73 source.n12 source.t7 1.3205
R74 source.n12 source.t6 1.3205
R75 source.n10 source.t10 1.3205
R76 source.n10 source.t12 1.3205
R77 source.n1 source.t8 1.3205
R78 source.n1 source.t15 1.3205
R79 source.n3 source.t11 1.3205
R80 source.n3 source.t14 1.3205
R81 source.n6 source.t3 1.3205
R82 source.n6 source.t4 1.3205
R83 source.n8 source.t1 1.3205
R84 source.n8 source.t0 1.3205
R85 source.n5 source.n4 0.720328
R86 source.n16 source.n14 0.720328
R87 source.n9 source.n7 0.5005
R88 source.n7 source.n5 0.5005
R89 source.n4 source.n2 0.5005
R90 source.n2 source.n0 0.5005
R91 source.n13 source.n11 0.5005
R92 source.n14 source.n13 0.5005
R93 source.n18 source.n16 0.5005
R94 source.n19 source.n18 0.5005
R95 source source.n20 0.188
R96 minus.n8 minus.t8 1631.2
R97 minus.n2 minus.t6 1631.2
R98 minus.n18 minus.t4 1631.2
R99 minus.n12 minus.t2 1631.2
R100 minus.n7 minus.t0 1571.32
R101 minus.n5 minus.t5 1571.32
R102 minus.n1 minus.t1 1571.32
R103 minus.n17 minus.t7 1571.32
R104 minus.n15 minus.t9 1571.32
R105 minus.n11 minus.t3 1571.32
R106 minus.n3 minus.n2 161.489
R107 minus.n13 minus.n12 161.489
R108 minus.n9 minus.n8 161.3
R109 minus.n6 minus.n0 161.3
R110 minus.n4 minus.n3 161.3
R111 minus.n19 minus.n18 161.3
R112 minus.n16 minus.n10 161.3
R113 minus.n14 minus.n13 161.3
R114 minus.n7 minus.n6 48.2005
R115 minus.n4 minus.n1 48.2005
R116 minus.n14 minus.n11 48.2005
R117 minus.n17 minus.n16 48.2005
R118 minus.n20 minus.n9 36.7581
R119 minus.n6 minus.n5 36.5157
R120 minus.n5 minus.n4 36.5157
R121 minus.n15 minus.n14 36.5157
R122 minus.n16 minus.n15 36.5157
R123 minus.n8 minus.n7 24.8308
R124 minus.n2 minus.n1 24.8308
R125 minus.n12 minus.n11 24.8308
R126 minus.n18 minus.n17 24.8308
R127 minus.n20 minus.n19 6.51565
R128 minus.n9 minus.n0 0.189894
R129 minus.n3 minus.n0 0.189894
R130 minus.n13 minus.n10 0.189894
R131 minus.n19 minus.n10 0.189894
R132 minus minus.n20 0.188
R133 drain_right.n1 drain_right.t7 62.6996
R134 drain_right.n7 drain_right.t1 62.1998
R135 drain_right.n6 drain_right.n4 61.3796
R136 drain_right.n3 drain_right.n2 61.1992
R137 drain_right.n6 drain_right.n5 60.8798
R138 drain_right.n1 drain_right.n0 60.8796
R139 drain_right drain_right.n3 31.2116
R140 drain_right drain_right.n7 5.90322
R141 drain_right.n2 drain_right.t2 1.3205
R142 drain_right.n2 drain_right.t5 1.3205
R143 drain_right.n0 drain_right.t6 1.3205
R144 drain_right.n0 drain_right.t0 1.3205
R145 drain_right.n4 drain_right.t8 1.3205
R146 drain_right.n4 drain_right.t3 1.3205
R147 drain_right.n5 drain_right.t9 1.3205
R148 drain_right.n5 drain_right.t4 1.3205
R149 drain_right.n7 drain_right.n6 0.5005
R150 drain_right.n3 drain_right.n1 0.070154
C0 drain_right plus 0.290745f
C1 drain_left drain_right 0.695203f
C2 minus source 3.77831f
C3 plus minus 5.46562f
C4 plus source 3.7932f
C5 drain_left minus 0.171039f
C6 drain_right minus 4.34033f
C7 drain_left source 27.9289f
C8 drain_right source 27.9147f
C9 drain_left plus 4.47088f
C10 drain_right a_n1412_n3888# 7.88277f
C11 drain_left a_n1412_n3888# 8.126981f
C12 source a_n1412_n3888# 7.070911f
C13 minus a_n1412_n3888# 5.642716f
C14 plus a_n1412_n3888# 7.91656f
C15 drain_right.t7 a_n1412_n3888# 4.28396f
C16 drain_right.t6 a_n1412_n3888# 0.371024f
C17 drain_right.t0 a_n1412_n3888# 0.371024f
C18 drain_right.n0 a_n1412_n3888# 3.35362f
C19 drain_right.n1 a_n1412_n3888# 0.725204f
C20 drain_right.t2 a_n1412_n3888# 0.371024f
C21 drain_right.t5 a_n1412_n3888# 0.371024f
C22 drain_right.n2 a_n1412_n3888# 3.35547f
C23 drain_right.n3 a_n1412_n3888# 1.89182f
C24 drain_right.t8 a_n1412_n3888# 0.371024f
C25 drain_right.t3 a_n1412_n3888# 0.371024f
C26 drain_right.n4 a_n1412_n3888# 3.35662f
C27 drain_right.t9 a_n1412_n3888# 0.371024f
C28 drain_right.t4 a_n1412_n3888# 0.371024f
C29 drain_right.n5 a_n1412_n3888# 3.35362f
C30 drain_right.n6 a_n1412_n3888# 0.724064f
C31 drain_right.t1 a_n1412_n3888# 4.28073f
C32 drain_right.n7 a_n1412_n3888# 0.661949f
C33 minus.n0 a_n1412_n3888# 0.055637f
C34 minus.t8 a_n1412_n3888# 0.597209f
C35 minus.t0 a_n1412_n3888# 0.588602f
C36 minus.t5 a_n1412_n3888# 0.588602f
C37 minus.t1 a_n1412_n3888# 0.588602f
C38 minus.n1 a_n1412_n3888# 0.228944f
C39 minus.t6 a_n1412_n3888# 0.597209f
C40 minus.n2 a_n1412_n3888# 0.247115f
C41 minus.n3 a_n1412_n3888# 0.130738f
C42 minus.n4 a_n1412_n3888# 0.021201f
C43 minus.n5 a_n1412_n3888# 0.228944f
C44 minus.n6 a_n1412_n3888# 0.021201f
C45 minus.n7 a_n1412_n3888# 0.228944f
C46 minus.n8 a_n1412_n3888# 0.247027f
C47 minus.n9 a_n1412_n3888# 2.01492f
C48 minus.n10 a_n1412_n3888# 0.055637f
C49 minus.t7 a_n1412_n3888# 0.588602f
C50 minus.t9 a_n1412_n3888# 0.588602f
C51 minus.t3 a_n1412_n3888# 0.588602f
C52 minus.n11 a_n1412_n3888# 0.228944f
C53 minus.t2 a_n1412_n3888# 0.597209f
C54 minus.n12 a_n1412_n3888# 0.247115f
C55 minus.n13 a_n1412_n3888# 0.130738f
C56 minus.n14 a_n1412_n3888# 0.021201f
C57 minus.n15 a_n1412_n3888# 0.228944f
C58 minus.n16 a_n1412_n3888# 0.021201f
C59 minus.n17 a_n1412_n3888# 0.228944f
C60 minus.t4 a_n1412_n3888# 0.597209f
C61 minus.n18 a_n1412_n3888# 0.247027f
C62 minus.n19 a_n1412_n3888# 0.365791f
C63 minus.n20 a_n1412_n3888# 2.44281f
C64 source.t9 a_n1412_n3888# 4.25666f
C65 source.n0 a_n1412_n3888# 1.96442f
C66 source.t8 a_n1412_n3888# 0.379835f
C67 source.t15 a_n1412_n3888# 0.379835f
C68 source.n1 a_n1412_n3888# 3.33653f
C69 source.n2 a_n1412_n3888# 0.418893f
C70 source.t11 a_n1412_n3888# 0.379835f
C71 source.t14 a_n1412_n3888# 0.379835f
C72 source.n3 a_n1412_n3888# 3.33653f
C73 source.n4 a_n1412_n3888# 0.441591f
C74 source.t2 a_n1412_n3888# 4.25666f
C75 source.n5 a_n1412_n3888# 0.557368f
C76 source.t3 a_n1412_n3888# 0.379835f
C77 source.t4 a_n1412_n3888# 0.379835f
C78 source.n6 a_n1412_n3888# 3.33653f
C79 source.n7 a_n1412_n3888# 0.418893f
C80 source.t1 a_n1412_n3888# 0.379835f
C81 source.t0 a_n1412_n3888# 0.379835f
C82 source.n8 a_n1412_n3888# 3.33653f
C83 source.n9 a_n1412_n3888# 2.43131f
C84 source.t10 a_n1412_n3888# 0.379835f
C85 source.t12 a_n1412_n3888# 0.379835f
C86 source.n10 a_n1412_n3888# 3.33652f
C87 source.n11 a_n1412_n3888# 2.43131f
C88 source.t7 a_n1412_n3888# 0.379835f
C89 source.t6 a_n1412_n3888# 0.379835f
C90 source.n12 a_n1412_n3888# 3.33652f
C91 source.n13 a_n1412_n3888# 0.418897f
C92 source.t13 a_n1412_n3888# 4.25666f
C93 source.n14 a_n1412_n3888# 0.557373f
C94 source.t17 a_n1412_n3888# 0.379835f
C95 source.t18 a_n1412_n3888# 0.379835f
C96 source.n15 a_n1412_n3888# 3.33652f
C97 source.n16 a_n1412_n3888# 0.441595f
C98 source.t16 a_n1412_n3888# 0.379835f
C99 source.t5 a_n1412_n3888# 0.379835f
C100 source.n17 a_n1412_n3888# 3.33652f
C101 source.n18 a_n1412_n3888# 0.418897f
C102 source.t19 a_n1412_n3888# 4.25666f
C103 source.n19 a_n1412_n3888# 0.708887f
C104 source.n20 a_n1412_n3888# 2.34042f
C105 drain_left.t4 a_n1412_n3888# 4.29423f
C106 drain_left.t5 a_n1412_n3888# 0.371914f
C107 drain_left.t8 a_n1412_n3888# 0.371914f
C108 drain_left.n0 a_n1412_n3888# 3.36167f
C109 drain_left.n1 a_n1412_n3888# 0.726944f
C110 drain_left.t0 a_n1412_n3888# 0.371914f
C111 drain_left.t2 a_n1412_n3888# 0.371914f
C112 drain_left.n2 a_n1412_n3888# 3.36352f
C113 drain_left.n3 a_n1412_n3888# 1.96216f
C114 drain_left.t1 a_n1412_n3888# 4.29424f
C115 drain_left.t3 a_n1412_n3888# 0.371914f
C116 drain_left.t7 a_n1412_n3888# 0.371914f
C117 drain_left.n4 a_n1412_n3888# 3.36167f
C118 drain_left.n5 a_n1412_n3888# 0.760003f
C119 drain_left.t9 a_n1412_n3888# 0.371914f
C120 drain_left.t6 a_n1412_n3888# 0.371914f
C121 drain_left.n6 a_n1412_n3888# 3.36166f
C122 drain_left.n7 a_n1412_n3888# 0.617086f
C123 plus.n0 a_n1412_n3888# 0.056926f
C124 plus.t0 a_n1412_n3888# 0.60224f
C125 plus.t7 a_n1412_n3888# 0.60224f
C126 plus.t1 a_n1412_n3888# 0.60224f
C127 plus.n1 a_n1412_n3888# 0.234249f
C128 plus.t4 a_n1412_n3888# 0.611046f
C129 plus.n2 a_n1412_n3888# 0.252841f
C130 plus.n3 a_n1412_n3888# 0.133768f
C131 plus.n4 a_n1412_n3888# 0.021692f
C132 plus.n5 a_n1412_n3888# 0.234249f
C133 plus.n6 a_n1412_n3888# 0.021692f
C134 plus.n7 a_n1412_n3888# 0.234249f
C135 plus.t6 a_n1412_n3888# 0.611046f
C136 plus.n8 a_n1412_n3888# 0.252751f
C137 plus.n9 a_n1412_n3888# 0.721465f
C138 plus.n10 a_n1412_n3888# 0.056926f
C139 plus.t5 a_n1412_n3888# 0.611046f
C140 plus.t3 a_n1412_n3888# 0.60224f
C141 plus.t8 a_n1412_n3888# 0.60224f
C142 plus.t9 a_n1412_n3888# 0.60224f
C143 plus.n11 a_n1412_n3888# 0.234249f
C144 plus.t2 a_n1412_n3888# 0.611046f
C145 plus.n12 a_n1412_n3888# 0.252841f
C146 plus.n13 a_n1412_n3888# 0.133768f
C147 plus.n14 a_n1412_n3888# 0.021692f
C148 plus.n15 a_n1412_n3888# 0.234249f
C149 plus.n16 a_n1412_n3888# 0.021692f
C150 plus.n17 a_n1412_n3888# 0.234249f
C151 plus.n18 a_n1412_n3888# 0.252751f
C152 plus.n19 a_n1412_n3888# 1.68891f
.ends

