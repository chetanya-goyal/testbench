* NGSPICE file created from diffpair373.ext - technology: sky130A

.subckt diffpair373 minus drain_right drain_left source plus
X0 a_n1646_n2688# a_n1646_n2688# a_n1646_n2688# a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.6
X1 a_n1646_n2688# a_n1646_n2688# a_n1646_n2688# a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X2 source.t15 minus.t0 drain_right.t7 a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X3 source.t1 plus.t0 drain_left.t7 a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X4 source.t14 minus.t1 drain_right.t2 a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X5 drain_left.t6 plus.t1 source.t3 a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X6 source.t13 minus.t2 drain_right.t4 a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X7 drain_right.t0 minus.t3 source.t12 a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X8 drain_left.t5 plus.t2 source.t0 a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X9 source.t11 minus.t4 drain_right.t3 a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X10 source.t7 plus.t3 drain_left.t4 a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X11 drain_right.t1 minus.t5 source.t10 a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X12 drain_left.t3 plus.t4 source.t6 a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X13 source.t5 plus.t5 drain_left.t2 a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X14 drain_right.t5 minus.t6 source.t9 a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X15 drain_left.t1 plus.t6 source.t2 a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X16 source.t4 plus.t7 drain_left.t0 a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X17 a_n1646_n2688# a_n1646_n2688# a_n1646_n2688# a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X18 drain_right.t6 minus.t7 source.t8 a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X19 a_n1646_n2688# a_n1646_n2688# a_n1646_n2688# a_n1646_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
R0 minus.n1 minus.t5 453.793
R1 minus.n7 minus.t1 453.793
R2 minus.n2 minus.t4 426.973
R3 minus.n3 minus.t3 426.973
R4 minus.n4 minus.t2 426.973
R5 minus.n8 minus.t7 426.973
R6 minus.n9 minus.t0 426.973
R7 minus.n10 minus.t6 426.973
R8 minus.n5 minus.n4 161.3
R9 minus.n11 minus.n10 161.3
R10 minus.n3 minus.n0 80.6037
R11 minus.n9 minus.n6 80.6037
R12 minus.n3 minus.n2 48.2005
R13 minus.n4 minus.n3 48.2005
R14 minus.n9 minus.n8 48.2005
R15 minus.n10 minus.n9 48.2005
R16 minus.n1 minus.n0 45.2318
R17 minus.n7 minus.n6 45.2318
R18 minus.n12 minus.n5 33.1975
R19 minus.n2 minus.n1 13.3799
R20 minus.n8 minus.n7 13.3799
R21 minus.n12 minus.n11 6.61414
R22 minus.n5 minus.n0 0.285035
R23 minus.n11 minus.n6 0.285035
R24 minus minus.n12 0.188
R25 drain_right.n5 drain_right.n3 66.3391
R26 drain_right.n2 drain_right.n1 65.8829
R27 drain_right.n2 drain_right.n0 65.8829
R28 drain_right.n5 drain_right.n4 65.5376
R29 drain_right drain_right.n2 27.3472
R30 drain_right drain_right.n5 6.45494
R31 drain_right.n1 drain_right.t7 2.2005
R32 drain_right.n1 drain_right.t5 2.2005
R33 drain_right.n0 drain_right.t2 2.2005
R34 drain_right.n0 drain_right.t6 2.2005
R35 drain_right.n3 drain_right.t3 2.2005
R36 drain_right.n3 drain_right.t1 2.2005
R37 drain_right.n4 drain_right.t4 2.2005
R38 drain_right.n4 drain_right.t0 2.2005
R39 source.n3 source.t5 51.0588
R40 source.n4 source.t10 51.0588
R41 source.n7 source.t13 51.0588
R42 source.n15 source.t9 51.0586
R43 source.n12 source.t14 51.0586
R44 source.n11 source.t2 51.0586
R45 source.n8 source.t4 51.0586
R46 source.n0 source.t0 51.0586
R47 source.n2 source.n1 48.8588
R48 source.n6 source.n5 48.8588
R49 source.n14 source.n13 48.8586
R50 source.n10 source.n9 48.8586
R51 source.n8 source.n7 19.8167
R52 source.n16 source.n0 14.1529
R53 source.n16 source.n15 5.66429
R54 source.n13 source.t8 2.2005
R55 source.n13 source.t15 2.2005
R56 source.n9 source.t3 2.2005
R57 source.n9 source.t1 2.2005
R58 source.n1 source.t6 2.2005
R59 source.n1 source.t7 2.2005
R60 source.n5 source.t12 2.2005
R61 source.n5 source.t11 2.2005
R62 source.n7 source.n6 0.802224
R63 source.n6 source.n4 0.802224
R64 source.n3 source.n2 0.802224
R65 source.n2 source.n0 0.802224
R66 source.n10 source.n8 0.802224
R67 source.n11 source.n10 0.802224
R68 source.n14 source.n12 0.802224
R69 source.n15 source.n14 0.802224
R70 source.n4 source.n3 0.470328
R71 source.n12 source.n11 0.470328
R72 source source.n16 0.188
R73 plus.n1 plus.t5 453.793
R74 plus.n7 plus.t6 453.793
R75 plus.n4 plus.t2 426.973
R76 plus.n3 plus.t3 426.973
R77 plus.n2 plus.t4 426.973
R78 plus.n10 plus.t7 426.973
R79 plus.n9 plus.t1 426.973
R80 plus.n8 plus.t0 426.973
R81 plus.n5 plus.n4 161.3
R82 plus.n11 plus.n10 161.3
R83 plus.n3 plus.n0 80.6037
R84 plus.n9 plus.n6 80.6037
R85 plus.n4 plus.n3 48.2005
R86 plus.n3 plus.n2 48.2005
R87 plus.n10 plus.n9 48.2005
R88 plus.n9 plus.n8 48.2005
R89 plus.n1 plus.n0 45.2318
R90 plus.n7 plus.n6 45.2318
R91 plus plus.n11 28.2149
R92 plus.n2 plus.n1 13.3799
R93 plus.n8 plus.n7 13.3799
R94 plus plus.n5 11.1217
R95 plus.n5 plus.n0 0.285035
R96 plus.n11 plus.n6 0.285035
R97 drain_left.n5 drain_left.n3 66.3393
R98 drain_left.n2 drain_left.n1 65.8829
R99 drain_left.n2 drain_left.n0 65.8829
R100 drain_left.n5 drain_left.n4 65.5374
R101 drain_left drain_left.n2 27.9004
R102 drain_left drain_left.n5 6.45494
R103 drain_left.n1 drain_left.t7 2.2005
R104 drain_left.n1 drain_left.t1 2.2005
R105 drain_left.n0 drain_left.t0 2.2005
R106 drain_left.n0 drain_left.t6 2.2005
R107 drain_left.n4 drain_left.t4 2.2005
R108 drain_left.n4 drain_left.t5 2.2005
R109 drain_left.n3 drain_left.t2 2.2005
R110 drain_left.n3 drain_left.t3 2.2005
C0 drain_right plus 0.312845f
C1 source drain_left 9.543f
C2 drain_right source 9.54415f
C3 source plus 3.75445f
C4 minus drain_left 0.171399f
C5 drain_right minus 3.90667f
C6 minus plus 4.63999f
C7 drain_right drain_left 0.775958f
C8 plus drain_left 4.0651f
C9 source minus 3.74041f
C10 drain_right a_n1646_n2688# 5.03732f
C11 drain_left a_n1646_n2688# 5.29179f
C12 source a_n1646_n2688# 7.178778f
C13 minus a_n1646_n2688# 6.15536f
C14 plus a_n1646_n2688# 7.74815f
C15 drain_left.t0 a_n1646_n2688# 0.19703f
C16 drain_left.t6 a_n1646_n2688# 0.19703f
C17 drain_left.n0 a_n1646_n2688# 1.72512f
C18 drain_left.t7 a_n1646_n2688# 0.19703f
C19 drain_left.t1 a_n1646_n2688# 0.19703f
C20 drain_left.n1 a_n1646_n2688# 1.72512f
C21 drain_left.n2 a_n1646_n2688# 1.8032f
C22 drain_left.t2 a_n1646_n2688# 0.19703f
C23 drain_left.t3 a_n1646_n2688# 0.19703f
C24 drain_left.n3 a_n1646_n2688# 1.7279f
C25 drain_left.t4 a_n1646_n2688# 0.19703f
C26 drain_left.t5 a_n1646_n2688# 0.19703f
C27 drain_left.n4 a_n1646_n2688# 1.72335f
C28 drain_left.n5 a_n1646_n2688# 0.978271f
C29 plus.n0 a_n1646_n2688# 0.232836f
C30 plus.t2 a_n1646_n2688# 0.73948f
C31 plus.t3 a_n1646_n2688# 0.73948f
C32 plus.t4 a_n1646_n2688# 0.73948f
C33 plus.t5 a_n1646_n2688# 0.757987f
C34 plus.n1 a_n1646_n2688# 0.29592f
C35 plus.n2 a_n1646_n2688# 0.323833f
C36 plus.n3 a_n1646_n2688# 0.323833f
C37 plus.n4 a_n1646_n2688# 0.312997f
C38 plus.n5 a_n1646_n2688# 0.498191f
C39 plus.n6 a_n1646_n2688# 0.232836f
C40 plus.t7 a_n1646_n2688# 0.73948f
C41 plus.t1 a_n1646_n2688# 0.73948f
C42 plus.t6 a_n1646_n2688# 0.757987f
C43 plus.n7 a_n1646_n2688# 0.29592f
C44 plus.t0 a_n1646_n2688# 0.73948f
C45 plus.n8 a_n1646_n2688# 0.323833f
C46 plus.n9 a_n1646_n2688# 0.323833f
C47 plus.n10 a_n1646_n2688# 0.312997f
C48 plus.n11 a_n1646_n2688# 1.30284f
C49 source.t0 a_n1646_n2688# 1.58575f
C50 source.n0 a_n1646_n2688# 0.940992f
C51 source.t6 a_n1646_n2688# 0.148709f
C52 source.t7 a_n1646_n2688# 0.148709f
C53 source.n1 a_n1646_n2688# 1.24489f
C54 source.n2 a_n1646_n2688# 0.30291f
C55 source.t5 a_n1646_n2688# 1.58575f
C56 source.n3 a_n1646_n2688# 0.345256f
C57 source.t10 a_n1646_n2688# 1.58575f
C58 source.n4 a_n1646_n2688# 0.345256f
C59 source.t12 a_n1646_n2688# 0.148709f
C60 source.t11 a_n1646_n2688# 0.148709f
C61 source.n5 a_n1646_n2688# 1.24489f
C62 source.n6 a_n1646_n2688# 0.30291f
C63 source.t13 a_n1646_n2688# 1.58575f
C64 source.n7 a_n1646_n2688# 1.25051f
C65 source.t4 a_n1646_n2688# 1.58575f
C66 source.n8 a_n1646_n2688# 1.25051f
C67 source.t3 a_n1646_n2688# 0.148709f
C68 source.t1 a_n1646_n2688# 0.148709f
C69 source.n9 a_n1646_n2688# 1.24489f
C70 source.n10 a_n1646_n2688# 0.302914f
C71 source.t2 a_n1646_n2688# 1.58575f
C72 source.n11 a_n1646_n2688# 0.34526f
C73 source.t14 a_n1646_n2688# 1.58575f
C74 source.n12 a_n1646_n2688# 0.34526f
C75 source.t8 a_n1646_n2688# 0.148709f
C76 source.t15 a_n1646_n2688# 0.148709f
C77 source.n13 a_n1646_n2688# 1.24489f
C78 source.n14 a_n1646_n2688# 0.302914f
C79 source.t9 a_n1646_n2688# 1.58575f
C80 source.n15 a_n1646_n2688# 0.477101f
C81 source.n16 a_n1646_n2688# 1.0978f
C82 drain_right.t2 a_n1646_n2688# 0.195691f
C83 drain_right.t6 a_n1646_n2688# 0.195691f
C84 drain_right.n0 a_n1646_n2688# 1.7134f
C85 drain_right.t7 a_n1646_n2688# 0.195691f
C86 drain_right.t5 a_n1646_n2688# 0.195691f
C87 drain_right.n1 a_n1646_n2688# 1.7134f
C88 drain_right.n2 a_n1646_n2688# 1.73409f
C89 drain_right.t3 a_n1646_n2688# 0.195691f
C90 drain_right.t1 a_n1646_n2688# 0.195691f
C91 drain_right.n3 a_n1646_n2688# 1.71616f
C92 drain_right.t4 a_n1646_n2688# 0.195691f
C93 drain_right.t0 a_n1646_n2688# 0.195691f
C94 drain_right.n4 a_n1646_n2688# 1.71165f
C95 drain_right.n5 a_n1646_n2688# 0.971628f
C96 minus.n0 a_n1646_n2688# 0.225506f
C97 minus.t4 a_n1646_n2688# 0.7162f
C98 minus.t5 a_n1646_n2688# 0.734124f
C99 minus.n1 a_n1646_n2688# 0.286604f
C100 minus.n2 a_n1646_n2688# 0.313638f
C101 minus.t3 a_n1646_n2688# 0.7162f
C102 minus.n3 a_n1646_n2688# 0.313638f
C103 minus.t2 a_n1646_n2688# 0.7162f
C104 minus.n4 a_n1646_n2688# 0.303143f
C105 minus.n5 a_n1646_n2688# 1.44403f
C106 minus.n6 a_n1646_n2688# 0.225506f
C107 minus.t1 a_n1646_n2688# 0.734124f
C108 minus.n7 a_n1646_n2688# 0.286604f
C109 minus.t7 a_n1646_n2688# 0.7162f
C110 minus.n8 a_n1646_n2688# 0.313638f
C111 minus.t0 a_n1646_n2688# 0.7162f
C112 minus.n9 a_n1646_n2688# 0.313638f
C113 minus.t6 a_n1646_n2688# 0.7162f
C114 minus.n10 a_n1646_n2688# 0.303143f
C115 minus.n11 a_n1646_n2688# 0.330183f
C116 minus.n12 a_n1646_n2688# 1.74492f
.ends

