* NGSPICE file created from diffpair629.ext - technology: sky130A

.subckt diffpair629 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t25 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X1 a_n3394_n4888# a_n3394_n4888# a_n3394_n4888# a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.7
X2 source.t12 minus.t0 drain_right.t23 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X3 source.t33 plus.t1 drain_left.t22 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X4 drain_left.t21 plus.t2 source.t44 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X5 source.t42 plus.t3 drain_left.t20 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X6 drain_right.t22 minus.t1 source.t6 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X7 source.t29 plus.t4 drain_left.t19 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X8 source.t8 minus.t2 drain_right.t21 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X9 drain_left.t18 plus.t5 source.t28 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X10 source.t20 minus.t3 drain_right.t20 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X11 source.t19 minus.t4 drain_right.t19 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X12 source.t39 plus.t6 drain_left.t17 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X13 source.t40 plus.t7 drain_left.t16 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X14 drain_right.t18 minus.t5 source.t13 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X15 drain_right.t17 minus.t6 source.t2 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X16 source.t41 plus.t8 drain_left.t15 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X17 drain_left.t14 plus.t9 source.t43 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X18 drain_right.t16 minus.t7 source.t11 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X19 source.t14 minus.t8 drain_right.t15 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X20 drain_right.t14 minus.t9 source.t0 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X21 drain_right.t13 minus.t10 source.t18 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X22 drain_right.t12 minus.t11 source.t1 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X23 drain_right.t11 minus.t12 source.t10 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X24 drain_left.t13 plus.t10 source.t27 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X25 a_n3394_n4888# a_n3394_n4888# a_n3394_n4888# a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X26 drain_right.t10 minus.t13 source.t17 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X27 drain_left.t12 plus.t11 source.t26 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X28 source.t37 plus.t12 drain_left.t11 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X29 drain_left.t10 plus.t13 source.t36 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X30 source.t35 plus.t14 drain_left.t9 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X31 drain_left.t8 plus.t15 source.t22 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X32 drain_right.t9 minus.t14 source.t15 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.7
X33 a_n3394_n4888# a_n3394_n4888# a_n3394_n4888# a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X34 drain_left.t7 plus.t16 source.t34 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X35 source.t5 minus.t15 drain_right.t8 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X36 drain_right.t7 minus.t16 source.t9 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X37 source.t7 minus.t17 drain_right.t6 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X38 source.t47 minus.t18 drain_right.t5 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X39 drain_left.t6 plus.t17 source.t32 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X40 source.t31 plus.t18 drain_left.t5 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X41 drain_left.t4 plus.t19 source.t30 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X42 source.t38 plus.t20 drain_left.t3 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.7
X43 drain_left.t2 plus.t21 source.t24 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X44 source.t16 minus.t19 drain_right.t4 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X45 a_n3394_n4888# a_n3394_n4888# a_n3394_n4888# a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.7
X46 drain_right.t3 minus.t20 source.t45 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X47 source.t3 minus.t21 drain_right.t2 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X48 source.t4 minus.t22 drain_right.t1 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X49 source.t46 minus.t23 drain_right.t0 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X50 source.t21 plus.t22 drain_left.t1 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
X51 source.t23 plus.t23 drain_left.t0 a_n3394_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.7
R0 plus.n11 plus.t7 771.048
R1 plus.n53 plus.t0 771.048
R2 plus.n40 plus.t2 744.691
R3 plus.n38 plus.t12 744.691
R4 plus.n2 plus.t5 744.691
R5 plus.n32 plus.t22 744.691
R6 plus.n4 plus.t10 744.691
R7 plus.n26 plus.t3 744.691
R8 plus.n6 plus.t13 744.691
R9 plus.n20 plus.t6 744.691
R10 plus.n8 plus.t11 744.691
R11 plus.n14 plus.t4 744.691
R12 plus.n10 plus.t16 744.691
R13 plus.n82 plus.t20 744.691
R14 plus.n80 plus.t19 744.691
R15 plus.n44 plus.t18 744.691
R16 plus.n74 plus.t17 744.691
R17 plus.n46 plus.t23 744.691
R18 plus.n68 plus.t9 744.691
R19 plus.n48 plus.t8 744.691
R20 plus.n62 plus.t15 744.691
R21 plus.n50 plus.t14 744.691
R22 plus.n56 plus.t21 744.691
R23 plus.n52 plus.t1 744.691
R24 plus.n13 plus.n12 161.3
R25 plus.n14 plus.n9 161.3
R26 plus.n16 plus.n15 161.3
R27 plus.n17 plus.n8 161.3
R28 plus.n19 plus.n18 161.3
R29 plus.n20 plus.n7 161.3
R30 plus.n22 plus.n21 161.3
R31 plus.n23 plus.n6 161.3
R32 plus.n25 plus.n24 161.3
R33 plus.n26 plus.n5 161.3
R34 plus.n28 plus.n27 161.3
R35 plus.n29 plus.n4 161.3
R36 plus.n31 plus.n30 161.3
R37 plus.n32 plus.n3 161.3
R38 plus.n34 plus.n33 161.3
R39 plus.n35 plus.n2 161.3
R40 plus.n37 plus.n36 161.3
R41 plus.n38 plus.n1 161.3
R42 plus.n39 plus.n0 161.3
R43 plus.n41 plus.n40 161.3
R44 plus.n55 plus.n54 161.3
R45 plus.n56 plus.n51 161.3
R46 plus.n58 plus.n57 161.3
R47 plus.n59 plus.n50 161.3
R48 plus.n61 plus.n60 161.3
R49 plus.n62 plus.n49 161.3
R50 plus.n64 plus.n63 161.3
R51 plus.n65 plus.n48 161.3
R52 plus.n67 plus.n66 161.3
R53 plus.n68 plus.n47 161.3
R54 plus.n70 plus.n69 161.3
R55 plus.n71 plus.n46 161.3
R56 plus.n73 plus.n72 161.3
R57 plus.n74 plus.n45 161.3
R58 plus.n76 plus.n75 161.3
R59 plus.n77 plus.n44 161.3
R60 plus.n79 plus.n78 161.3
R61 plus.n80 plus.n43 161.3
R62 plus.n81 plus.n42 161.3
R63 plus.n83 plus.n82 161.3
R64 plus.n40 plus.n39 46.0096
R65 plus.n82 plus.n81 46.0096
R66 plus.n12 plus.n11 45.0871
R67 plus.n54 plus.n53 45.0871
R68 plus.n38 plus.n37 41.6278
R69 plus.n13 plus.n10 41.6278
R70 plus.n80 plus.n79 41.6278
R71 plus.n55 plus.n52 41.6278
R72 plus plus.n83 39.0672
R73 plus.n33 plus.n2 37.246
R74 plus.n15 plus.n14 37.246
R75 plus.n75 plus.n44 37.246
R76 plus.n57 plus.n56 37.246
R77 plus.n32 plus.n31 32.8641
R78 plus.n19 plus.n8 32.8641
R79 plus.n74 plus.n73 32.8641
R80 plus.n61 plus.n50 32.8641
R81 plus.n27 plus.n4 28.4823
R82 plus.n21 plus.n20 28.4823
R83 plus.n69 plus.n46 28.4823
R84 plus.n63 plus.n62 28.4823
R85 plus.n25 plus.n6 24.1005
R86 plus.n26 plus.n25 24.1005
R87 plus.n68 plus.n67 24.1005
R88 plus.n67 plus.n48 24.1005
R89 plus.n27 plus.n26 19.7187
R90 plus.n21 plus.n6 19.7187
R91 plus.n69 plus.n68 19.7187
R92 plus.n63 plus.n48 19.7187
R93 plus plus.n41 15.3528
R94 plus.n31 plus.n4 15.3369
R95 plus.n20 plus.n19 15.3369
R96 plus.n73 plus.n46 15.3369
R97 plus.n62 plus.n61 15.3369
R98 plus.n11 plus.n10 14.1472
R99 plus.n53 plus.n52 14.1472
R100 plus.n33 plus.n32 10.955
R101 plus.n15 plus.n8 10.955
R102 plus.n75 plus.n74 10.955
R103 plus.n57 plus.n50 10.955
R104 plus.n37 plus.n2 6.57323
R105 plus.n14 plus.n13 6.57323
R106 plus.n79 plus.n44 6.57323
R107 plus.n56 plus.n55 6.57323
R108 plus.n39 plus.n38 2.19141
R109 plus.n81 plus.n80 2.19141
R110 plus.n12 plus.n9 0.189894
R111 plus.n16 plus.n9 0.189894
R112 plus.n17 plus.n16 0.189894
R113 plus.n18 plus.n17 0.189894
R114 plus.n18 plus.n7 0.189894
R115 plus.n22 plus.n7 0.189894
R116 plus.n23 plus.n22 0.189894
R117 plus.n24 plus.n23 0.189894
R118 plus.n24 plus.n5 0.189894
R119 plus.n28 plus.n5 0.189894
R120 plus.n29 plus.n28 0.189894
R121 plus.n30 plus.n29 0.189894
R122 plus.n30 plus.n3 0.189894
R123 plus.n34 plus.n3 0.189894
R124 plus.n35 plus.n34 0.189894
R125 plus.n36 plus.n35 0.189894
R126 plus.n36 plus.n1 0.189894
R127 plus.n1 plus.n0 0.189894
R128 plus.n41 plus.n0 0.189894
R129 plus.n83 plus.n42 0.189894
R130 plus.n43 plus.n42 0.189894
R131 plus.n78 plus.n43 0.189894
R132 plus.n78 plus.n77 0.189894
R133 plus.n77 plus.n76 0.189894
R134 plus.n76 plus.n45 0.189894
R135 plus.n72 plus.n45 0.189894
R136 plus.n72 plus.n71 0.189894
R137 plus.n71 plus.n70 0.189894
R138 plus.n70 plus.n47 0.189894
R139 plus.n66 plus.n47 0.189894
R140 plus.n66 plus.n65 0.189894
R141 plus.n65 plus.n64 0.189894
R142 plus.n64 plus.n49 0.189894
R143 plus.n60 plus.n49 0.189894
R144 plus.n60 plus.n59 0.189894
R145 plus.n59 plus.n58 0.189894
R146 plus.n58 plus.n51 0.189894
R147 plus.n54 plus.n51 0.189894
R148 source.n0 source.t44 44.1297
R149 source.n11 source.t40 44.1296
R150 source.n12 source.t15 44.1296
R151 source.n23 source.t5 44.1296
R152 source.n47 source.t2 44.1295
R153 source.n36 source.t14 44.1295
R154 source.n35 source.t25 44.1295
R155 source.n24 source.t38 44.1295
R156 source.n2 source.n1 43.1397
R157 source.n4 source.n3 43.1397
R158 source.n6 source.n5 43.1397
R159 source.n8 source.n7 43.1397
R160 source.n10 source.n9 43.1397
R161 source.n14 source.n13 43.1397
R162 source.n16 source.n15 43.1397
R163 source.n18 source.n17 43.1397
R164 source.n20 source.n19 43.1397
R165 source.n22 source.n21 43.1397
R166 source.n46 source.n45 43.1396
R167 source.n44 source.n43 43.1396
R168 source.n42 source.n41 43.1396
R169 source.n40 source.n39 43.1396
R170 source.n38 source.n37 43.1396
R171 source.n34 source.n33 43.1396
R172 source.n32 source.n31 43.1396
R173 source.n30 source.n29 43.1396
R174 source.n28 source.n27 43.1396
R175 source.n26 source.n25 43.1396
R176 source.n24 source.n23 28.2363
R177 source.n48 source.n0 22.5294
R178 source.n48 source.n47 5.7074
R179 source.n45 source.t1 0.9905
R180 source.n45 source.t20 0.9905
R181 source.n43 source.t9 0.9905
R182 source.n43 source.t47 0.9905
R183 source.n41 source.t45 0.9905
R184 source.n41 source.t46 0.9905
R185 source.n39 source.t6 0.9905
R186 source.n39 source.t19 0.9905
R187 source.n37 source.t11 0.9905
R188 source.n37 source.t12 0.9905
R189 source.n33 source.t24 0.9905
R190 source.n33 source.t33 0.9905
R191 source.n31 source.t22 0.9905
R192 source.n31 source.t35 0.9905
R193 source.n29 source.t43 0.9905
R194 source.n29 source.t41 0.9905
R195 source.n27 source.t32 0.9905
R196 source.n27 source.t23 0.9905
R197 source.n25 source.t30 0.9905
R198 source.n25 source.t31 0.9905
R199 source.n1 source.t28 0.9905
R200 source.n1 source.t37 0.9905
R201 source.n3 source.t27 0.9905
R202 source.n3 source.t21 0.9905
R203 source.n5 source.t36 0.9905
R204 source.n5 source.t42 0.9905
R205 source.n7 source.t26 0.9905
R206 source.n7 source.t39 0.9905
R207 source.n9 source.t34 0.9905
R208 source.n9 source.t29 0.9905
R209 source.n13 source.t17 0.9905
R210 source.n13 source.t8 0.9905
R211 source.n15 source.t10 0.9905
R212 source.n15 source.t3 0.9905
R213 source.n17 source.t18 0.9905
R214 source.n17 source.t4 0.9905
R215 source.n19 source.t0 0.9905
R216 source.n19 source.t16 0.9905
R217 source.n21 source.t13 0.9905
R218 source.n21 source.t7 0.9905
R219 source.n23 source.n22 0.888431
R220 source.n22 source.n20 0.888431
R221 source.n20 source.n18 0.888431
R222 source.n18 source.n16 0.888431
R223 source.n16 source.n14 0.888431
R224 source.n14 source.n12 0.888431
R225 source.n11 source.n10 0.888431
R226 source.n10 source.n8 0.888431
R227 source.n8 source.n6 0.888431
R228 source.n6 source.n4 0.888431
R229 source.n4 source.n2 0.888431
R230 source.n2 source.n0 0.888431
R231 source.n26 source.n24 0.888431
R232 source.n28 source.n26 0.888431
R233 source.n30 source.n28 0.888431
R234 source.n32 source.n30 0.888431
R235 source.n34 source.n32 0.888431
R236 source.n35 source.n34 0.888431
R237 source.n38 source.n36 0.888431
R238 source.n40 source.n38 0.888431
R239 source.n42 source.n40 0.888431
R240 source.n44 source.n42 0.888431
R241 source.n46 source.n44 0.888431
R242 source.n47 source.n46 0.888431
R243 source.n12 source.n11 0.470328
R244 source.n36 source.n35 0.470328
R245 source source.n48 0.188
R246 drain_left.n13 drain_left.n11 60.7064
R247 drain_left.n7 drain_left.n5 60.7063
R248 drain_left.n2 drain_left.n0 60.7063
R249 drain_left.n21 drain_left.n20 59.8185
R250 drain_left.n19 drain_left.n18 59.8185
R251 drain_left.n17 drain_left.n16 59.8185
R252 drain_left.n15 drain_left.n14 59.8185
R253 drain_left.n13 drain_left.n12 59.8185
R254 drain_left.n7 drain_left.n6 59.8184
R255 drain_left.n9 drain_left.n8 59.8184
R256 drain_left.n4 drain_left.n3 59.8184
R257 drain_left.n2 drain_left.n1 59.8184
R258 drain_left drain_left.n10 41.863
R259 drain_left drain_left.n21 6.54115
R260 drain_left.n5 drain_left.t22 0.9905
R261 drain_left.n5 drain_left.t23 0.9905
R262 drain_left.n6 drain_left.t9 0.9905
R263 drain_left.n6 drain_left.t2 0.9905
R264 drain_left.n8 drain_left.t15 0.9905
R265 drain_left.n8 drain_left.t8 0.9905
R266 drain_left.n3 drain_left.t0 0.9905
R267 drain_left.n3 drain_left.t14 0.9905
R268 drain_left.n1 drain_left.t5 0.9905
R269 drain_left.n1 drain_left.t6 0.9905
R270 drain_left.n0 drain_left.t3 0.9905
R271 drain_left.n0 drain_left.t4 0.9905
R272 drain_left.n20 drain_left.t11 0.9905
R273 drain_left.n20 drain_left.t21 0.9905
R274 drain_left.n18 drain_left.t1 0.9905
R275 drain_left.n18 drain_left.t18 0.9905
R276 drain_left.n16 drain_left.t20 0.9905
R277 drain_left.n16 drain_left.t13 0.9905
R278 drain_left.n14 drain_left.t17 0.9905
R279 drain_left.n14 drain_left.t10 0.9905
R280 drain_left.n12 drain_left.t19 0.9905
R281 drain_left.n12 drain_left.t12 0.9905
R282 drain_left.n11 drain_left.t16 0.9905
R283 drain_left.n11 drain_left.t7 0.9905
R284 drain_left.n9 drain_left.n7 0.888431
R285 drain_left.n4 drain_left.n2 0.888431
R286 drain_left.n15 drain_left.n13 0.888431
R287 drain_left.n17 drain_left.n15 0.888431
R288 drain_left.n19 drain_left.n17 0.888431
R289 drain_left.n21 drain_left.n19 0.888431
R290 drain_left.n10 drain_left.n9 0.389119
R291 drain_left.n10 drain_left.n4 0.389119
R292 minus.n11 minus.t14 771.048
R293 minus.n53 minus.t8 771.048
R294 minus.n10 minus.t2 744.691
R295 minus.n14 minus.t13 744.691
R296 minus.n16 minus.t21 744.691
R297 minus.n20 minus.t12 744.691
R298 minus.n22 minus.t22 744.691
R299 minus.n26 minus.t10 744.691
R300 minus.n28 minus.t19 744.691
R301 minus.n32 minus.t9 744.691
R302 minus.n34 minus.t17 744.691
R303 minus.n38 minus.t5 744.691
R304 minus.n40 minus.t15 744.691
R305 minus.n52 minus.t7 744.691
R306 minus.n56 minus.t0 744.691
R307 minus.n58 minus.t1 744.691
R308 minus.n62 minus.t4 744.691
R309 minus.n64 minus.t20 744.691
R310 minus.n68 minus.t23 744.691
R311 minus.n70 minus.t16 744.691
R312 minus.n74 minus.t18 744.691
R313 minus.n76 minus.t11 744.691
R314 minus.n80 minus.t3 744.691
R315 minus.n82 minus.t6 744.691
R316 minus.n41 minus.n40 161.3
R317 minus.n39 minus.n0 161.3
R318 minus.n38 minus.n37 161.3
R319 minus.n36 minus.n1 161.3
R320 minus.n35 minus.n34 161.3
R321 minus.n33 minus.n2 161.3
R322 minus.n32 minus.n31 161.3
R323 minus.n30 minus.n3 161.3
R324 minus.n29 minus.n28 161.3
R325 minus.n27 minus.n4 161.3
R326 minus.n26 minus.n25 161.3
R327 minus.n24 minus.n5 161.3
R328 minus.n23 minus.n22 161.3
R329 minus.n21 minus.n6 161.3
R330 minus.n20 minus.n19 161.3
R331 minus.n18 minus.n7 161.3
R332 minus.n17 minus.n16 161.3
R333 minus.n15 minus.n8 161.3
R334 minus.n14 minus.n13 161.3
R335 minus.n12 minus.n9 161.3
R336 minus.n83 minus.n82 161.3
R337 minus.n81 minus.n42 161.3
R338 minus.n80 minus.n79 161.3
R339 minus.n78 minus.n43 161.3
R340 minus.n77 minus.n76 161.3
R341 minus.n75 minus.n44 161.3
R342 minus.n74 minus.n73 161.3
R343 minus.n72 minus.n45 161.3
R344 minus.n71 minus.n70 161.3
R345 minus.n69 minus.n46 161.3
R346 minus.n68 minus.n67 161.3
R347 minus.n66 minus.n47 161.3
R348 minus.n65 minus.n64 161.3
R349 minus.n63 minus.n48 161.3
R350 minus.n62 minus.n61 161.3
R351 minus.n60 minus.n49 161.3
R352 minus.n59 minus.n58 161.3
R353 minus.n57 minus.n50 161.3
R354 minus.n56 minus.n55 161.3
R355 minus.n54 minus.n51 161.3
R356 minus.n84 minus.n41 48.2164
R357 minus.n40 minus.n39 46.0096
R358 minus.n82 minus.n81 46.0096
R359 minus.n12 minus.n11 45.0871
R360 minus.n54 minus.n53 45.0871
R361 minus.n10 minus.n9 41.6278
R362 minus.n38 minus.n1 41.6278
R363 minus.n52 minus.n51 41.6278
R364 minus.n80 minus.n43 41.6278
R365 minus.n15 minus.n14 37.246
R366 minus.n34 minus.n33 37.246
R367 minus.n57 minus.n56 37.246
R368 minus.n76 minus.n75 37.246
R369 minus.n16 minus.n7 32.8641
R370 minus.n32 minus.n3 32.8641
R371 minus.n58 minus.n49 32.8641
R372 minus.n74 minus.n45 32.8641
R373 minus.n21 minus.n20 28.4823
R374 minus.n28 minus.n27 28.4823
R375 minus.n63 minus.n62 28.4823
R376 minus.n70 minus.n69 28.4823
R377 minus.n26 minus.n5 24.1005
R378 minus.n22 minus.n5 24.1005
R379 minus.n64 minus.n47 24.1005
R380 minus.n68 minus.n47 24.1005
R381 minus.n22 minus.n21 19.7187
R382 minus.n27 minus.n26 19.7187
R383 minus.n64 minus.n63 19.7187
R384 minus.n69 minus.n68 19.7187
R385 minus.n20 minus.n7 15.3369
R386 minus.n28 minus.n3 15.3369
R387 minus.n62 minus.n49 15.3369
R388 minus.n70 minus.n45 15.3369
R389 minus.n11 minus.n10 14.1472
R390 minus.n53 minus.n52 14.1472
R391 minus.n16 minus.n15 10.955
R392 minus.n33 minus.n32 10.955
R393 minus.n58 minus.n57 10.955
R394 minus.n75 minus.n74 10.955
R395 minus.n84 minus.n83 6.67853
R396 minus.n14 minus.n9 6.57323
R397 minus.n34 minus.n1 6.57323
R398 minus.n56 minus.n51 6.57323
R399 minus.n76 minus.n43 6.57323
R400 minus.n39 minus.n38 2.19141
R401 minus.n81 minus.n80 2.19141
R402 minus.n41 minus.n0 0.189894
R403 minus.n37 minus.n0 0.189894
R404 minus.n37 minus.n36 0.189894
R405 minus.n36 minus.n35 0.189894
R406 minus.n35 minus.n2 0.189894
R407 minus.n31 minus.n2 0.189894
R408 minus.n31 minus.n30 0.189894
R409 minus.n30 minus.n29 0.189894
R410 minus.n29 minus.n4 0.189894
R411 minus.n25 minus.n4 0.189894
R412 minus.n25 minus.n24 0.189894
R413 minus.n24 minus.n23 0.189894
R414 minus.n23 minus.n6 0.189894
R415 minus.n19 minus.n6 0.189894
R416 minus.n19 minus.n18 0.189894
R417 minus.n18 minus.n17 0.189894
R418 minus.n17 minus.n8 0.189894
R419 minus.n13 minus.n8 0.189894
R420 minus.n13 minus.n12 0.189894
R421 minus.n55 minus.n54 0.189894
R422 minus.n55 minus.n50 0.189894
R423 minus.n59 minus.n50 0.189894
R424 minus.n60 minus.n59 0.189894
R425 minus.n61 minus.n60 0.189894
R426 minus.n61 minus.n48 0.189894
R427 minus.n65 minus.n48 0.189894
R428 minus.n66 minus.n65 0.189894
R429 minus.n67 minus.n66 0.189894
R430 minus.n67 minus.n46 0.189894
R431 minus.n71 minus.n46 0.189894
R432 minus.n72 minus.n71 0.189894
R433 minus.n73 minus.n72 0.189894
R434 minus.n73 minus.n44 0.189894
R435 minus.n77 minus.n44 0.189894
R436 minus.n78 minus.n77 0.189894
R437 minus.n79 minus.n78 0.189894
R438 minus.n79 minus.n42 0.189894
R439 minus.n83 minus.n42 0.189894
R440 minus minus.n84 0.188
R441 drain_right.n13 drain_right.n11 60.7064
R442 drain_right.n7 drain_right.n5 60.7063
R443 drain_right.n2 drain_right.n0 60.7063
R444 drain_right.n13 drain_right.n12 59.8185
R445 drain_right.n15 drain_right.n14 59.8185
R446 drain_right.n17 drain_right.n16 59.8185
R447 drain_right.n19 drain_right.n18 59.8185
R448 drain_right.n21 drain_right.n20 59.8185
R449 drain_right.n7 drain_right.n6 59.8184
R450 drain_right.n9 drain_right.n8 59.8184
R451 drain_right.n4 drain_right.n3 59.8184
R452 drain_right.n2 drain_right.n1 59.8184
R453 drain_right drain_right.n10 41.3098
R454 drain_right drain_right.n21 6.54115
R455 drain_right.n5 drain_right.t20 0.9905
R456 drain_right.n5 drain_right.t17 0.9905
R457 drain_right.n6 drain_right.t5 0.9905
R458 drain_right.n6 drain_right.t12 0.9905
R459 drain_right.n8 drain_right.t0 0.9905
R460 drain_right.n8 drain_right.t7 0.9905
R461 drain_right.n3 drain_right.t19 0.9905
R462 drain_right.n3 drain_right.t3 0.9905
R463 drain_right.n1 drain_right.t23 0.9905
R464 drain_right.n1 drain_right.t22 0.9905
R465 drain_right.n0 drain_right.t15 0.9905
R466 drain_right.n0 drain_right.t16 0.9905
R467 drain_right.n11 drain_right.t21 0.9905
R468 drain_right.n11 drain_right.t9 0.9905
R469 drain_right.n12 drain_right.t2 0.9905
R470 drain_right.n12 drain_right.t10 0.9905
R471 drain_right.n14 drain_right.t1 0.9905
R472 drain_right.n14 drain_right.t11 0.9905
R473 drain_right.n16 drain_right.t4 0.9905
R474 drain_right.n16 drain_right.t13 0.9905
R475 drain_right.n18 drain_right.t6 0.9905
R476 drain_right.n18 drain_right.t14 0.9905
R477 drain_right.n20 drain_right.t8 0.9905
R478 drain_right.n20 drain_right.t18 0.9905
R479 drain_right.n9 drain_right.n7 0.888431
R480 drain_right.n4 drain_right.n2 0.888431
R481 drain_right.n21 drain_right.n19 0.888431
R482 drain_right.n19 drain_right.n17 0.888431
R483 drain_right.n17 drain_right.n15 0.888431
R484 drain_right.n15 drain_right.n13 0.888431
R485 drain_right.n10 drain_right.n9 0.389119
R486 drain_right.n10 drain_right.n4 0.389119
C0 drain_right drain_left 1.87044f
C1 drain_left minus 0.174517f
C2 drain_left source 44.0863f
C3 drain_right plus 0.498726f
C4 plus minus 8.86237f
C5 plus source 24.3699f
C6 plus drain_left 24.717598f
C7 drain_right minus 24.3772f
C8 drain_right source 44.0888f
C9 minus source 24.3559f
C10 drain_right a_n3394_n4888# 9.331349f
C11 drain_left a_n3394_n4888# 9.79634f
C12 source a_n3394_n4888# 14.040558f
C13 minus a_n3394_n4888# 14.28508f
C14 plus a_n3394_n4888# 16.557669f
C15 drain_right.t15 a_n3394_n4888# 0.429989f
C16 drain_right.t16 a_n3394_n4888# 0.429989f
C17 drain_right.n0 a_n3394_n4888# 3.93685f
C18 drain_right.t23 a_n3394_n4888# 0.429989f
C19 drain_right.t22 a_n3394_n4888# 0.429989f
C20 drain_right.n1 a_n3394_n4888# 3.93105f
C21 drain_right.n2 a_n3394_n4888# 0.775696f
C22 drain_right.t19 a_n3394_n4888# 0.429989f
C23 drain_right.t3 a_n3394_n4888# 0.429989f
C24 drain_right.n3 a_n3394_n4888# 3.93105f
C25 drain_right.n4 a_n3394_n4888# 0.343117f
C26 drain_right.t20 a_n3394_n4888# 0.429989f
C27 drain_right.t17 a_n3394_n4888# 0.429989f
C28 drain_right.n5 a_n3394_n4888# 3.93685f
C29 drain_right.t5 a_n3394_n4888# 0.429989f
C30 drain_right.t12 a_n3394_n4888# 0.429989f
C31 drain_right.n6 a_n3394_n4888# 3.93105f
C32 drain_right.n7 a_n3394_n4888# 0.775696f
C33 drain_right.t0 a_n3394_n4888# 0.429989f
C34 drain_right.t7 a_n3394_n4888# 0.429989f
C35 drain_right.n8 a_n3394_n4888# 3.93105f
C36 drain_right.n9 a_n3394_n4888# 0.343117f
C37 drain_right.n10 a_n3394_n4888# 2.27434f
C38 drain_right.t21 a_n3394_n4888# 0.429989f
C39 drain_right.t9 a_n3394_n4888# 0.429989f
C40 drain_right.n11 a_n3394_n4888# 3.93684f
C41 drain_right.t2 a_n3394_n4888# 0.429989f
C42 drain_right.t10 a_n3394_n4888# 0.429989f
C43 drain_right.n12 a_n3394_n4888# 3.93105f
C44 drain_right.n13 a_n3394_n4888# 0.775707f
C45 drain_right.t1 a_n3394_n4888# 0.429989f
C46 drain_right.t11 a_n3394_n4888# 0.429989f
C47 drain_right.n14 a_n3394_n4888# 3.93105f
C48 drain_right.n15 a_n3394_n4888# 0.385272f
C49 drain_right.t4 a_n3394_n4888# 0.429989f
C50 drain_right.t13 a_n3394_n4888# 0.429989f
C51 drain_right.n16 a_n3394_n4888# 3.93105f
C52 drain_right.n17 a_n3394_n4888# 0.385272f
C53 drain_right.t6 a_n3394_n4888# 0.429989f
C54 drain_right.t14 a_n3394_n4888# 0.429989f
C55 drain_right.n18 a_n3394_n4888# 3.93105f
C56 drain_right.n19 a_n3394_n4888# 0.385272f
C57 drain_right.t8 a_n3394_n4888# 0.429989f
C58 drain_right.t18 a_n3394_n4888# 0.429989f
C59 drain_right.n20 a_n3394_n4888# 3.93105f
C60 drain_right.n21 a_n3394_n4888# 0.625916f
C61 minus.n0 a_n3394_n4888# 0.038955f
C62 minus.n1 a_n3394_n4888# 0.00884f
C63 minus.t5 a_n3394_n4888# 1.54443f
C64 minus.n2 a_n3394_n4888# 0.038955f
C65 minus.n3 a_n3394_n4888# 0.00884f
C66 minus.t9 a_n3394_n4888# 1.54443f
C67 minus.n4 a_n3394_n4888# 0.038955f
C68 minus.n5 a_n3394_n4888# 0.00884f
C69 minus.t10 a_n3394_n4888# 1.54443f
C70 minus.n6 a_n3394_n4888# 0.038955f
C71 minus.n7 a_n3394_n4888# 0.00884f
C72 minus.t12 a_n3394_n4888# 1.54443f
C73 minus.n8 a_n3394_n4888# 0.038955f
C74 minus.n9 a_n3394_n4888# 0.00884f
C75 minus.t13 a_n3394_n4888# 1.54443f
C76 minus.t14 a_n3394_n4888# 1.56414f
C77 minus.t2 a_n3394_n4888# 1.54443f
C78 minus.n10 a_n3394_n4888# 0.583883f
C79 minus.n11 a_n3394_n4888# 0.558275f
C80 minus.n12 a_n3394_n4888# 0.167703f
C81 minus.n13 a_n3394_n4888# 0.038955f
C82 minus.n14 a_n3394_n4888# 0.575911f
C83 minus.n15 a_n3394_n4888# 0.00884f
C84 minus.t21 a_n3394_n4888# 1.54443f
C85 minus.n16 a_n3394_n4888# 0.575911f
C86 minus.n17 a_n3394_n4888# 0.038955f
C87 minus.n18 a_n3394_n4888# 0.038955f
C88 minus.n19 a_n3394_n4888# 0.038955f
C89 minus.n20 a_n3394_n4888# 0.575911f
C90 minus.n21 a_n3394_n4888# 0.00884f
C91 minus.t22 a_n3394_n4888# 1.54443f
C92 minus.n22 a_n3394_n4888# 0.575911f
C93 minus.n23 a_n3394_n4888# 0.038955f
C94 minus.n24 a_n3394_n4888# 0.038955f
C95 minus.n25 a_n3394_n4888# 0.038955f
C96 minus.n26 a_n3394_n4888# 0.575911f
C97 minus.n27 a_n3394_n4888# 0.00884f
C98 minus.t19 a_n3394_n4888# 1.54443f
C99 minus.n28 a_n3394_n4888# 0.575911f
C100 minus.n29 a_n3394_n4888# 0.038955f
C101 minus.n30 a_n3394_n4888# 0.038955f
C102 minus.n31 a_n3394_n4888# 0.038955f
C103 minus.n32 a_n3394_n4888# 0.575911f
C104 minus.n33 a_n3394_n4888# 0.00884f
C105 minus.t17 a_n3394_n4888# 1.54443f
C106 minus.n34 a_n3394_n4888# 0.575911f
C107 minus.n35 a_n3394_n4888# 0.038955f
C108 minus.n36 a_n3394_n4888# 0.038955f
C109 minus.n37 a_n3394_n4888# 0.038955f
C110 minus.n38 a_n3394_n4888# 0.575911f
C111 minus.n39 a_n3394_n4888# 0.00884f
C112 minus.t15 a_n3394_n4888# 1.54443f
C113 minus.n40 a_n3394_n4888# 0.576272f
C114 minus.n41 a_n3394_n4888# 2.10754f
C115 minus.n42 a_n3394_n4888# 0.038955f
C116 minus.n43 a_n3394_n4888# 0.00884f
C117 minus.n44 a_n3394_n4888# 0.038955f
C118 minus.n45 a_n3394_n4888# 0.00884f
C119 minus.n46 a_n3394_n4888# 0.038955f
C120 minus.n47 a_n3394_n4888# 0.00884f
C121 minus.n48 a_n3394_n4888# 0.038955f
C122 minus.n49 a_n3394_n4888# 0.00884f
C123 minus.n50 a_n3394_n4888# 0.038955f
C124 minus.n51 a_n3394_n4888# 0.00884f
C125 minus.t8 a_n3394_n4888# 1.56414f
C126 minus.t7 a_n3394_n4888# 1.54443f
C127 minus.n52 a_n3394_n4888# 0.583883f
C128 minus.n53 a_n3394_n4888# 0.558275f
C129 minus.n54 a_n3394_n4888# 0.167703f
C130 minus.n55 a_n3394_n4888# 0.038955f
C131 minus.t0 a_n3394_n4888# 1.54443f
C132 minus.n56 a_n3394_n4888# 0.575911f
C133 minus.n57 a_n3394_n4888# 0.00884f
C134 minus.t1 a_n3394_n4888# 1.54443f
C135 minus.n58 a_n3394_n4888# 0.575911f
C136 minus.n59 a_n3394_n4888# 0.038955f
C137 minus.n60 a_n3394_n4888# 0.038955f
C138 minus.n61 a_n3394_n4888# 0.038955f
C139 minus.t4 a_n3394_n4888# 1.54443f
C140 minus.n62 a_n3394_n4888# 0.575911f
C141 minus.n63 a_n3394_n4888# 0.00884f
C142 minus.t20 a_n3394_n4888# 1.54443f
C143 minus.n64 a_n3394_n4888# 0.575911f
C144 minus.n65 a_n3394_n4888# 0.038955f
C145 minus.n66 a_n3394_n4888# 0.038955f
C146 minus.n67 a_n3394_n4888# 0.038955f
C147 minus.t23 a_n3394_n4888# 1.54443f
C148 minus.n68 a_n3394_n4888# 0.575911f
C149 minus.n69 a_n3394_n4888# 0.00884f
C150 minus.t16 a_n3394_n4888# 1.54443f
C151 minus.n70 a_n3394_n4888# 0.575911f
C152 minus.n71 a_n3394_n4888# 0.038955f
C153 minus.n72 a_n3394_n4888# 0.038955f
C154 minus.n73 a_n3394_n4888# 0.038955f
C155 minus.t18 a_n3394_n4888# 1.54443f
C156 minus.n74 a_n3394_n4888# 0.575911f
C157 minus.n75 a_n3394_n4888# 0.00884f
C158 minus.t11 a_n3394_n4888# 1.54443f
C159 minus.n76 a_n3394_n4888# 0.575911f
C160 minus.n77 a_n3394_n4888# 0.038955f
C161 minus.n78 a_n3394_n4888# 0.038955f
C162 minus.n79 a_n3394_n4888# 0.038955f
C163 minus.t3 a_n3394_n4888# 1.54443f
C164 minus.n80 a_n3394_n4888# 0.575911f
C165 minus.n81 a_n3394_n4888# 0.00884f
C166 minus.t6 a_n3394_n4888# 1.54443f
C167 minus.n82 a_n3394_n4888# 0.576272f
C168 minus.n83 a_n3394_n4888# 0.270926f
C169 minus.n84 a_n3394_n4888# 2.47248f
C170 drain_left.t3 a_n3394_n4888# 0.431202f
C171 drain_left.t4 a_n3394_n4888# 0.431202f
C172 drain_left.n0 a_n3394_n4888# 3.94796f
C173 drain_left.t5 a_n3394_n4888# 0.431202f
C174 drain_left.t6 a_n3394_n4888# 0.431202f
C175 drain_left.n1 a_n3394_n4888# 3.94214f
C176 drain_left.n2 a_n3394_n4888# 0.777884f
C177 drain_left.t0 a_n3394_n4888# 0.431202f
C178 drain_left.t14 a_n3394_n4888# 0.431202f
C179 drain_left.n3 a_n3394_n4888# 3.94214f
C180 drain_left.n4 a_n3394_n4888# 0.344085f
C181 drain_left.t22 a_n3394_n4888# 0.431202f
C182 drain_left.t23 a_n3394_n4888# 0.431202f
C183 drain_left.n5 a_n3394_n4888# 3.94796f
C184 drain_left.t9 a_n3394_n4888# 0.431202f
C185 drain_left.t2 a_n3394_n4888# 0.431202f
C186 drain_left.n6 a_n3394_n4888# 3.94214f
C187 drain_left.n7 a_n3394_n4888# 0.777884f
C188 drain_left.t15 a_n3394_n4888# 0.431202f
C189 drain_left.t8 a_n3394_n4888# 0.431202f
C190 drain_left.n8 a_n3394_n4888# 3.94214f
C191 drain_left.n9 a_n3394_n4888# 0.344085f
C192 drain_left.n10 a_n3394_n4888# 2.33638f
C193 drain_left.t16 a_n3394_n4888# 0.431202f
C194 drain_left.t7 a_n3394_n4888# 0.431202f
C195 drain_left.n11 a_n3394_n4888# 3.94795f
C196 drain_left.t19 a_n3394_n4888# 0.431202f
C197 drain_left.t12 a_n3394_n4888# 0.431202f
C198 drain_left.n12 a_n3394_n4888# 3.94214f
C199 drain_left.n13 a_n3394_n4888# 0.777895f
C200 drain_left.t17 a_n3394_n4888# 0.431202f
C201 drain_left.t10 a_n3394_n4888# 0.431202f
C202 drain_left.n14 a_n3394_n4888# 3.94214f
C203 drain_left.n15 a_n3394_n4888# 0.386359f
C204 drain_left.t20 a_n3394_n4888# 0.431202f
C205 drain_left.t13 a_n3394_n4888# 0.431202f
C206 drain_left.n16 a_n3394_n4888# 3.94214f
C207 drain_left.n17 a_n3394_n4888# 0.386359f
C208 drain_left.t1 a_n3394_n4888# 0.431202f
C209 drain_left.t18 a_n3394_n4888# 0.431202f
C210 drain_left.n18 a_n3394_n4888# 3.94214f
C211 drain_left.n19 a_n3394_n4888# 0.386359f
C212 drain_left.t11 a_n3394_n4888# 0.431202f
C213 drain_left.t21 a_n3394_n4888# 0.431202f
C214 drain_left.n20 a_n3394_n4888# 3.94214f
C215 drain_left.n21 a_n3394_n4888# 0.627682f
C216 source.t44 a_n3394_n4888# 4.35183f
C217 source.n0 a_n3394_n4888# 1.89317f
C218 source.t28 a_n3394_n4888# 0.380791f
C219 source.t37 a_n3394_n4888# 0.380791f
C220 source.n1 a_n3394_n4888# 3.40444f
C221 source.n2 a_n3394_n4888# 0.385278f
C222 source.t27 a_n3394_n4888# 0.380791f
C223 source.t21 a_n3394_n4888# 0.380791f
C224 source.n3 a_n3394_n4888# 3.40444f
C225 source.n4 a_n3394_n4888# 0.385278f
C226 source.t36 a_n3394_n4888# 0.380791f
C227 source.t42 a_n3394_n4888# 0.380791f
C228 source.n5 a_n3394_n4888# 3.40444f
C229 source.n6 a_n3394_n4888# 0.385278f
C230 source.t26 a_n3394_n4888# 0.380791f
C231 source.t39 a_n3394_n4888# 0.380791f
C232 source.n7 a_n3394_n4888# 3.40444f
C233 source.n8 a_n3394_n4888# 0.385278f
C234 source.t34 a_n3394_n4888# 0.380791f
C235 source.t29 a_n3394_n4888# 0.380791f
C236 source.n9 a_n3394_n4888# 3.40444f
C237 source.n10 a_n3394_n4888# 0.385278f
C238 source.t40 a_n3394_n4888# 4.35183f
C239 source.n11 a_n3394_n4888# 0.443941f
C240 source.t15 a_n3394_n4888# 4.35183f
C241 source.n12 a_n3394_n4888# 0.443941f
C242 source.t17 a_n3394_n4888# 0.380791f
C243 source.t8 a_n3394_n4888# 0.380791f
C244 source.n13 a_n3394_n4888# 3.40444f
C245 source.n14 a_n3394_n4888# 0.385278f
C246 source.t10 a_n3394_n4888# 0.380791f
C247 source.t3 a_n3394_n4888# 0.380791f
C248 source.n15 a_n3394_n4888# 3.40444f
C249 source.n16 a_n3394_n4888# 0.385278f
C250 source.t18 a_n3394_n4888# 0.380791f
C251 source.t4 a_n3394_n4888# 0.380791f
C252 source.n17 a_n3394_n4888# 3.40444f
C253 source.n18 a_n3394_n4888# 0.385278f
C254 source.t0 a_n3394_n4888# 0.380791f
C255 source.t16 a_n3394_n4888# 0.380791f
C256 source.n19 a_n3394_n4888# 3.40444f
C257 source.n20 a_n3394_n4888# 0.385278f
C258 source.t13 a_n3394_n4888# 0.380791f
C259 source.t7 a_n3394_n4888# 0.380791f
C260 source.n21 a_n3394_n4888# 3.40444f
C261 source.n22 a_n3394_n4888# 0.385278f
C262 source.t5 a_n3394_n4888# 4.35183f
C263 source.n23 a_n3394_n4888# 2.33149f
C264 source.t38 a_n3394_n4888# 4.35181f
C265 source.n24 a_n3394_n4888# 2.33151f
C266 source.t30 a_n3394_n4888# 0.380791f
C267 source.t31 a_n3394_n4888# 0.380791f
C268 source.n25 a_n3394_n4888# 3.40444f
C269 source.n26 a_n3394_n4888# 0.385272f
C270 source.t32 a_n3394_n4888# 0.380791f
C271 source.t23 a_n3394_n4888# 0.380791f
C272 source.n27 a_n3394_n4888# 3.40444f
C273 source.n28 a_n3394_n4888# 0.385272f
C274 source.t43 a_n3394_n4888# 0.380791f
C275 source.t41 a_n3394_n4888# 0.380791f
C276 source.n29 a_n3394_n4888# 3.40444f
C277 source.n30 a_n3394_n4888# 0.385272f
C278 source.t22 a_n3394_n4888# 0.380791f
C279 source.t35 a_n3394_n4888# 0.380791f
C280 source.n31 a_n3394_n4888# 3.40444f
C281 source.n32 a_n3394_n4888# 0.385272f
C282 source.t24 a_n3394_n4888# 0.380791f
C283 source.t33 a_n3394_n4888# 0.380791f
C284 source.n33 a_n3394_n4888# 3.40444f
C285 source.n34 a_n3394_n4888# 0.385272f
C286 source.t25 a_n3394_n4888# 4.35181f
C287 source.n35 a_n3394_n4888# 0.443965f
C288 source.t14 a_n3394_n4888# 4.35181f
C289 source.n36 a_n3394_n4888# 0.443965f
C290 source.t11 a_n3394_n4888# 0.380791f
C291 source.t12 a_n3394_n4888# 0.380791f
C292 source.n37 a_n3394_n4888# 3.40444f
C293 source.n38 a_n3394_n4888# 0.385272f
C294 source.t6 a_n3394_n4888# 0.380791f
C295 source.t19 a_n3394_n4888# 0.380791f
C296 source.n39 a_n3394_n4888# 3.40444f
C297 source.n40 a_n3394_n4888# 0.385272f
C298 source.t45 a_n3394_n4888# 0.380791f
C299 source.t46 a_n3394_n4888# 0.380791f
C300 source.n41 a_n3394_n4888# 3.40444f
C301 source.n42 a_n3394_n4888# 0.385272f
C302 source.t9 a_n3394_n4888# 0.380791f
C303 source.t47 a_n3394_n4888# 0.380791f
C304 source.n43 a_n3394_n4888# 3.40444f
C305 source.n44 a_n3394_n4888# 0.385272f
C306 source.t1 a_n3394_n4888# 0.380791f
C307 source.t20 a_n3394_n4888# 0.380791f
C308 source.n45 a_n3394_n4888# 3.40444f
C309 source.n46 a_n3394_n4888# 0.385272f
C310 source.t2 a_n3394_n4888# 4.35181f
C311 source.n47 a_n3394_n4888# 0.601129f
C312 source.n48 a_n3394_n4888# 2.18585f
C313 plus.n0 a_n3394_n4888# 0.039211f
C314 plus.t2 a_n3394_n4888# 1.55458f
C315 plus.t12 a_n3394_n4888# 1.55458f
C316 plus.n1 a_n3394_n4888# 0.039211f
C317 plus.t5 a_n3394_n4888# 1.55458f
C318 plus.n2 a_n3394_n4888# 0.579697f
C319 plus.n3 a_n3394_n4888# 0.039211f
C320 plus.t22 a_n3394_n4888# 1.55458f
C321 plus.t10 a_n3394_n4888# 1.55458f
C322 plus.n4 a_n3394_n4888# 0.579697f
C323 plus.n5 a_n3394_n4888# 0.039211f
C324 plus.t3 a_n3394_n4888# 1.55458f
C325 plus.t13 a_n3394_n4888# 1.55458f
C326 plus.n6 a_n3394_n4888# 0.579697f
C327 plus.n7 a_n3394_n4888# 0.039211f
C328 plus.t6 a_n3394_n4888# 1.55458f
C329 plus.t11 a_n3394_n4888# 1.55458f
C330 plus.n8 a_n3394_n4888# 0.579697f
C331 plus.n9 a_n3394_n4888# 0.039211f
C332 plus.t4 a_n3394_n4888# 1.55458f
C333 plus.t16 a_n3394_n4888# 1.55458f
C334 plus.n10 a_n3394_n4888# 0.587721f
C335 plus.t7 a_n3394_n4888# 1.57442f
C336 plus.n11 a_n3394_n4888# 0.561944f
C337 plus.n12 a_n3394_n4888# 0.168805f
C338 plus.n13 a_n3394_n4888# 0.008898f
C339 plus.n14 a_n3394_n4888# 0.579697f
C340 plus.n15 a_n3394_n4888# 0.008898f
C341 plus.n16 a_n3394_n4888# 0.039211f
C342 plus.n17 a_n3394_n4888# 0.039211f
C343 plus.n18 a_n3394_n4888# 0.039211f
C344 plus.n19 a_n3394_n4888# 0.008898f
C345 plus.n20 a_n3394_n4888# 0.579697f
C346 plus.n21 a_n3394_n4888# 0.008898f
C347 plus.n22 a_n3394_n4888# 0.039211f
C348 plus.n23 a_n3394_n4888# 0.039211f
C349 plus.n24 a_n3394_n4888# 0.039211f
C350 plus.n25 a_n3394_n4888# 0.008898f
C351 plus.n26 a_n3394_n4888# 0.579697f
C352 plus.n27 a_n3394_n4888# 0.008898f
C353 plus.n28 a_n3394_n4888# 0.039211f
C354 plus.n29 a_n3394_n4888# 0.039211f
C355 plus.n30 a_n3394_n4888# 0.039211f
C356 plus.n31 a_n3394_n4888# 0.008898f
C357 plus.n32 a_n3394_n4888# 0.579697f
C358 plus.n33 a_n3394_n4888# 0.008898f
C359 plus.n34 a_n3394_n4888# 0.039211f
C360 plus.n35 a_n3394_n4888# 0.039211f
C361 plus.n36 a_n3394_n4888# 0.039211f
C362 plus.n37 a_n3394_n4888# 0.008898f
C363 plus.n38 a_n3394_n4888# 0.579697f
C364 plus.n39 a_n3394_n4888# 0.008898f
C365 plus.n40 a_n3394_n4888# 0.58006f
C366 plus.n41 a_n3394_n4888# 0.61144f
C367 plus.n42 a_n3394_n4888# 0.039211f
C368 plus.t20 a_n3394_n4888# 1.55458f
C369 plus.n43 a_n3394_n4888# 0.039211f
C370 plus.t19 a_n3394_n4888# 1.55458f
C371 plus.t18 a_n3394_n4888# 1.55458f
C372 plus.n44 a_n3394_n4888# 0.579697f
C373 plus.n45 a_n3394_n4888# 0.039211f
C374 plus.t17 a_n3394_n4888# 1.55458f
C375 plus.t23 a_n3394_n4888# 1.55458f
C376 plus.n46 a_n3394_n4888# 0.579697f
C377 plus.n47 a_n3394_n4888# 0.039211f
C378 plus.t9 a_n3394_n4888# 1.55458f
C379 plus.t8 a_n3394_n4888# 1.55458f
C380 plus.n48 a_n3394_n4888# 0.579697f
C381 plus.n49 a_n3394_n4888# 0.039211f
C382 plus.t15 a_n3394_n4888# 1.55458f
C383 plus.t14 a_n3394_n4888# 1.55458f
C384 plus.n50 a_n3394_n4888# 0.579697f
C385 plus.n51 a_n3394_n4888# 0.039211f
C386 plus.t21 a_n3394_n4888# 1.55458f
C387 plus.t1 a_n3394_n4888# 1.55458f
C388 plus.n52 a_n3394_n4888# 0.587721f
C389 plus.t0 a_n3394_n4888# 1.57442f
C390 plus.n53 a_n3394_n4888# 0.561944f
C391 plus.n54 a_n3394_n4888# 0.168805f
C392 plus.n55 a_n3394_n4888# 0.008898f
C393 plus.n56 a_n3394_n4888# 0.579697f
C394 plus.n57 a_n3394_n4888# 0.008898f
C395 plus.n58 a_n3394_n4888# 0.039211f
C396 plus.n59 a_n3394_n4888# 0.039211f
C397 plus.n60 a_n3394_n4888# 0.039211f
C398 plus.n61 a_n3394_n4888# 0.008898f
C399 plus.n62 a_n3394_n4888# 0.579697f
C400 plus.n63 a_n3394_n4888# 0.008898f
C401 plus.n64 a_n3394_n4888# 0.039211f
C402 plus.n65 a_n3394_n4888# 0.039211f
C403 plus.n66 a_n3394_n4888# 0.039211f
C404 plus.n67 a_n3394_n4888# 0.008898f
C405 plus.n68 a_n3394_n4888# 0.579697f
C406 plus.n69 a_n3394_n4888# 0.008898f
C407 plus.n70 a_n3394_n4888# 0.039211f
C408 plus.n71 a_n3394_n4888# 0.039211f
C409 plus.n72 a_n3394_n4888# 0.039211f
C410 plus.n73 a_n3394_n4888# 0.008898f
C411 plus.n74 a_n3394_n4888# 0.579697f
C412 plus.n75 a_n3394_n4888# 0.008898f
C413 plus.n76 a_n3394_n4888# 0.039211f
C414 plus.n77 a_n3394_n4888# 0.039211f
C415 plus.n78 a_n3394_n4888# 0.039211f
C416 plus.n79 a_n3394_n4888# 0.008898f
C417 plus.n80 a_n3394_n4888# 0.579697f
C418 plus.n81 a_n3394_n4888# 0.008898f
C419 plus.n82 a_n3394_n4888# 0.58006f
C420 plus.n83 a_n3394_n4888# 1.71967f
.ends

