* NGSPICE file created from diffpair576.ext - technology: sky130A

.subckt diffpair576 minus drain_right drain_left source plus
X0 drain_left.t13 plus.t0 source.t16 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X1 drain_left.t12 plus.t1 source.t25 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X2 drain_right.t13 minus.t0 source.t0 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X3 drain_right.t12 minus.t1 source.t8 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X4 source.t17 plus.t2 drain_left.t11 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X5 drain_left.t10 plus.t3 source.t20 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X6 source.t22 plus.t4 drain_left.t9 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X7 drain_right.t11 minus.t2 source.t3 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X8 source.t9 minus.t3 drain_right.t10 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X9 drain_right.t9 minus.t4 source.t12 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X10 source.t1 minus.t5 drain_right.t8 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X11 a_n1564_n4888# a_n1564_n4888# a_n1564_n4888# a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.2
X12 a_n1564_n4888# a_n1564_n4888# a_n1564_n4888# a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X13 source.t11 minus.t6 drain_right.t7 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X14 source.t2 minus.t7 drain_right.t6 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X15 source.t26 plus.t5 drain_left.t8 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X16 drain_left.t7 plus.t6 source.t14 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X17 source.t5 minus.t8 drain_right.t5 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X18 drain_right.t4 minus.t9 source.t13 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X19 drain_right.t3 minus.t10 source.t7 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X20 drain_right.t2 minus.t11 source.t10 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X21 drain_right.t1 minus.t12 source.t4 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X22 a_n1564_n4888# a_n1564_n4888# a_n1564_n4888# a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X23 drain_left.t6 plus.t7 source.t18 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X24 source.t21 plus.t8 drain_left.t5 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X25 source.t6 minus.t13 drain_right.t0 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X26 source.t24 plus.t9 drain_left.t4 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X27 source.t19 plus.t10 drain_left.t3 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X28 a_n1564_n4888# a_n1564_n4888# a_n1564_n4888# a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X29 drain_left.t2 plus.t11 source.t27 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X30 drain_left.t1 plus.t12 source.t15 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X31 drain_left.t0 plus.t13 source.t23 a_n1564_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
R0 plus.n3 plus.t6 2616.31
R1 plus.n14 plus.t3 2616.31
R2 plus.n19 plus.t0 2616.31
R3 plus.n30 plus.t11 2616.31
R4 plus.n4 plus.t4 2566.65
R5 plus.n6 plus.t12 2566.65
R6 plus.n1 plus.t8 2566.65
R7 plus.n11 plus.t7 2566.65
R8 plus.n13 plus.t5 2566.65
R9 plus.n20 plus.t2 2566.65
R10 plus.n22 plus.t1 2566.65
R11 plus.n17 plus.t9 2566.65
R12 plus.n27 plus.t13 2566.65
R13 plus.n29 plus.t10 2566.65
R14 plus.n3 plus.n2 161.489
R15 plus.n19 plus.n18 161.489
R16 plus.n5 plus.n2 161.3
R17 plus.n8 plus.n7 161.3
R18 plus.n10 plus.n9 161.3
R19 plus.n12 plus.n0 161.3
R20 plus.n15 plus.n14 161.3
R21 plus.n21 plus.n18 161.3
R22 plus.n24 plus.n23 161.3
R23 plus.n26 plus.n25 161.3
R24 plus.n28 plus.n16 161.3
R25 plus.n31 plus.n30 161.3
R26 plus.n5 plus.n4 45.2793
R27 plus.n13 plus.n12 45.2793
R28 plus.n29 plus.n28 45.2793
R29 plus.n21 plus.n20 45.2793
R30 plus.n7 plus.n6 40.8975
R31 plus.n11 plus.n10 40.8975
R32 plus.n27 plus.n26 40.8975
R33 plus.n23 plus.n22 40.8975
R34 plus.n7 plus.n1 36.5157
R35 plus.n10 plus.n1 36.5157
R36 plus.n26 plus.n17 36.5157
R37 plus.n23 plus.n17 36.5157
R38 plus.n6 plus.n5 32.1338
R39 plus.n12 plus.n11 32.1338
R40 plus.n28 plus.n27 32.1338
R41 plus.n22 plus.n21 32.1338
R42 plus plus.n31 31.9176
R43 plus.n4 plus.n3 27.752
R44 plus.n14 plus.n13 27.752
R45 plus.n30 plus.n29 27.752
R46 plus.n20 plus.n19 27.752
R47 plus plus.n15 15.135
R48 plus.n8 plus.n2 0.189894
R49 plus.n9 plus.n8 0.189894
R50 plus.n9 plus.n0 0.189894
R51 plus.n15 plus.n0 0.189894
R52 plus.n31 plus.n16 0.189894
R53 plus.n25 plus.n16 0.189894
R54 plus.n25 plus.n24 0.189894
R55 plus.n24 plus.n18 0.189894
R56 source.n0 source.t20 44.1297
R57 source.n7 source.t7 44.1296
R58 source.n27 source.t13 44.1295
R59 source.n20 source.t16 44.1295
R60 source.n2 source.n1 43.1397
R61 source.n4 source.n3 43.1397
R62 source.n6 source.n5 43.1397
R63 source.n9 source.n8 43.1397
R64 source.n11 source.n10 43.1397
R65 source.n13 source.n12 43.1397
R66 source.n26 source.n25 43.1396
R67 source.n24 source.n23 43.1396
R68 source.n22 source.n21 43.1396
R69 source.n19 source.n18 43.1396
R70 source.n17 source.n16 43.1396
R71 source.n15 source.n14 43.1396
R72 source.n15 source.n13 28.2621
R73 source.n28 source.n0 22.3138
R74 source.n28 source.n27 5.49188
R75 source.n25 source.t4 0.9905
R76 source.n25 source.t5 0.9905
R77 source.n23 source.t3 0.9905
R78 source.n23 source.t11 0.9905
R79 source.n21 source.t12 0.9905
R80 source.n21 source.t2 0.9905
R81 source.n18 source.t25 0.9905
R82 source.n18 source.t17 0.9905
R83 source.n16 source.t23 0.9905
R84 source.n16 source.t24 0.9905
R85 source.n14 source.t27 0.9905
R86 source.n14 source.t19 0.9905
R87 source.n1 source.t18 0.9905
R88 source.n1 source.t26 0.9905
R89 source.n3 source.t15 0.9905
R90 source.n3 source.t21 0.9905
R91 source.n5 source.t14 0.9905
R92 source.n5 source.t22 0.9905
R93 source.n8 source.t0 0.9905
R94 source.n8 source.t1 0.9905
R95 source.n10 source.t10 0.9905
R96 source.n10 source.t6 0.9905
R97 source.n12 source.t8 0.9905
R98 source.n12 source.t9 0.9905
R99 source.n7 source.n6 0.698776
R100 source.n22 source.n20 0.698776
R101 source.n13 source.n11 0.457397
R102 source.n11 source.n9 0.457397
R103 source.n9 source.n7 0.457397
R104 source.n6 source.n4 0.457397
R105 source.n4 source.n2 0.457397
R106 source.n2 source.n0 0.457397
R107 source.n17 source.n15 0.457397
R108 source.n19 source.n17 0.457397
R109 source.n20 source.n19 0.457397
R110 source.n24 source.n22 0.457397
R111 source.n26 source.n24 0.457397
R112 source.n27 source.n26 0.457397
R113 source source.n28 0.188
R114 drain_left.n7 drain_left.t7 61.2653
R115 drain_left.n1 drain_left.t2 61.2652
R116 drain_left.n4 drain_left.n2 60.2753
R117 drain_left.n11 drain_left.n10 59.8185
R118 drain_left.n9 drain_left.n8 59.8185
R119 drain_left.n7 drain_left.n6 59.8185
R120 drain_left.n4 drain_left.n3 59.8184
R121 drain_left.n1 drain_left.n0 59.8184
R122 drain_left drain_left.n5 36.0548
R123 drain_left drain_left.n11 6.11011
R124 drain_left.n2 drain_left.t11 0.9905
R125 drain_left.n2 drain_left.t13 0.9905
R126 drain_left.n3 drain_left.t4 0.9905
R127 drain_left.n3 drain_left.t12 0.9905
R128 drain_left.n0 drain_left.t3 0.9905
R129 drain_left.n0 drain_left.t0 0.9905
R130 drain_left.n10 drain_left.t8 0.9905
R131 drain_left.n10 drain_left.t10 0.9905
R132 drain_left.n8 drain_left.t5 0.9905
R133 drain_left.n8 drain_left.t6 0.9905
R134 drain_left.n6 drain_left.t9 0.9905
R135 drain_left.n6 drain_left.t1 0.9905
R136 drain_left.n9 drain_left.n7 0.457397
R137 drain_left.n11 drain_left.n9 0.457397
R138 drain_left.n5 drain_left.n1 0.287826
R139 drain_left.n5 drain_left.n4 0.0593781
R140 minus.n14 minus.t1 2616.31
R141 minus.n3 minus.t10 2616.31
R142 minus.n30 minus.t9 2616.31
R143 minus.n19 minus.t4 2616.31
R144 minus.n13 minus.t3 2566.65
R145 minus.n11 minus.t11 2566.65
R146 minus.n1 minus.t13 2566.65
R147 minus.n6 minus.t0 2566.65
R148 minus.n4 minus.t5 2566.65
R149 minus.n29 minus.t8 2566.65
R150 minus.n27 minus.t12 2566.65
R151 minus.n17 minus.t6 2566.65
R152 minus.n22 minus.t2 2566.65
R153 minus.n20 minus.t7 2566.65
R154 minus.n3 minus.n2 161.489
R155 minus.n19 minus.n18 161.489
R156 minus.n15 minus.n14 161.3
R157 minus.n12 minus.n0 161.3
R158 minus.n10 minus.n9 161.3
R159 minus.n8 minus.n7 161.3
R160 minus.n5 minus.n2 161.3
R161 minus.n31 minus.n30 161.3
R162 minus.n28 minus.n16 161.3
R163 minus.n26 minus.n25 161.3
R164 minus.n24 minus.n23 161.3
R165 minus.n21 minus.n18 161.3
R166 minus.n13 minus.n12 45.2793
R167 minus.n5 minus.n4 45.2793
R168 minus.n21 minus.n20 45.2793
R169 minus.n29 minus.n28 45.2793
R170 minus.n32 minus.n15 41.0668
R171 minus.n11 minus.n10 40.8975
R172 minus.n7 minus.n6 40.8975
R173 minus.n23 minus.n22 40.8975
R174 minus.n27 minus.n26 40.8975
R175 minus.n10 minus.n1 36.5157
R176 minus.n7 minus.n1 36.5157
R177 minus.n23 minus.n17 36.5157
R178 minus.n26 minus.n17 36.5157
R179 minus.n12 minus.n11 32.1338
R180 minus.n6 minus.n5 32.1338
R181 minus.n22 minus.n21 32.1338
R182 minus.n28 minus.n27 32.1338
R183 minus.n14 minus.n13 27.752
R184 minus.n4 minus.n3 27.752
R185 minus.n20 minus.n19 27.752
R186 minus.n30 minus.n29 27.752
R187 minus.n32 minus.n31 6.46073
R188 minus.n15 minus.n0 0.189894
R189 minus.n9 minus.n0 0.189894
R190 minus.n9 minus.n8 0.189894
R191 minus.n8 minus.n2 0.189894
R192 minus.n24 minus.n18 0.189894
R193 minus.n25 minus.n24 0.189894
R194 minus.n25 minus.n16 0.189894
R195 minus.n31 minus.n16 0.189894
R196 minus minus.n32 0.188
R197 drain_right.n1 drain_right.t9 61.2652
R198 drain_right.n11 drain_right.t12 60.8084
R199 drain_right.n8 drain_right.n6 60.2753
R200 drain_right.n4 drain_right.n2 60.2753
R201 drain_right.n8 drain_right.n7 59.8185
R202 drain_right.n10 drain_right.n9 59.8185
R203 drain_right.n4 drain_right.n3 59.8184
R204 drain_right.n1 drain_right.n0 59.8184
R205 drain_right drain_right.n5 35.5016
R206 drain_right drain_right.n11 5.88166
R207 drain_right.n2 drain_right.t5 0.9905
R208 drain_right.n2 drain_right.t4 0.9905
R209 drain_right.n3 drain_right.t7 0.9905
R210 drain_right.n3 drain_right.t1 0.9905
R211 drain_right.n0 drain_right.t6 0.9905
R212 drain_right.n0 drain_right.t11 0.9905
R213 drain_right.n6 drain_right.t8 0.9905
R214 drain_right.n6 drain_right.t3 0.9905
R215 drain_right.n7 drain_right.t0 0.9905
R216 drain_right.n7 drain_right.t13 0.9905
R217 drain_right.n9 drain_right.t10 0.9905
R218 drain_right.n9 drain_right.t2 0.9905
R219 drain_right.n11 drain_right.n10 0.457397
R220 drain_right.n10 drain_right.n8 0.457397
R221 drain_right.n5 drain_right.n1 0.287826
R222 drain_right.n5 drain_right.n4 0.0593781
C0 drain_left minus 0.171065f
C1 source drain_right 54.0062f
C2 source drain_left 54.025f
C3 plus drain_right 0.307632f
C4 drain_left plus 6.46827f
C5 source minus 5.54413f
C6 plus minus 6.58649f
C7 drain_left drain_right 0.79887f
C8 source plus 5.55934f
C9 drain_right minus 6.32319f
C10 drain_right a_n1564_n4888# 10.077031f
C11 drain_left a_n1564_n4888# 10.345241f
C12 source a_n1564_n4888# 8.740211f
C13 minus a_n1564_n4888# 6.592106f
C14 plus a_n1564_n4888# 9.25426f
C15 drain_right.t9 a_n1564_n4888# 6.4981f
C16 drain_right.t6 a_n1564_n4888# 0.555456f
C17 drain_right.t11 a_n1564_n4888# 0.555456f
C18 drain_right.n0 a_n1564_n4888# 5.0781f
C19 drain_right.n1 a_n1564_n4888# 0.841044f
C20 drain_right.t5 a_n1564_n4888# 0.555456f
C21 drain_right.t4 a_n1564_n4888# 0.555456f
C22 drain_right.n2 a_n1564_n4888# 5.08124f
C23 drain_right.t7 a_n1564_n4888# 0.555456f
C24 drain_right.t1 a_n1564_n4888# 0.555456f
C25 drain_right.n3 a_n1564_n4888# 5.0781f
C26 drain_right.n4 a_n1564_n4888# 0.779896f
C27 drain_right.n5 a_n1564_n4888# 2.21904f
C28 drain_right.t8 a_n1564_n4888# 0.555456f
C29 drain_right.t3 a_n1564_n4888# 0.555456f
C30 drain_right.n6 a_n1564_n4888# 5.08123f
C31 drain_right.t0 a_n1564_n4888# 0.555456f
C32 drain_right.t13 a_n1564_n4888# 0.555456f
C33 drain_right.n7 a_n1564_n4888# 5.07809f
C34 drain_right.n8 a_n1564_n4888# 0.811146f
C35 drain_right.t10 a_n1564_n4888# 0.555456f
C36 drain_right.t2 a_n1564_n4888# 0.555456f
C37 drain_right.n9 a_n1564_n4888# 5.07809f
C38 drain_right.n10 a_n1564_n4888# 0.400065f
C39 drain_right.t12 a_n1564_n4888# 6.49468f
C40 drain_right.n11 a_n1564_n4888# 0.746417f
C41 minus.n0 a_n1564_n4888# 0.055136f
C42 minus.t1 a_n1564_n4888# 0.625668f
C43 minus.t3 a_n1564_n4888# 0.621155f
C44 minus.t11 a_n1564_n4888# 0.621155f
C45 minus.t13 a_n1564_n4888# 0.621155f
C46 minus.n1 a_n1564_n4888# 0.23641f
C47 minus.n2 a_n1564_n4888# 0.123109f
C48 minus.t0 a_n1564_n4888# 0.621155f
C49 minus.t5 a_n1564_n4888# 0.621155f
C50 minus.t10 a_n1564_n4888# 0.625668f
C51 minus.n3 a_n1564_n4888# 0.252646f
C52 minus.n4 a_n1564_n4888# 0.23641f
C53 minus.n5 a_n1564_n4888# 0.01931f
C54 minus.n6 a_n1564_n4888# 0.23641f
C55 minus.n7 a_n1564_n4888# 0.01931f
C56 minus.n8 a_n1564_n4888# 0.055136f
C57 minus.n9 a_n1564_n4888# 0.055136f
C58 minus.n10 a_n1564_n4888# 0.01931f
C59 minus.n11 a_n1564_n4888# 0.23641f
C60 minus.n12 a_n1564_n4888# 0.01931f
C61 minus.n13 a_n1564_n4888# 0.23641f
C62 minus.n14 a_n1564_n4888# 0.252566f
C63 minus.n15 a_n1564_n4888# 2.36049f
C64 minus.n16 a_n1564_n4888# 0.055136f
C65 minus.t8 a_n1564_n4888# 0.621155f
C66 minus.t12 a_n1564_n4888# 0.621155f
C67 minus.t6 a_n1564_n4888# 0.621155f
C68 minus.n17 a_n1564_n4888# 0.23641f
C69 minus.n18 a_n1564_n4888# 0.123109f
C70 minus.t2 a_n1564_n4888# 0.621155f
C71 minus.t7 a_n1564_n4888# 0.621155f
C72 minus.t4 a_n1564_n4888# 0.625668f
C73 minus.n19 a_n1564_n4888# 0.252646f
C74 minus.n20 a_n1564_n4888# 0.23641f
C75 minus.n21 a_n1564_n4888# 0.01931f
C76 minus.n22 a_n1564_n4888# 0.23641f
C77 minus.n23 a_n1564_n4888# 0.01931f
C78 minus.n24 a_n1564_n4888# 0.055136f
C79 minus.n25 a_n1564_n4888# 0.055136f
C80 minus.n26 a_n1564_n4888# 0.01931f
C81 minus.n27 a_n1564_n4888# 0.23641f
C82 minus.n28 a_n1564_n4888# 0.01931f
C83 minus.n29 a_n1564_n4888# 0.23641f
C84 minus.t9 a_n1564_n4888# 0.625668f
C85 minus.n30 a_n1564_n4888# 0.252566f
C86 minus.n31 a_n1564_n4888# 0.355352f
C87 minus.n32 a_n1564_n4888# 2.8277f
C88 drain_left.t2 a_n1564_n4888# 6.50482f
C89 drain_left.t3 a_n1564_n4888# 0.55603f
C90 drain_left.t0 a_n1564_n4888# 0.55603f
C91 drain_left.n0 a_n1564_n4888# 5.08335f
C92 drain_left.n1 a_n1564_n4888# 0.841914f
C93 drain_left.t11 a_n1564_n4888# 0.55603f
C94 drain_left.t13 a_n1564_n4888# 0.55603f
C95 drain_left.n2 a_n1564_n4888# 5.08649f
C96 drain_left.t4 a_n1564_n4888# 0.55603f
C97 drain_left.t12 a_n1564_n4888# 0.55603f
C98 drain_left.n3 a_n1564_n4888# 5.08335f
C99 drain_left.n4 a_n1564_n4888# 0.780703f
C100 drain_left.n5 a_n1564_n4888# 2.29487f
C101 drain_left.t7 a_n1564_n4888# 6.50484f
C102 drain_left.t9 a_n1564_n4888# 0.55603f
C103 drain_left.t1 a_n1564_n4888# 0.55603f
C104 drain_left.n6 a_n1564_n4888# 5.08334f
C105 drain_left.n7 a_n1564_n4888# 0.85828f
C106 drain_left.t5 a_n1564_n4888# 0.55603f
C107 drain_left.t6 a_n1564_n4888# 0.55603f
C108 drain_left.n8 a_n1564_n4888# 5.08334f
C109 drain_left.n9 a_n1564_n4888# 0.400479f
C110 drain_left.t8 a_n1564_n4888# 0.55603f
C111 drain_left.t10 a_n1564_n4888# 0.55603f
C112 drain_left.n10 a_n1564_n4888# 5.08334f
C113 drain_left.n11 a_n1564_n4888# 0.688406f
C114 source.t20 a_n1564_n4888# 6.44001f
C115 source.n0 a_n1564_n4888# 2.72354f
C116 source.t18 a_n1564_n4888# 0.56351f
C117 source.t26 a_n1564_n4888# 0.56351f
C118 source.n1 a_n1564_n4888# 5.03802f
C119 source.n2 a_n1564_n4888# 0.47111f
C120 source.t15 a_n1564_n4888# 0.56351f
C121 source.t21 a_n1564_n4888# 0.56351f
C122 source.n3 a_n1564_n4888# 5.03802f
C123 source.n4 a_n1564_n4888# 0.47111f
C124 source.t14 a_n1564_n4888# 0.56351f
C125 source.t22 a_n1564_n4888# 0.56351f
C126 source.n5 a_n1564_n4888# 5.03802f
C127 source.n6 a_n1564_n4888# 0.498841f
C128 source.t7 a_n1564_n4888# 6.44002f
C129 source.n7 a_n1564_n4888# 0.633687f
C130 source.t0 a_n1564_n4888# 0.56351f
C131 source.t1 a_n1564_n4888# 0.56351f
C132 source.n8 a_n1564_n4888# 5.03802f
C133 source.n9 a_n1564_n4888# 0.47111f
C134 source.t10 a_n1564_n4888# 0.56351f
C135 source.t6 a_n1564_n4888# 0.56351f
C136 source.n10 a_n1564_n4888# 5.03802f
C137 source.n11 a_n1564_n4888# 0.47111f
C138 source.t8 a_n1564_n4888# 0.56351f
C139 source.t9 a_n1564_n4888# 0.56351f
C140 source.n12 a_n1564_n4888# 5.03802f
C141 source.n13 a_n1564_n4888# 3.26884f
C142 source.t27 a_n1564_n4888# 0.56351f
C143 source.t19 a_n1564_n4888# 0.56351f
C144 source.n14 a_n1564_n4888# 5.03803f
C145 source.n15 a_n1564_n4888# 3.26883f
C146 source.t23 a_n1564_n4888# 0.56351f
C147 source.t24 a_n1564_n4888# 0.56351f
C148 source.n16 a_n1564_n4888# 5.03803f
C149 source.n17 a_n1564_n4888# 0.4711f
C150 source.t25 a_n1564_n4888# 0.56351f
C151 source.t17 a_n1564_n4888# 0.56351f
C152 source.n18 a_n1564_n4888# 5.03803f
C153 source.n19 a_n1564_n4888# 0.4711f
C154 source.t16 a_n1564_n4888# 6.43999f
C155 source.n20 a_n1564_n4888# 0.633722f
C156 source.t12 a_n1564_n4888# 0.56351f
C157 source.t2 a_n1564_n4888# 0.56351f
C158 source.n21 a_n1564_n4888# 5.03803f
C159 source.n22 a_n1564_n4888# 0.498831f
C160 source.t3 a_n1564_n4888# 0.56351f
C161 source.t11 a_n1564_n4888# 0.56351f
C162 source.n23 a_n1564_n4888# 5.03803f
C163 source.n24 a_n1564_n4888# 0.4711f
C164 source.t4 a_n1564_n4888# 0.56351f
C165 source.t5 a_n1564_n4888# 0.56351f
C166 source.n25 a_n1564_n4888# 5.03803f
C167 source.n26 a_n1564_n4888# 0.4711f
C168 source.t13 a_n1564_n4888# 6.43999f
C169 source.n27 a_n1564_n4888# 0.800808f
C170 source.n28 a_n1564_n4888# 3.20344f
C171 plus.n0 a_n1564_n4888# 0.056376f
C172 plus.t5 a_n1564_n4888# 0.635131f
C173 plus.t7 a_n1564_n4888# 0.635131f
C174 plus.t8 a_n1564_n4888# 0.635131f
C175 plus.n1 a_n1564_n4888# 0.241729f
C176 plus.n2 a_n1564_n4888# 0.125879f
C177 plus.t12 a_n1564_n4888# 0.635131f
C178 plus.t4 a_n1564_n4888# 0.635131f
C179 plus.t6 a_n1564_n4888# 0.639745f
C180 plus.n3 a_n1564_n4888# 0.258331f
C181 plus.n4 a_n1564_n4888# 0.241729f
C182 plus.n5 a_n1564_n4888# 0.019745f
C183 plus.n6 a_n1564_n4888# 0.241729f
C184 plus.n7 a_n1564_n4888# 0.019745f
C185 plus.n8 a_n1564_n4888# 0.056376f
C186 plus.n9 a_n1564_n4888# 0.056376f
C187 plus.n10 a_n1564_n4888# 0.019745f
C188 plus.n11 a_n1564_n4888# 0.241729f
C189 plus.n12 a_n1564_n4888# 0.019745f
C190 plus.n13 a_n1564_n4888# 0.241729f
C191 plus.t3 a_n1564_n4888# 0.639745f
C192 plus.n14 a_n1564_n4888# 0.258249f
C193 plus.n15 a_n1564_n4888# 0.850939f
C194 plus.n16 a_n1564_n4888# 0.056376f
C195 plus.t11 a_n1564_n4888# 0.639745f
C196 plus.t10 a_n1564_n4888# 0.635131f
C197 plus.t13 a_n1564_n4888# 0.635131f
C198 plus.t9 a_n1564_n4888# 0.635131f
C199 plus.n17 a_n1564_n4888# 0.241729f
C200 plus.n18 a_n1564_n4888# 0.125879f
C201 plus.t1 a_n1564_n4888# 0.635131f
C202 plus.t2 a_n1564_n4888# 0.635131f
C203 plus.t0 a_n1564_n4888# 0.639745f
C204 plus.n19 a_n1564_n4888# 0.258331f
C205 plus.n20 a_n1564_n4888# 0.241729f
C206 plus.n21 a_n1564_n4888# 0.019745f
C207 plus.n22 a_n1564_n4888# 0.241729f
C208 plus.n23 a_n1564_n4888# 0.019745f
C209 plus.n24 a_n1564_n4888# 0.056376f
C210 plus.n25 a_n1564_n4888# 0.056376f
C211 plus.n26 a_n1564_n4888# 0.019745f
C212 plus.n27 a_n1564_n4888# 0.241729f
C213 plus.n28 a_n1564_n4888# 0.019745f
C214 plus.n29 a_n1564_n4888# 0.241729f
C215 plus.n30 a_n1564_n4888# 0.258249f
C216 plus.n31 a_n1564_n4888# 1.90032f
.ends

