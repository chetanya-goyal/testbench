* NGSPICE file created from diffpair343.ext - technology: sky130A

.subckt diffpair343 minus drain_right drain_left source plus
X0 a_n1296_n2688# a_n1296_n2688# a_n1296_n2688# a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.25
X1 drain_left.t7 plus.t0 source.t8 a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X2 drain_left.t6 plus.t1 source.t4 a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X3 drain_right.t7 minus.t0 source.t12 a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X4 a_n1296_n2688# a_n1296_n2688# a_n1296_n2688# a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
X5 source.t0 minus.t1 drain_right.t6 a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X6 source.t15 minus.t2 drain_right.t5 a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X7 drain_left.t5 plus.t2 source.t11 a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X8 source.t10 plus.t3 drain_left.t4 a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X9 a_n1296_n2688# a_n1296_n2688# a_n1296_n2688# a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
X10 source.t9 plus.t4 drain_left.t3 a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X11 drain_right.t4 minus.t3 source.t2 a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X12 source.t6 plus.t5 drain_left.t2 a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X13 drain_right.t3 minus.t4 source.t1 a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X14 source.t13 minus.t5 drain_right.t2 a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X15 drain_right.t1 minus.t6 source.t14 a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X16 drain_left.t1 plus.t6 source.t5 a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X17 source.t3 minus.t7 drain_right.t0 a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X18 source.t7 plus.t7 drain_left.t0 a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X19 a_n1296_n2688# a_n1296_n2688# a_n1296_n2688# a_n1296_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
R0 plus.n1 plus.t3 1046.96
R1 plus.n5 plus.t0 1046.96
R2 plus.n8 plus.t6 1046.96
R3 plus.n12 plus.t7 1046.96
R4 plus.n2 plus.t1 992.92
R5 plus.n4 plus.t4 992.92
R6 plus.n9 plus.t5 992.92
R7 plus.n11 plus.t2 992.92
R8 plus.n1 plus.n0 161.489
R9 plus.n8 plus.n7 161.489
R10 plus.n3 plus.n0 161.3
R11 plus.n6 plus.n5 161.3
R12 plus.n10 plus.n7 161.3
R13 plus.n13 plus.n12 161.3
R14 plus.n3 plus.n2 42.3581
R15 plus.n4 plus.n3 42.3581
R16 plus.n11 plus.n10 42.3581
R17 plus.n10 plus.n9 42.3581
R18 plus.n2 plus.n1 30.6732
R19 plus.n5 plus.n4 30.6732
R20 plus.n12 plus.n11 30.6732
R21 plus.n9 plus.n8 30.6732
R22 plus plus.n13 26.7755
R23 plus plus.n6 11.0081
R24 plus.n6 plus.n0 0.189894
R25 plus.n13 plus.n7 0.189894
R26 source.n3 source.t10 51.0588
R27 source.n4 source.t14 51.0588
R28 source.n7 source.t0 51.0588
R29 source.n15 source.t2 51.0586
R30 source.n12 source.t3 51.0586
R31 source.n11 source.t5 51.0586
R32 source.n8 source.t7 51.0586
R33 source.n0 source.t8 51.0586
R34 source.n2 source.n1 48.8588
R35 source.n6 source.n5 48.8588
R36 source.n14 source.n13 48.8586
R37 source.n10 source.n9 48.8586
R38 source.n8 source.n7 19.515
R39 source.n16 source.n0 14.0021
R40 source.n16 source.n15 5.51343
R41 source.n13 source.t12 2.2005
R42 source.n13 source.t13 2.2005
R43 source.n9 source.t11 2.2005
R44 source.n9 source.t6 2.2005
R45 source.n1 source.t4 2.2005
R46 source.n1 source.t9 2.2005
R47 source.n5 source.t1 2.2005
R48 source.n5 source.t15 2.2005
R49 source.n7 source.n6 0.5005
R50 source.n6 source.n4 0.5005
R51 source.n3 source.n2 0.5005
R52 source.n2 source.n0 0.5005
R53 source.n10 source.n8 0.5005
R54 source.n11 source.n10 0.5005
R55 source.n14 source.n12 0.5005
R56 source.n15 source.n14 0.5005
R57 source.n4 source.n3 0.470328
R58 source.n12 source.n11 0.470328
R59 source source.n16 0.188
R60 drain_left.n5 drain_left.n3 66.0376
R61 drain_left.n2 drain_left.n1 65.732
R62 drain_left.n2 drain_left.n0 65.732
R63 drain_left.n5 drain_left.n4 65.5374
R64 drain_left drain_left.n2 26.8443
R65 drain_left drain_left.n5 6.15322
R66 drain_left.n1 drain_left.t2 2.2005
R67 drain_left.n1 drain_left.t1 2.2005
R68 drain_left.n0 drain_left.t0 2.2005
R69 drain_left.n0 drain_left.t5 2.2005
R70 drain_left.n4 drain_left.t3 2.2005
R71 drain_left.n4 drain_left.t7 2.2005
R72 drain_left.n3 drain_left.t4 2.2005
R73 drain_left.n3 drain_left.t6 2.2005
R74 minus.n5 minus.t1 1046.96
R75 minus.n1 minus.t6 1046.96
R76 minus.n12 minus.t3 1046.96
R77 minus.n8 minus.t7 1046.96
R78 minus.n4 minus.t4 992.92
R79 minus.n2 minus.t2 992.92
R80 minus.n11 minus.t5 992.92
R81 minus.n9 minus.t0 992.92
R82 minus.n1 minus.n0 161.489
R83 minus.n8 minus.n7 161.489
R84 minus.n6 minus.n5 161.3
R85 minus.n3 minus.n0 161.3
R86 minus.n13 minus.n12 161.3
R87 minus.n10 minus.n7 161.3
R88 minus.n4 minus.n3 42.3581
R89 minus.n3 minus.n2 42.3581
R90 minus.n10 minus.n9 42.3581
R91 minus.n11 minus.n10 42.3581
R92 minus.n14 minus.n6 31.7581
R93 minus.n5 minus.n4 30.6732
R94 minus.n2 minus.n1 30.6732
R95 minus.n9 minus.n8 30.6732
R96 minus.n12 minus.n11 30.6732
R97 minus.n14 minus.n13 6.5005
R98 minus.n6 minus.n0 0.189894
R99 minus.n13 minus.n7 0.189894
R100 minus minus.n14 0.188
R101 drain_right.n5 drain_right.n3 66.0374
R102 drain_right.n2 drain_right.n1 65.732
R103 drain_right.n2 drain_right.n0 65.732
R104 drain_right.n5 drain_right.n4 65.5376
R105 drain_right drain_right.n2 26.2911
R106 drain_right drain_right.n5 6.15322
R107 drain_right.n1 drain_right.t2 2.2005
R108 drain_right.n1 drain_right.t4 2.2005
R109 drain_right.n0 drain_right.t0 2.2005
R110 drain_right.n0 drain_right.t7 2.2005
R111 drain_right.n3 drain_right.t5 2.2005
R112 drain_right.n3 drain_right.t1 2.2005
R113 drain_right.n4 drain_right.t6 2.2005
R114 drain_right.n4 drain_right.t3 2.2005
C0 source minus 2.00805f
C1 minus plus 4.21057f
C2 drain_right drain_left 0.605638f
C3 drain_right source 13.8981f
C4 drain_right plus 0.275273f
C5 drain_right minus 2.33765f
C6 source drain_left 13.899199f
C7 drain_left plus 2.45965f
C8 drain_left minus 0.170438f
C9 source plus 2.02209f
C10 drain_right a_n1296_n2688# 5.15236f
C11 drain_left a_n1296_n2688# 5.36262f
C12 source a_n1296_n2688# 6.819076f
C13 minus a_n1296_n2688# 4.776173f
C14 plus a_n1296_n2688# 6.60713f
C15 drain_right.t0 a_n1296_n2688# 0.244388f
C16 drain_right.t7 a_n1296_n2688# 0.244388f
C17 drain_right.n0 a_n1296_n2688# 2.13868f
C18 drain_right.t2 a_n1296_n2688# 0.244388f
C19 drain_right.t4 a_n1296_n2688# 0.244388f
C20 drain_right.n1 a_n1296_n2688# 2.13868f
C21 drain_right.n2 a_n1296_n2688# 1.91795f
C22 drain_right.t5 a_n1296_n2688# 0.244388f
C23 drain_right.t1 a_n1296_n2688# 0.244388f
C24 drain_right.n3 a_n1296_n2688# 2.1406f
C25 drain_right.t6 a_n1296_n2688# 0.244388f
C26 drain_right.t3 a_n1296_n2688# 0.244388f
C27 drain_right.n4 a_n1296_n2688# 2.13759f
C28 drain_right.n5 a_n1296_n2688# 1.06639f
C29 minus.n0 a_n1296_n2688# 0.129565f
C30 minus.t1 a_n1296_n2688# 0.367168f
C31 minus.t4 a_n1296_n2688# 0.359064f
C32 minus.t2 a_n1296_n2688# 0.359064f
C33 minus.t6 a_n1296_n2688# 0.367168f
C34 minus.n1 a_n1296_n2688# 0.170441f
C35 minus.n2 a_n1296_n2688# 0.152832f
C36 minus.n3 a_n1296_n2688# 0.021461f
C37 minus.n4 a_n1296_n2688# 0.152832f
C38 minus.n5 a_n1296_n2688# 0.170355f
C39 minus.n6 a_n1296_n2688# 1.61251f
C40 minus.n7 a_n1296_n2688# 0.129565f
C41 minus.t5 a_n1296_n2688# 0.359064f
C42 minus.t0 a_n1296_n2688# 0.359064f
C43 minus.t7 a_n1296_n2688# 0.367168f
C44 minus.n8 a_n1296_n2688# 0.170441f
C45 minus.n9 a_n1296_n2688# 0.152832f
C46 minus.n10 a_n1296_n2688# 0.021461f
C47 minus.n11 a_n1296_n2688# 0.152832f
C48 minus.t3 a_n1296_n2688# 0.367168f
C49 minus.n12 a_n1296_n2688# 0.170355f
C50 minus.n13 a_n1296_n2688# 0.368261f
C51 minus.n14 a_n1296_n2688# 1.98234f
C52 drain_left.t0 a_n1296_n2688# 0.245369f
C53 drain_left.t5 a_n1296_n2688# 0.245369f
C54 drain_left.n0 a_n1296_n2688# 2.14726f
C55 drain_left.t2 a_n1296_n2688# 0.245369f
C56 drain_left.t1 a_n1296_n2688# 0.245369f
C57 drain_left.n1 a_n1296_n2688# 2.14726f
C58 drain_left.n2 a_n1296_n2688# 1.9974f
C59 drain_left.t4 a_n1296_n2688# 0.245369f
C60 drain_left.t6 a_n1296_n2688# 0.245369f
C61 drain_left.n3 a_n1296_n2688# 2.14921f
C62 drain_left.t3 a_n1296_n2688# 0.245369f
C63 drain_left.t7 a_n1296_n2688# 0.245369f
C64 drain_left.n4 a_n1296_n2688# 2.14616f
C65 drain_left.n5 a_n1296_n2688# 1.07068f
C66 source.t8 a_n1296_n2688# 1.93255f
C67 source.n0 a_n1296_n2688# 1.10534f
C68 source.t4 a_n1296_n2688# 0.181231f
C69 source.t9 a_n1296_n2688# 0.181231f
C70 source.n1 a_n1296_n2688# 1.51715f
C71 source.n2 a_n1296_n2688# 0.319607f
C72 source.t10 a_n1296_n2688# 1.93255f
C73 source.n3 a_n1296_n2688# 0.395988f
C74 source.t14 a_n1296_n2688# 1.93255f
C75 source.n4 a_n1296_n2688# 0.395988f
C76 source.t1 a_n1296_n2688# 0.181231f
C77 source.t15 a_n1296_n2688# 0.181231f
C78 source.n5 a_n1296_n2688# 1.51715f
C79 source.n6 a_n1296_n2688# 0.319607f
C80 source.t0 a_n1296_n2688# 1.93255f
C81 source.n7 a_n1296_n2688# 1.47444f
C82 source.t7 a_n1296_n2688# 1.93255f
C83 source.n8 a_n1296_n2688# 1.47444f
C84 source.t11 a_n1296_n2688# 0.181231f
C85 source.t6 a_n1296_n2688# 0.181231f
C86 source.n9 a_n1296_n2688# 1.51714f
C87 source.n10 a_n1296_n2688# 0.319611f
C88 source.t5 a_n1296_n2688# 1.93255f
C89 source.n11 a_n1296_n2688# 0.395993f
C90 source.t3 a_n1296_n2688# 1.93255f
C91 source.n12 a_n1296_n2688# 0.395993f
C92 source.t12 a_n1296_n2688# 0.181231f
C93 source.t13 a_n1296_n2688# 0.181231f
C94 source.n13 a_n1296_n2688# 1.51714f
C95 source.n14 a_n1296_n2688# 0.319611f
C96 source.t2 a_n1296_n2688# 1.93255f
C97 source.n15 a_n1296_n2688# 0.537006f
C98 source.n16 a_n1296_n2688# 1.32467f
C99 plus.n0 a_n1296_n2688# 0.134414f
C100 plus.t4 a_n1296_n2688# 0.372503f
C101 plus.t1 a_n1296_n2688# 0.372503f
C102 plus.t3 a_n1296_n2688# 0.380911f
C103 plus.n1 a_n1296_n2688# 0.176821f
C104 plus.n2 a_n1296_n2688# 0.158553f
C105 plus.n3 a_n1296_n2688# 0.022264f
C106 plus.n4 a_n1296_n2688# 0.158553f
C107 plus.t0 a_n1296_n2688# 0.380911f
C108 plus.n5 a_n1296_n2688# 0.176732f
C109 plus.n6 a_n1296_n2688# 0.573991f
C110 plus.n7 a_n1296_n2688# 0.134414f
C111 plus.t7 a_n1296_n2688# 0.380911f
C112 plus.t2 a_n1296_n2688# 0.372503f
C113 plus.t5 a_n1296_n2688# 0.372503f
C114 plus.t6 a_n1296_n2688# 0.380911f
C115 plus.n8 a_n1296_n2688# 0.176821f
C116 plus.n9 a_n1296_n2688# 0.158553f
C117 plus.n10 a_n1296_n2688# 0.022264f
C118 plus.n11 a_n1296_n2688# 0.158553f
C119 plus.n12 a_n1296_n2688# 0.176732f
C120 plus.n13 a_n1296_n2688# 1.45671f
.ends

