* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t16 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X1 drain_left.t18 plus.t1 source.t14 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X2 source.t4 minus.t0 drain_right.t19 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X3 drain_right.t18 minus.t1 source.t3 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X4 drain_right.t17 minus.t2 source.t8 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X5 drain_right.t16 minus.t3 source.t6 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X6 a_n2102_n1088# a_n2102_n1088# a_n2102_n1088# a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.3
X7 source.t5 minus.t4 drain_right.t15 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X8 source.t22 plus.t2 drain_left.t17 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X9 source.t31 plus.t3 drain_left.t16 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X10 source.t32 plus.t4 drain_left.t15 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X11 source.t7 minus.t5 drain_right.t14 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X12 drain_right.t13 minus.t6 source.t2 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X13 drain_right.t12 minus.t7 source.t1 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X14 drain_left.t14 plus.t5 source.t20 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X15 drain_left.t13 plus.t6 source.t24 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X16 drain_right.t11 minus.t8 source.t0 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X17 source.t34 minus.t9 drain_right.t10 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X18 a_n2102_n1088# a_n2102_n1088# a_n2102_n1088# a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X19 source.t39 minus.t10 drain_right.t9 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X20 source.t25 plus.t7 drain_left.t12 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X21 source.t21 plus.t8 drain_left.t11 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X22 drain_left.t10 plus.t9 source.t23 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X23 drain_left.t9 plus.t10 source.t29 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X24 source.t37 minus.t11 drain_right.t8 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X25 a_n2102_n1088# a_n2102_n1088# a_n2102_n1088# a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X26 source.t17 plus.t11 drain_left.t8 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X27 drain_right.t7 minus.t12 source.t33 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X28 source.t12 minus.t13 drain_right.t6 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X29 drain_left.t7 plus.t12 source.t19 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X30 source.t30 plus.t13 drain_left.t6 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X31 source.t18 plus.t14 drain_left.t5 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X32 drain_right.t5 minus.t14 source.t11 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X33 drain_left.t4 plus.t15 source.t27 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X34 drain_left.t3 plus.t16 source.t28 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X35 drain_right.t4 minus.t15 source.t38 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X36 drain_right.t3 minus.t16 source.t36 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X37 source.t35 minus.t17 drain_right.t2 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X38 source.t9 minus.t18 drain_right.t1 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X39 source.t10 minus.t19 drain_right.t0 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X40 source.t15 plus.t17 drain_left.t2 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X41 source.t13 plus.t18 drain_left.t1 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X42 drain_left.t0 plus.t19 source.t26 a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X43 a_n2102_n1088# a_n2102_n1088# a_n2102_n1088# a_n2102_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
R0 plus.n6 plus.t4 233.697
R1 plus.n27 plus.t16 233.697
R2 plus.n36 plus.t10 233.697
R3 plus.n56 plus.t17 233.697
R4 plus.n5 plus.t9 184.768
R5 plus.n9 plus.t14 184.768
R6 plus.n3 plus.t19 184.768
R7 plus.n15 plus.t8 184.768
R8 plus.n17 plus.t12 184.768
R9 plus.n18 plus.t18 184.768
R10 plus.n24 plus.t1 184.768
R11 plus.n26 plus.t11 184.768
R12 plus.n35 plus.t2 184.768
R13 plus.n39 plus.t0 184.768
R14 plus.n33 plus.t13 184.768
R15 plus.n45 plus.t5 184.768
R16 plus.n47 plus.t3 184.768
R17 plus.n32 plus.t15 184.768
R18 plus.n53 plus.t7 184.768
R19 plus.n55 plus.t6 184.768
R20 plus.n7 plus.n6 161.489
R21 plus.n37 plus.n36 161.489
R22 plus.n8 plus.n7 161.3
R23 plus.n10 plus.n4 161.3
R24 plus.n12 plus.n11 161.3
R25 plus.n14 plus.n13 161.3
R26 plus.n16 plus.n2 161.3
R27 plus.n20 plus.n19 161.3
R28 plus.n21 plus.n1 161.3
R29 plus.n23 plus.n22 161.3
R30 plus.n25 plus.n0 161.3
R31 plus.n28 plus.n27 161.3
R32 plus.n38 plus.n37 161.3
R33 plus.n40 plus.n34 161.3
R34 plus.n42 plus.n41 161.3
R35 plus.n44 plus.n43 161.3
R36 plus.n46 plus.n31 161.3
R37 plus.n49 plus.n48 161.3
R38 plus.n50 plus.n30 161.3
R39 plus.n52 plus.n51 161.3
R40 plus.n54 plus.n29 161.3
R41 plus.n57 plus.n56 161.3
R42 plus.n11 plus.n10 73.0308
R43 plus.n23 plus.n1 73.0308
R44 plus.n52 plus.n30 73.0308
R45 plus.n41 plus.n40 73.0308
R46 plus.n14 plus.n3 64.9975
R47 plus.n19 plus.n18 64.9975
R48 plus.n48 plus.n32 64.9975
R49 plus.n44 plus.n33 64.9975
R50 plus.n9 plus.n8 62.0763
R51 plus.n25 plus.n24 62.0763
R52 plus.n54 plus.n53 62.0763
R53 plus.n39 plus.n38 62.0763
R54 plus.n16 plus.n15 46.0096
R55 plus.n17 plus.n16 46.0096
R56 plus.n47 plus.n46 46.0096
R57 plus.n46 plus.n45 46.0096
R58 plus.n6 plus.n5 43.0884
R59 plus.n27 plus.n26 43.0884
R60 plus.n56 plus.n55 43.0884
R61 plus.n36 plus.n35 43.0884
R62 plus.n8 plus.n5 29.9429
R63 plus.n26 plus.n25 29.9429
R64 plus.n55 plus.n54 29.9429
R65 plus.n38 plus.n35 29.9429
R66 plus.n15 plus.n14 27.0217
R67 plus.n19 plus.n17 27.0217
R68 plus.n48 plus.n47 27.0217
R69 plus.n45 plus.n44 27.0217
R70 plus plus.n57 26.8134
R71 plus.n10 plus.n9 10.955
R72 plus.n24 plus.n23 10.955
R73 plus.n53 plus.n52 10.955
R74 plus.n40 plus.n39 10.955
R75 plus.n11 plus.n3 8.03383
R76 plus.n18 plus.n1 8.03383
R77 plus.n32 plus.n30 8.03383
R78 plus.n41 plus.n33 8.03383
R79 plus plus.n28 7.99292
R80 plus.n7 plus.n4 0.189894
R81 plus.n12 plus.n4 0.189894
R82 plus.n13 plus.n12 0.189894
R83 plus.n13 plus.n2 0.189894
R84 plus.n20 plus.n2 0.189894
R85 plus.n21 plus.n20 0.189894
R86 plus.n22 plus.n21 0.189894
R87 plus.n22 plus.n0 0.189894
R88 plus.n28 plus.n0 0.189894
R89 plus.n57 plus.n29 0.189894
R90 plus.n51 plus.n29 0.189894
R91 plus.n51 plus.n50 0.189894
R92 plus.n50 plus.n49 0.189894
R93 plus.n49 plus.n31 0.189894
R94 plus.n43 plus.n31 0.189894
R95 plus.n43 plus.n42 0.189894
R96 plus.n42 plus.n34 0.189894
R97 plus.n37 plus.n34 0.189894
R98 source.n0 source.t28 243.255
R99 source.n9 source.t32 243.255
R100 source.n10 source.t33 243.255
R101 source.n19 source.t34 243.255
R102 source.n39 source.t6 243.254
R103 source.n30 source.t12 243.254
R104 source.n29 source.t29 243.254
R105 source.n20 source.t15 243.254
R106 source.n2 source.n1 223.454
R107 source.n4 source.n3 223.454
R108 source.n6 source.n5 223.454
R109 source.n8 source.n7 223.454
R110 source.n12 source.n11 223.454
R111 source.n14 source.n13 223.454
R112 source.n16 source.n15 223.454
R113 source.n18 source.n17 223.454
R114 source.n38 source.n37 223.453
R115 source.n36 source.n35 223.453
R116 source.n34 source.n33 223.453
R117 source.n32 source.n31 223.453
R118 source.n28 source.n27 223.453
R119 source.n26 source.n25 223.453
R120 source.n24 source.n23 223.453
R121 source.n22 source.n21 223.453
R122 source.n37 source.t36 19.8005
R123 source.n37 source.t7 19.8005
R124 source.n35 source.t1 19.8005
R125 source.n35 source.t10 19.8005
R126 source.n33 source.t11 19.8005
R127 source.n33 source.t39 19.8005
R128 source.n31 source.t2 19.8005
R129 source.n31 source.t5 19.8005
R130 source.n27 source.t16 19.8005
R131 source.n27 source.t22 19.8005
R132 source.n25 source.t20 19.8005
R133 source.n25 source.t30 19.8005
R134 source.n23 source.t27 19.8005
R135 source.n23 source.t31 19.8005
R136 source.n21 source.t24 19.8005
R137 source.n21 source.t25 19.8005
R138 source.n1 source.t14 19.8005
R139 source.n1 source.t17 19.8005
R140 source.n3 source.t19 19.8005
R141 source.n3 source.t13 19.8005
R142 source.n5 source.t26 19.8005
R143 source.n5 source.t21 19.8005
R144 source.n7 source.t23 19.8005
R145 source.n7 source.t18 19.8005
R146 source.n11 source.t3 19.8005
R147 source.n11 source.t35 19.8005
R148 source.n13 source.t38 19.8005
R149 source.n13 source.t37 19.8005
R150 source.n15 source.t0 19.8005
R151 source.n15 source.t4 19.8005
R152 source.n17 source.t8 19.8005
R153 source.n17 source.t9 19.8005
R154 source.n20 source.n19 13.4975
R155 source.n40 source.n0 7.96301
R156 source.n40 source.n39 5.53498
R157 source.n19 source.n18 0.543603
R158 source.n18 source.n16 0.543603
R159 source.n16 source.n14 0.543603
R160 source.n14 source.n12 0.543603
R161 source.n12 source.n10 0.543603
R162 source.n9 source.n8 0.543603
R163 source.n8 source.n6 0.543603
R164 source.n6 source.n4 0.543603
R165 source.n4 source.n2 0.543603
R166 source.n2 source.n0 0.543603
R167 source.n22 source.n20 0.543603
R168 source.n24 source.n22 0.543603
R169 source.n26 source.n24 0.543603
R170 source.n28 source.n26 0.543603
R171 source.n29 source.n28 0.543603
R172 source.n32 source.n30 0.543603
R173 source.n34 source.n32 0.543603
R174 source.n36 source.n34 0.543603
R175 source.n38 source.n36 0.543603
R176 source.n39 source.n38 0.543603
R177 source.n10 source.n9 0.470328
R178 source.n30 source.n29 0.470328
R179 source source.n40 0.188
R180 drain_left.n10 drain_left.n8 240.675
R181 drain_left.n6 drain_left.n4 240.674
R182 drain_left.n2 drain_left.n0 240.674
R183 drain_left.n16 drain_left.n15 240.132
R184 drain_left.n14 drain_left.n13 240.132
R185 drain_left.n12 drain_left.n11 240.132
R186 drain_left.n10 drain_left.n9 240.132
R187 drain_left.n7 drain_left.n3 240.131
R188 drain_left.n6 drain_left.n5 240.131
R189 drain_left.n2 drain_left.n1 240.131
R190 drain_left drain_left.n7 23.3786
R191 drain_left.n3 drain_left.t16 19.8005
R192 drain_left.n3 drain_left.t14 19.8005
R193 drain_left.n4 drain_left.t17 19.8005
R194 drain_left.n4 drain_left.t9 19.8005
R195 drain_left.n5 drain_left.t6 19.8005
R196 drain_left.n5 drain_left.t19 19.8005
R197 drain_left.n1 drain_left.t12 19.8005
R198 drain_left.n1 drain_left.t4 19.8005
R199 drain_left.n0 drain_left.t2 19.8005
R200 drain_left.n0 drain_left.t13 19.8005
R201 drain_left.n15 drain_left.t8 19.8005
R202 drain_left.n15 drain_left.t3 19.8005
R203 drain_left.n13 drain_left.t1 19.8005
R204 drain_left.n13 drain_left.t18 19.8005
R205 drain_left.n11 drain_left.t11 19.8005
R206 drain_left.n11 drain_left.t7 19.8005
R207 drain_left.n9 drain_left.t5 19.8005
R208 drain_left.n9 drain_left.t0 19.8005
R209 drain_left.n8 drain_left.t15 19.8005
R210 drain_left.n8 drain_left.t10 19.8005
R211 drain_left drain_left.n16 6.19632
R212 drain_left.n12 drain_left.n10 0.543603
R213 drain_left.n14 drain_left.n12 0.543603
R214 drain_left.n16 drain_left.n14 0.543603
R215 drain_left.n7 drain_left.n6 0.488257
R216 drain_left.n7 drain_left.n2 0.488257
R217 minus.n27 minus.t9 233.697
R218 minus.n7 minus.t12 233.697
R219 minus.n56 minus.t3 233.697
R220 minus.n35 minus.t13 233.697
R221 minus.n26 minus.t2 184.768
R222 minus.n24 minus.t18 184.768
R223 minus.n3 minus.t8 184.768
R224 minus.n18 minus.t0 184.768
R225 minus.n16 minus.t15 184.768
R226 minus.n4 minus.t11 184.768
R227 minus.n10 minus.t1 184.768
R228 minus.n6 minus.t17 184.768
R229 minus.n55 minus.t5 184.768
R230 minus.n53 minus.t16 184.768
R231 minus.n47 minus.t19 184.768
R232 minus.n46 minus.t7 184.768
R233 minus.n44 minus.t10 184.768
R234 minus.n32 minus.t14 184.768
R235 minus.n38 minus.t4 184.768
R236 minus.n34 minus.t6 184.768
R237 minus.n8 minus.n7 161.489
R238 minus.n36 minus.n35 161.489
R239 minus.n28 minus.n27 161.3
R240 minus.n25 minus.n0 161.3
R241 minus.n23 minus.n22 161.3
R242 minus.n21 minus.n1 161.3
R243 minus.n20 minus.n19 161.3
R244 minus.n17 minus.n2 161.3
R245 minus.n15 minus.n14 161.3
R246 minus.n13 minus.n12 161.3
R247 minus.n11 minus.n5 161.3
R248 minus.n9 minus.n8 161.3
R249 minus.n57 minus.n56 161.3
R250 minus.n54 minus.n29 161.3
R251 minus.n52 minus.n51 161.3
R252 minus.n50 minus.n30 161.3
R253 minus.n49 minus.n48 161.3
R254 minus.n45 minus.n31 161.3
R255 minus.n43 minus.n42 161.3
R256 minus.n41 minus.n40 161.3
R257 minus.n39 minus.n33 161.3
R258 minus.n37 minus.n36 161.3
R259 minus.n23 minus.n1 73.0308
R260 minus.n12 minus.n11 73.0308
R261 minus.n40 minus.n39 73.0308
R262 minus.n52 minus.n30 73.0308
R263 minus.n19 minus.n3 64.9975
R264 minus.n15 minus.n4 64.9975
R265 minus.n43 minus.n32 64.9975
R266 minus.n48 minus.n47 64.9975
R267 minus.n25 minus.n24 62.0763
R268 minus.n10 minus.n9 62.0763
R269 minus.n38 minus.n37 62.0763
R270 minus.n54 minus.n53 62.0763
R271 minus.n18 minus.n17 46.0096
R272 minus.n17 minus.n16 46.0096
R273 minus.n45 minus.n44 46.0096
R274 minus.n46 minus.n45 46.0096
R275 minus.n27 minus.n26 43.0884
R276 minus.n7 minus.n6 43.0884
R277 minus.n35 minus.n34 43.0884
R278 minus.n56 minus.n55 43.0884
R279 minus.n26 minus.n25 29.9429
R280 minus.n9 minus.n6 29.9429
R281 minus.n37 minus.n34 29.9429
R282 minus.n55 minus.n54 29.9429
R283 minus.n58 minus.n28 28.7657
R284 minus.n19 minus.n18 27.0217
R285 minus.n16 minus.n15 27.0217
R286 minus.n44 minus.n43 27.0217
R287 minus.n48 minus.n46 27.0217
R288 minus.n24 minus.n23 10.955
R289 minus.n11 minus.n10 10.955
R290 minus.n39 minus.n38 10.955
R291 minus.n53 minus.n52 10.955
R292 minus.n3 minus.n1 8.03383
R293 minus.n12 minus.n4 8.03383
R294 minus.n40 minus.n32 8.03383
R295 minus.n47 minus.n30 8.03383
R296 minus.n58 minus.n57 6.51565
R297 minus.n28 minus.n0 0.189894
R298 minus.n22 minus.n0 0.189894
R299 minus.n22 minus.n21 0.189894
R300 minus.n21 minus.n20 0.189894
R301 minus.n20 minus.n2 0.189894
R302 minus.n14 minus.n2 0.189894
R303 minus.n14 minus.n13 0.189894
R304 minus.n13 minus.n5 0.189894
R305 minus.n8 minus.n5 0.189894
R306 minus.n36 minus.n33 0.189894
R307 minus.n41 minus.n33 0.189894
R308 minus.n42 minus.n41 0.189894
R309 minus.n42 minus.n31 0.189894
R310 minus.n49 minus.n31 0.189894
R311 minus.n50 minus.n49 0.189894
R312 minus.n51 minus.n50 0.189894
R313 minus.n51 minus.n29 0.189894
R314 minus.n57 minus.n29 0.189894
R315 minus minus.n58 0.188
R316 drain_right.n10 drain_right.n8 240.675
R317 drain_right.n6 drain_right.n4 240.674
R318 drain_right.n2 drain_right.n0 240.674
R319 drain_right.n10 drain_right.n9 240.132
R320 drain_right.n12 drain_right.n11 240.132
R321 drain_right.n14 drain_right.n13 240.132
R322 drain_right.n16 drain_right.n15 240.132
R323 drain_right.n7 drain_right.n3 240.131
R324 drain_right.n6 drain_right.n5 240.131
R325 drain_right.n2 drain_right.n1 240.131
R326 drain_right drain_right.n7 22.8253
R327 drain_right.n3 drain_right.t9 19.8005
R328 drain_right.n3 drain_right.t12 19.8005
R329 drain_right.n4 drain_right.t14 19.8005
R330 drain_right.n4 drain_right.t16 19.8005
R331 drain_right.n5 drain_right.t0 19.8005
R332 drain_right.n5 drain_right.t3 19.8005
R333 drain_right.n1 drain_right.t15 19.8005
R334 drain_right.n1 drain_right.t5 19.8005
R335 drain_right.n0 drain_right.t6 19.8005
R336 drain_right.n0 drain_right.t13 19.8005
R337 drain_right.n8 drain_right.t2 19.8005
R338 drain_right.n8 drain_right.t7 19.8005
R339 drain_right.n9 drain_right.t8 19.8005
R340 drain_right.n9 drain_right.t18 19.8005
R341 drain_right.n11 drain_right.t19 19.8005
R342 drain_right.n11 drain_right.t4 19.8005
R343 drain_right.n13 drain_right.t1 19.8005
R344 drain_right.n13 drain_right.t11 19.8005
R345 drain_right.n15 drain_right.t10 19.8005
R346 drain_right.n15 drain_right.t17 19.8005
R347 drain_right drain_right.n16 6.19632
R348 drain_right.n16 drain_right.n14 0.543603
R349 drain_right.n14 drain_right.n12 0.543603
R350 drain_right.n12 drain_right.n10 0.543603
R351 drain_right.n7 drain_right.n6 0.488257
R352 drain_right.n7 drain_right.n2 0.488257
C0 drain_right source 6.15332f
C1 drain_left plus 1.35853f
C2 drain_left minus 0.179105f
C3 plus minus 3.74723f
C4 drain_left source 6.1529f
C5 plus source 1.52861f
C6 minus source 1.51475f
C7 drain_left drain_right 1.10881f
C8 drain_right plus 0.3693f
C9 drain_right minus 1.15266f
C10 drain_right a_n2102_n1088# 4.06542f
C11 drain_left a_n2102_n1088# 4.34638f
C12 source a_n2102_n1088# 2.645866f
C13 minus a_n2102_n1088# 7.337873f
C14 plus a_n2102_n1088# 7.987417f
C15 drain_right.t6 a_n2102_n1088# 0.020541f
C16 drain_right.t13 a_n2102_n1088# 0.020541f
C17 drain_right.n0 a_n2102_n1088# 0.080455f
C18 drain_right.t15 a_n2102_n1088# 0.020541f
C19 drain_right.t5 a_n2102_n1088# 0.020541f
C20 drain_right.n1 a_n2102_n1088# 0.079816f
C21 drain_right.n2 a_n2102_n1088# 0.55194f
C22 drain_right.t9 a_n2102_n1088# 0.020541f
C23 drain_right.t12 a_n2102_n1088# 0.020541f
C24 drain_right.n3 a_n2102_n1088# 0.079816f
C25 drain_right.t14 a_n2102_n1088# 0.020541f
C26 drain_right.t16 a_n2102_n1088# 0.020541f
C27 drain_right.n4 a_n2102_n1088# 0.080455f
C28 drain_right.t0 a_n2102_n1088# 0.020541f
C29 drain_right.t3 a_n2102_n1088# 0.020541f
C30 drain_right.n5 a_n2102_n1088# 0.079816f
C31 drain_right.n6 a_n2102_n1088# 0.55194f
C32 drain_right.n7 a_n2102_n1088# 0.944131f
C33 drain_right.t2 a_n2102_n1088# 0.020541f
C34 drain_right.t7 a_n2102_n1088# 0.020541f
C35 drain_right.n8 a_n2102_n1088# 0.080455f
C36 drain_right.t8 a_n2102_n1088# 0.020541f
C37 drain_right.t18 a_n2102_n1088# 0.020541f
C38 drain_right.n9 a_n2102_n1088# 0.079816f
C39 drain_right.n10 a_n2102_n1088# 0.55534f
C40 drain_right.t19 a_n2102_n1088# 0.020541f
C41 drain_right.t4 a_n2102_n1088# 0.020541f
C42 drain_right.n11 a_n2102_n1088# 0.079816f
C43 drain_right.n12 a_n2102_n1088# 0.272755f
C44 drain_right.t1 a_n2102_n1088# 0.020541f
C45 drain_right.t11 a_n2102_n1088# 0.020541f
C46 drain_right.n13 a_n2102_n1088# 0.079816f
C47 drain_right.n14 a_n2102_n1088# 0.272755f
C48 drain_right.t10 a_n2102_n1088# 0.020541f
C49 drain_right.t17 a_n2102_n1088# 0.020541f
C50 drain_right.n15 a_n2102_n1088# 0.079816f
C51 drain_right.n16 a_n2102_n1088# 0.489116f
C52 minus.n0 a_n2102_n1088# 0.028785f
C53 minus.t9 a_n2102_n1088# 0.032865f
C54 minus.t2 a_n2102_n1088# 0.02662f
C55 minus.t18 a_n2102_n1088# 0.02662f
C56 minus.n1 a_n2102_n1088# 0.010525f
C57 minus.n2 a_n2102_n1088# 0.028785f
C58 minus.t8 a_n2102_n1088# 0.02662f
C59 minus.n3 a_n2102_n1088# 0.027427f
C60 minus.t0 a_n2102_n1088# 0.02662f
C61 minus.t15 a_n2102_n1088# 0.02662f
C62 minus.t11 a_n2102_n1088# 0.02662f
C63 minus.n4 a_n2102_n1088# 0.027427f
C64 minus.n5 a_n2102_n1088# 0.028785f
C65 minus.t1 a_n2102_n1088# 0.02662f
C66 minus.t17 a_n2102_n1088# 0.02662f
C67 minus.n6 a_n2102_n1088# 0.027427f
C68 minus.t12 a_n2102_n1088# 0.032865f
C69 minus.n7 a_n2102_n1088# 0.035478f
C70 minus.n8 a_n2102_n1088# 0.065867f
C71 minus.n9 a_n2102_n1088# 0.011856f
C72 minus.n10 a_n2102_n1088# 0.027427f
C73 minus.n11 a_n2102_n1088# 0.01088f
C74 minus.n12 a_n2102_n1088# 0.010525f
C75 minus.n13 a_n2102_n1088# 0.028785f
C76 minus.n14 a_n2102_n1088# 0.028785f
C77 minus.n15 a_n2102_n1088# 0.011856f
C78 minus.n16 a_n2102_n1088# 0.027427f
C79 minus.n17 a_n2102_n1088# 0.011856f
C80 minus.n18 a_n2102_n1088# 0.027427f
C81 minus.n19 a_n2102_n1088# 0.011856f
C82 minus.n20 a_n2102_n1088# 0.028785f
C83 minus.n21 a_n2102_n1088# 0.028785f
C84 minus.n22 a_n2102_n1088# 0.028785f
C85 minus.n23 a_n2102_n1088# 0.01088f
C86 minus.n24 a_n2102_n1088# 0.027427f
C87 minus.n25 a_n2102_n1088# 0.011856f
C88 minus.n26 a_n2102_n1088# 0.027427f
C89 minus.n27 a_n2102_n1088# 0.035435f
C90 minus.n28 a_n2102_n1088# 0.696861f
C91 minus.n29 a_n2102_n1088# 0.028785f
C92 minus.t5 a_n2102_n1088# 0.02662f
C93 minus.t16 a_n2102_n1088# 0.02662f
C94 minus.n30 a_n2102_n1088# 0.010525f
C95 minus.n31 a_n2102_n1088# 0.028785f
C96 minus.t7 a_n2102_n1088# 0.02662f
C97 minus.t10 a_n2102_n1088# 0.02662f
C98 minus.t14 a_n2102_n1088# 0.02662f
C99 minus.n32 a_n2102_n1088# 0.027427f
C100 minus.n33 a_n2102_n1088# 0.028785f
C101 minus.t4 a_n2102_n1088# 0.02662f
C102 minus.t6 a_n2102_n1088# 0.02662f
C103 minus.n34 a_n2102_n1088# 0.027427f
C104 minus.t13 a_n2102_n1088# 0.032865f
C105 minus.n35 a_n2102_n1088# 0.035478f
C106 minus.n36 a_n2102_n1088# 0.065867f
C107 minus.n37 a_n2102_n1088# 0.011856f
C108 minus.n38 a_n2102_n1088# 0.027427f
C109 minus.n39 a_n2102_n1088# 0.01088f
C110 minus.n40 a_n2102_n1088# 0.010525f
C111 minus.n41 a_n2102_n1088# 0.028785f
C112 minus.n42 a_n2102_n1088# 0.028785f
C113 minus.n43 a_n2102_n1088# 0.011856f
C114 minus.n44 a_n2102_n1088# 0.027427f
C115 minus.n45 a_n2102_n1088# 0.011856f
C116 minus.n46 a_n2102_n1088# 0.027427f
C117 minus.t19 a_n2102_n1088# 0.02662f
C118 minus.n47 a_n2102_n1088# 0.027427f
C119 minus.n48 a_n2102_n1088# 0.011856f
C120 minus.n49 a_n2102_n1088# 0.028785f
C121 minus.n50 a_n2102_n1088# 0.028785f
C122 minus.n51 a_n2102_n1088# 0.028785f
C123 minus.n52 a_n2102_n1088# 0.01088f
C124 minus.n53 a_n2102_n1088# 0.027427f
C125 minus.n54 a_n2102_n1088# 0.011856f
C126 minus.n55 a_n2102_n1088# 0.027427f
C127 minus.t3 a_n2102_n1088# 0.032865f
C128 minus.n56 a_n2102_n1088# 0.035435f
C129 minus.n57 a_n2102_n1088# 0.189247f
C130 minus.n58 a_n2102_n1088# 0.860482f
C131 drain_left.t2 a_n2102_n1088# 0.02021f
C132 drain_left.t13 a_n2102_n1088# 0.02021f
C133 drain_left.n0 a_n2102_n1088# 0.079157f
C134 drain_left.t12 a_n2102_n1088# 0.02021f
C135 drain_left.t4 a_n2102_n1088# 0.02021f
C136 drain_left.n1 a_n2102_n1088# 0.078528f
C137 drain_left.n2 a_n2102_n1088# 0.543034f
C138 drain_left.t16 a_n2102_n1088# 0.02021f
C139 drain_left.t14 a_n2102_n1088# 0.02021f
C140 drain_left.n3 a_n2102_n1088# 0.078528f
C141 drain_left.t17 a_n2102_n1088# 0.02021f
C142 drain_left.t9 a_n2102_n1088# 0.02021f
C143 drain_left.n4 a_n2102_n1088# 0.079157f
C144 drain_left.t6 a_n2102_n1088# 0.02021f
C145 drain_left.t19 a_n2102_n1088# 0.02021f
C146 drain_left.n5 a_n2102_n1088# 0.078528f
C147 drain_left.n6 a_n2102_n1088# 0.543034f
C148 drain_left.n7 a_n2102_n1088# 0.978236f
C149 drain_left.t15 a_n2102_n1088# 0.02021f
C150 drain_left.t10 a_n2102_n1088# 0.02021f
C151 drain_left.n8 a_n2102_n1088# 0.079157f
C152 drain_left.t5 a_n2102_n1088# 0.02021f
C153 drain_left.t0 a_n2102_n1088# 0.02021f
C154 drain_left.n9 a_n2102_n1088# 0.078528f
C155 drain_left.n10 a_n2102_n1088# 0.546379f
C156 drain_left.t11 a_n2102_n1088# 0.02021f
C157 drain_left.t7 a_n2102_n1088# 0.02021f
C158 drain_left.n11 a_n2102_n1088# 0.078528f
C159 drain_left.n12 a_n2102_n1088# 0.268353f
C160 drain_left.t1 a_n2102_n1088# 0.02021f
C161 drain_left.t18 a_n2102_n1088# 0.02021f
C162 drain_left.n13 a_n2102_n1088# 0.078528f
C163 drain_left.n14 a_n2102_n1088# 0.268353f
C164 drain_left.t8 a_n2102_n1088# 0.02021f
C165 drain_left.t3 a_n2102_n1088# 0.02021f
C166 drain_left.n15 a_n2102_n1088# 0.078528f
C167 drain_left.n16 a_n2102_n1088# 0.481224f
C168 source.t28 a_n2102_n1088# 0.134785f
C169 source.n0 a_n2102_n1088# 0.578747f
C170 source.t14 a_n2102_n1088# 0.024216f
C171 source.t17 a_n2102_n1088# 0.024216f
C172 source.n1 a_n2102_n1088# 0.078538f
C173 source.n2 a_n2102_n1088# 0.295467f
C174 source.t19 a_n2102_n1088# 0.024216f
C175 source.t13 a_n2102_n1088# 0.024216f
C176 source.n3 a_n2102_n1088# 0.078538f
C177 source.n4 a_n2102_n1088# 0.295467f
C178 source.t26 a_n2102_n1088# 0.024216f
C179 source.t21 a_n2102_n1088# 0.024216f
C180 source.n5 a_n2102_n1088# 0.078538f
C181 source.n6 a_n2102_n1088# 0.295467f
C182 source.t23 a_n2102_n1088# 0.024216f
C183 source.t18 a_n2102_n1088# 0.024216f
C184 source.n7 a_n2102_n1088# 0.078538f
C185 source.n8 a_n2102_n1088# 0.295467f
C186 source.t32 a_n2102_n1088# 0.134785f
C187 source.n9 a_n2102_n1088# 0.298029f
C188 source.t33 a_n2102_n1088# 0.134785f
C189 source.n10 a_n2102_n1088# 0.298029f
C190 source.t3 a_n2102_n1088# 0.024216f
C191 source.t35 a_n2102_n1088# 0.024216f
C192 source.n11 a_n2102_n1088# 0.078538f
C193 source.n12 a_n2102_n1088# 0.295467f
C194 source.t38 a_n2102_n1088# 0.024216f
C195 source.t37 a_n2102_n1088# 0.024216f
C196 source.n13 a_n2102_n1088# 0.078538f
C197 source.n14 a_n2102_n1088# 0.295467f
C198 source.t0 a_n2102_n1088# 0.024216f
C199 source.t4 a_n2102_n1088# 0.024216f
C200 source.n15 a_n2102_n1088# 0.078538f
C201 source.n16 a_n2102_n1088# 0.295467f
C202 source.t8 a_n2102_n1088# 0.024216f
C203 source.t9 a_n2102_n1088# 0.024216f
C204 source.n17 a_n2102_n1088# 0.078538f
C205 source.n18 a_n2102_n1088# 0.295467f
C206 source.t34 a_n2102_n1088# 0.134785f
C207 source.n19 a_n2102_n1088# 0.824304f
C208 source.t15 a_n2102_n1088# 0.134785f
C209 source.n20 a_n2102_n1088# 0.824304f
C210 source.t24 a_n2102_n1088# 0.024216f
C211 source.t25 a_n2102_n1088# 0.024216f
C212 source.n21 a_n2102_n1088# 0.078538f
C213 source.n22 a_n2102_n1088# 0.295467f
C214 source.t27 a_n2102_n1088# 0.024216f
C215 source.t31 a_n2102_n1088# 0.024216f
C216 source.n23 a_n2102_n1088# 0.078538f
C217 source.n24 a_n2102_n1088# 0.295467f
C218 source.t20 a_n2102_n1088# 0.024216f
C219 source.t30 a_n2102_n1088# 0.024216f
C220 source.n25 a_n2102_n1088# 0.078538f
C221 source.n26 a_n2102_n1088# 0.295467f
C222 source.t16 a_n2102_n1088# 0.024216f
C223 source.t22 a_n2102_n1088# 0.024216f
C224 source.n27 a_n2102_n1088# 0.078538f
C225 source.n28 a_n2102_n1088# 0.295467f
C226 source.t29 a_n2102_n1088# 0.134785f
C227 source.n29 a_n2102_n1088# 0.298029f
C228 source.t12 a_n2102_n1088# 0.134785f
C229 source.n30 a_n2102_n1088# 0.298029f
C230 source.t2 a_n2102_n1088# 0.024216f
C231 source.t5 a_n2102_n1088# 0.024216f
C232 source.n31 a_n2102_n1088# 0.078538f
C233 source.n32 a_n2102_n1088# 0.295467f
C234 source.t11 a_n2102_n1088# 0.024216f
C235 source.t39 a_n2102_n1088# 0.024216f
C236 source.n33 a_n2102_n1088# 0.078538f
C237 source.n34 a_n2102_n1088# 0.295467f
C238 source.t1 a_n2102_n1088# 0.024216f
C239 source.t10 a_n2102_n1088# 0.024216f
C240 source.n35 a_n2102_n1088# 0.078538f
C241 source.n36 a_n2102_n1088# 0.295467f
C242 source.t36 a_n2102_n1088# 0.024216f
C243 source.t7 a_n2102_n1088# 0.024216f
C244 source.n37 a_n2102_n1088# 0.078538f
C245 source.n38 a_n2102_n1088# 0.295467f
C246 source.t6 a_n2102_n1088# 0.134785f
C247 source.n39 a_n2102_n1088# 0.471019f
C248 source.n40 a_n2102_n1088# 0.62064f
C249 plus.n0 a_n2102_n1088# 0.029245f
C250 plus.t11 a_n2102_n1088# 0.027046f
C251 plus.t1 a_n2102_n1088# 0.027046f
C252 plus.n1 a_n2102_n1088# 0.010693f
C253 plus.n2 a_n2102_n1088# 0.029245f
C254 plus.t12 a_n2102_n1088# 0.027046f
C255 plus.t8 a_n2102_n1088# 0.027046f
C256 plus.t19 a_n2102_n1088# 0.027046f
C257 plus.n3 a_n2102_n1088# 0.027865f
C258 plus.n4 a_n2102_n1088# 0.029245f
C259 plus.t14 a_n2102_n1088# 0.027046f
C260 plus.t9 a_n2102_n1088# 0.027046f
C261 plus.n5 a_n2102_n1088# 0.027865f
C262 plus.t4 a_n2102_n1088# 0.03339f
C263 plus.n6 a_n2102_n1088# 0.036045f
C264 plus.n7 a_n2102_n1088# 0.066919f
C265 plus.n8 a_n2102_n1088# 0.012045f
C266 plus.n9 a_n2102_n1088# 0.027865f
C267 plus.n10 a_n2102_n1088# 0.011054f
C268 plus.n11 a_n2102_n1088# 0.010693f
C269 plus.n12 a_n2102_n1088# 0.029245f
C270 plus.n13 a_n2102_n1088# 0.029245f
C271 plus.n14 a_n2102_n1088# 0.012045f
C272 plus.n15 a_n2102_n1088# 0.027865f
C273 plus.n16 a_n2102_n1088# 0.012045f
C274 plus.n17 a_n2102_n1088# 0.027865f
C275 plus.t18 a_n2102_n1088# 0.027046f
C276 plus.n18 a_n2102_n1088# 0.027865f
C277 plus.n19 a_n2102_n1088# 0.012045f
C278 plus.n20 a_n2102_n1088# 0.029245f
C279 plus.n21 a_n2102_n1088# 0.029245f
C280 plus.n22 a_n2102_n1088# 0.029245f
C281 plus.n23 a_n2102_n1088# 0.011054f
C282 plus.n24 a_n2102_n1088# 0.027865f
C283 plus.n25 a_n2102_n1088# 0.012045f
C284 plus.n26 a_n2102_n1088# 0.027865f
C285 plus.t16 a_n2102_n1088# 0.03339f
C286 plus.n27 a_n2102_n1088# 0.036001f
C287 plus.n28 a_n2102_n1088# 0.201637f
C288 plus.n29 a_n2102_n1088# 0.029245f
C289 plus.t17 a_n2102_n1088# 0.03339f
C290 plus.t6 a_n2102_n1088# 0.027046f
C291 plus.t7 a_n2102_n1088# 0.027046f
C292 plus.n30 a_n2102_n1088# 0.010693f
C293 plus.n31 a_n2102_n1088# 0.029245f
C294 plus.t15 a_n2102_n1088# 0.027046f
C295 plus.n32 a_n2102_n1088# 0.027865f
C296 plus.t3 a_n2102_n1088# 0.027046f
C297 plus.t5 a_n2102_n1088# 0.027046f
C298 plus.t13 a_n2102_n1088# 0.027046f
C299 plus.n33 a_n2102_n1088# 0.027865f
C300 plus.n34 a_n2102_n1088# 0.029245f
C301 plus.t0 a_n2102_n1088# 0.027046f
C302 plus.t2 a_n2102_n1088# 0.027046f
C303 plus.n35 a_n2102_n1088# 0.027865f
C304 plus.t10 a_n2102_n1088# 0.03339f
C305 plus.n36 a_n2102_n1088# 0.036045f
C306 plus.n37 a_n2102_n1088# 0.066919f
C307 plus.n38 a_n2102_n1088# 0.012045f
C308 plus.n39 a_n2102_n1088# 0.027865f
C309 plus.n40 a_n2102_n1088# 0.011054f
C310 plus.n41 a_n2102_n1088# 0.010693f
C311 plus.n42 a_n2102_n1088# 0.029245f
C312 plus.n43 a_n2102_n1088# 0.029245f
C313 plus.n44 a_n2102_n1088# 0.012045f
C314 plus.n45 a_n2102_n1088# 0.027865f
C315 plus.n46 a_n2102_n1088# 0.012045f
C316 plus.n47 a_n2102_n1088# 0.027865f
C317 plus.n48 a_n2102_n1088# 0.012045f
C318 plus.n49 a_n2102_n1088# 0.029245f
C319 plus.n50 a_n2102_n1088# 0.029245f
C320 plus.n51 a_n2102_n1088# 0.029245f
C321 plus.n52 a_n2102_n1088# 0.011054f
C322 plus.n53 a_n2102_n1088# 0.027865f
C323 plus.n54 a_n2102_n1088# 0.012045f
C324 plus.n55 a_n2102_n1088# 0.027865f
C325 plus.n56 a_n2102_n1088# 0.036001f
C326 plus.n57 a_n2102_n1088# 0.684917f
.ends

