* NGSPICE file created from diffpair331.ext - technology: sky130A

.subckt diffpair331 minus drain_right drain_left source plus
X0 drain_right.t3 minus.t0 source.t4 a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X1 a_n1034_n2692# a_n1034_n2692# a_n1034_n2692# a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.2
X2 a_n1034_n2692# a_n1034_n2692# a_n1034_n2692# a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X3 drain_left.t3 plus.t0 source.t1 a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X4 a_n1034_n2692# a_n1034_n2692# a_n1034_n2692# a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X5 source.t3 plus.t1 drain_left.t2 a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X6 source.t7 minus.t1 drain_right.t2 a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X7 drain_right.t1 minus.t2 source.t5 a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X8 drain_left.t1 plus.t2 source.t2 a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.2
X9 a_n1034_n2692# a_n1034_n2692# a_n1034_n2692# a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.2
X10 source.t6 minus.t3 drain_right.t0 a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
X11 source.t0 plus.t3 drain_left.t0 a_n1034_n2692# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.2
R0 minus.n0 minus.t3 1279.86
R1 minus.n0 minus.t0 1279.86
R2 minus.n1 minus.t2 1279.86
R3 minus.n1 minus.t1 1279.86
R4 minus.n2 minus.n0 192.012
R5 minus.n2 minus.n1 167.732
R6 minus minus.n2 0.188
R7 source.n1 source.t0 51.0588
R8 source.n2 source.t4 51.0588
R9 source.n3 source.t6 51.0588
R10 source.n7 source.t5 51.0586
R11 source.n6 source.t7 51.0586
R12 source.n5 source.t1 51.0586
R13 source.n4 source.t3 51.0586
R14 source.n0 source.t2 51.0586
R15 source.n4 source.n3 19.487
R16 source.n8 source.n0 13.9957
R17 source.n8 source.n7 5.49188
R18 source.n2 source.n1 0.470328
R19 source.n6 source.n5 0.470328
R20 source.n3 source.n2 0.457397
R21 source.n1 source.n0 0.457397
R22 source.n5 source.n4 0.457397
R23 source.n7 source.n6 0.457397
R24 source source.n8 0.188
R25 drain_right drain_right.n0 91.0069
R26 drain_right drain_right.n1 71.647
R27 drain_right.n0 drain_right.t2 2.2005
R28 drain_right.n0 drain_right.t1 2.2005
R29 drain_right.n1 drain_right.t0 2.2005
R30 drain_right.n1 drain_right.t3 2.2005
R31 plus.n0 plus.t3 1279.86
R32 plus.n0 plus.t2 1279.86
R33 plus.n1 plus.t0 1279.86
R34 plus.n1 plus.t1 1279.86
R35 plus plus.n1 187.03
R36 plus plus.n0 172.239
R37 drain_left drain_left.n0 91.5601
R38 drain_left drain_left.n1 71.647
R39 drain_left.n0 drain_left.t2 2.2005
R40 drain_left.n0 drain_left.t3 2.2005
R41 drain_left.n1 drain_left.t0 2.2005
R42 drain_left.n1 drain_left.t1 2.2005
C0 source drain_right 8.6641f
C1 minus drain_right 1.35948f
C2 source minus 0.926542f
C3 plus drain_left 1.45419f
C4 plus drain_right 0.248706f
C5 plus source 0.940581f
C6 plus minus 3.88444f
C7 drain_left drain_right 0.457115f
C8 drain_left source 8.666151f
C9 drain_left minus 0.171239f
C10 drain_right a_n1034_n2692# 5.80617f
C11 drain_left a_n1034_n2692# 5.95363f
C12 source a_n1034_n2692# 6.440058f
C13 minus a_n1034_n2692# 3.739792f
C14 plus a_n1034_n2692# 6.10921f
C15 drain_left.t2 a_n1034_n2692# 0.214129f
C16 drain_left.t3 a_n1034_n2692# 0.214129f
C17 drain_left.n0 a_n1034_n2692# 2.2042f
C18 drain_left.t0 a_n1034_n2692# 0.214129f
C19 drain_left.t1 a_n1034_n2692# 0.214129f
C20 drain_left.n1 a_n1034_n2692# 1.92308f
C21 plus.t3 a_n1034_n2692# 0.210782f
C22 plus.t2 a_n1034_n2692# 0.210782f
C23 plus.n0 a_n1034_n2692# 0.214603f
C24 plus.t1 a_n1034_n2692# 0.210782f
C25 plus.t0 a_n1034_n2692# 0.210782f
C26 plus.n1 a_n1034_n2692# 0.321957f
C27 drain_right.t2 a_n1034_n2692# 0.217067f
C28 drain_right.t1 a_n1034_n2692# 0.217067f
C29 drain_right.n0 a_n1034_n2692# 2.21144f
C30 drain_right.t0 a_n1034_n2692# 0.217067f
C31 drain_right.t3 a_n1034_n2692# 0.217067f
C32 drain_right.n1 a_n1034_n2692# 1.94947f
C33 source.t2 a_n1034_n2692# 1.46411f
C34 source.n0 a_n1034_n2692# 0.833963f
C35 source.t0 a_n1034_n2692# 1.46411f
C36 source.n1 a_n1034_n2692# 0.297321f
C37 source.t4 a_n1034_n2692# 1.46411f
C38 source.n2 a_n1034_n2692# 0.297321f
C39 source.t6 a_n1034_n2692# 1.46411f
C40 source.n3 a_n1034_n2692# 1.1129f
C41 source.t3 a_n1034_n2692# 1.46411f
C42 source.n4 a_n1034_n2692# 1.1129f
C43 source.t1 a_n1034_n2692# 1.46411f
C44 source.n5 a_n1034_n2692# 0.297325f
C45 source.t7 a_n1034_n2692# 1.46411f
C46 source.n6 a_n1034_n2692# 0.297325f
C47 source.t5 a_n1034_n2692# 1.46411f
C48 source.n7 a_n1034_n2692# 0.402005f
C49 source.n8 a_n1034_n2692# 1.00357f
C50 minus.t3 a_n1034_n2692# 0.206416f
C51 minus.t0 a_n1034_n2692# 0.206416f
C52 minus.n0 a_n1034_n2692# 0.358734f
C53 minus.t1 a_n1034_n2692# 0.206416f
C54 minus.t2 a_n1034_n2692# 0.206416f
C55 minus.n1 a_n1034_n2692# 0.19528f
C56 minus.n2 a_n1034_n2692# 2.49409f
.ends

