* NGSPICE file created from diffpair676.ext - technology: sky130A

.subckt diffpair676 minus drain_right drain_left source plus
X0 source.t27 minus.t0 drain_right.t1 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X1 drain_right.t0 minus.t1 source.t26 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X2 a_n1724_n5888# a_n1724_n5888# a_n1724_n5888# a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.3
X3 drain_right.t3 minus.t2 source.t25 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X4 drain_right.t2 minus.t3 source.t24 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X5 drain_left.t13 plus.t0 source.t7 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X6 drain_right.t5 minus.t4 source.t23 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X7 drain_left.t12 plus.t1 source.t2 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X8 drain_left.t11 plus.t2 source.t0 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X9 a_n1724_n5888# a_n1724_n5888# a_n1724_n5888# a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X10 drain_left.t10 plus.t3 source.t1 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X11 source.t4 plus.t4 drain_left.t9 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X12 drain_right.t4 minus.t5 source.t22 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X13 drain_right.t11 minus.t6 source.t21 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X14 source.t20 minus.t7 drain_right.t10 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X15 source.t10 plus.t5 drain_left.t8 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X16 drain_right.t9 minus.t8 source.t19 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X17 source.t6 plus.t6 drain_left.t7 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X18 source.t12 plus.t7 drain_left.t6 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X19 drain_left.t5 plus.t8 source.t13 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X20 source.t5 plus.t9 drain_left.t4 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X21 source.t18 minus.t9 drain_right.t8 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X22 source.t17 minus.t10 drain_right.t7 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X23 a_n1724_n5888# a_n1724_n5888# a_n1724_n5888# a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X24 drain_right.t6 minus.t11 source.t16 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X25 a_n1724_n5888# a_n1724_n5888# a_n1724_n5888# a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X26 source.t15 minus.t12 drain_right.t13 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X27 source.t14 minus.t13 drain_right.t12 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X28 drain_left.t3 plus.t10 source.t8 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X29 source.t11 plus.t11 drain_left.t2 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X30 drain_left.t1 plus.t12 source.t3 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X31 drain_left.t0 plus.t13 source.t9 a_n1724_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
R0 minus.n15 minus.t4 2169.73
R1 minus.n3 minus.t8 2169.73
R2 minus.n32 minus.t5 2169.73
R3 minus.n20 minus.t3 2169.73
R4 minus.n1 minus.t7 2112.77
R5 minus.n14 minus.t0 2112.77
R6 minus.n12 minus.t11 2112.77
R7 minus.n6 minus.t1 2112.77
R8 minus.n4 minus.t12 2112.77
R9 minus.n18 minus.t9 2112.77
R10 minus.n31 minus.t13 2112.77
R11 minus.n29 minus.t6 2112.77
R12 minus.n23 minus.t2 2112.77
R13 minus.n21 minus.t10 2112.77
R14 minus.n3 minus.n2 161.489
R15 minus.n20 minus.n19 161.489
R16 minus.n16 minus.n15 161.3
R17 minus.n13 minus.n0 161.3
R18 minus.n11 minus.n10 161.3
R19 minus.n9 minus.n1 161.3
R20 minus.n8 minus.n7 161.3
R21 minus.n5 minus.n2 161.3
R22 minus.n33 minus.n32 161.3
R23 minus.n30 minus.n17 161.3
R24 minus.n28 minus.n27 161.3
R25 minus.n26 minus.n18 161.3
R26 minus.n25 minus.n24 161.3
R27 minus.n22 minus.n19 161.3
R28 minus.n11 minus.n1 73.0308
R29 minus.n7 minus.n1 73.0308
R30 minus.n24 minus.n18 73.0308
R31 minus.n28 minus.n18 73.0308
R32 minus.n13 minus.n12 54.0429
R33 minus.n6 minus.n5 54.0429
R34 minus.n23 minus.n22 54.0429
R35 minus.n30 minus.n29 54.0429
R36 minus.n34 minus.n16 45.5365
R37 minus.n14 minus.n13 37.9763
R38 minus.n5 minus.n4 37.9763
R39 minus.n22 minus.n21 37.9763
R40 minus.n31 minus.n30 37.9763
R41 minus.n15 minus.n14 35.055
R42 minus.n4 minus.n3 35.055
R43 minus.n21 minus.n20 35.055
R44 minus.n32 minus.n31 35.055
R45 minus.n12 minus.n11 18.9884
R46 minus.n7 minus.n6 18.9884
R47 minus.n24 minus.n23 18.9884
R48 minus.n29 minus.n28 18.9884
R49 minus.n34 minus.n33 6.53648
R50 minus.n16 minus.n0 0.189894
R51 minus.n10 minus.n0 0.189894
R52 minus.n10 minus.n9 0.189894
R53 minus.n9 minus.n8 0.189894
R54 minus.n8 minus.n2 0.189894
R55 minus.n25 minus.n19 0.189894
R56 minus.n26 minus.n25 0.189894
R57 minus.n27 minus.n26 0.189894
R58 minus.n27 minus.n17 0.189894
R59 minus.n33 minus.n17 0.189894
R60 minus minus.n34 0.188
R61 drain_right.n134 drain_right.n0 289.615
R62 drain_right.n284 drain_right.n150 289.615
R63 drain_right.n44 drain_right.n43 185
R64 drain_right.n49 drain_right.n48 185
R65 drain_right.n51 drain_right.n50 185
R66 drain_right.n40 drain_right.n39 185
R67 drain_right.n57 drain_right.n56 185
R68 drain_right.n59 drain_right.n58 185
R69 drain_right.n36 drain_right.n35 185
R70 drain_right.n66 drain_right.n65 185
R71 drain_right.n67 drain_right.n34 185
R72 drain_right.n69 drain_right.n68 185
R73 drain_right.n32 drain_right.n31 185
R74 drain_right.n75 drain_right.n74 185
R75 drain_right.n77 drain_right.n76 185
R76 drain_right.n28 drain_right.n27 185
R77 drain_right.n83 drain_right.n82 185
R78 drain_right.n85 drain_right.n84 185
R79 drain_right.n24 drain_right.n23 185
R80 drain_right.n91 drain_right.n90 185
R81 drain_right.n93 drain_right.n92 185
R82 drain_right.n20 drain_right.n19 185
R83 drain_right.n99 drain_right.n98 185
R84 drain_right.n101 drain_right.n100 185
R85 drain_right.n16 drain_right.n15 185
R86 drain_right.n107 drain_right.n106 185
R87 drain_right.n110 drain_right.n109 185
R88 drain_right.n108 drain_right.n12 185
R89 drain_right.n115 drain_right.n11 185
R90 drain_right.n117 drain_right.n116 185
R91 drain_right.n119 drain_right.n118 185
R92 drain_right.n8 drain_right.n7 185
R93 drain_right.n125 drain_right.n124 185
R94 drain_right.n127 drain_right.n126 185
R95 drain_right.n4 drain_right.n3 185
R96 drain_right.n133 drain_right.n132 185
R97 drain_right.n135 drain_right.n134 185
R98 drain_right.n285 drain_right.n284 185
R99 drain_right.n283 drain_right.n282 185
R100 drain_right.n154 drain_right.n153 185
R101 drain_right.n277 drain_right.n276 185
R102 drain_right.n275 drain_right.n274 185
R103 drain_right.n158 drain_right.n157 185
R104 drain_right.n269 drain_right.n268 185
R105 drain_right.n267 drain_right.n266 185
R106 drain_right.n265 drain_right.n161 185
R107 drain_right.n165 drain_right.n162 185
R108 drain_right.n260 drain_right.n259 185
R109 drain_right.n258 drain_right.n257 185
R110 drain_right.n167 drain_right.n166 185
R111 drain_right.n252 drain_right.n251 185
R112 drain_right.n250 drain_right.n249 185
R113 drain_right.n171 drain_right.n170 185
R114 drain_right.n244 drain_right.n243 185
R115 drain_right.n242 drain_right.n241 185
R116 drain_right.n175 drain_right.n174 185
R117 drain_right.n236 drain_right.n235 185
R118 drain_right.n234 drain_right.n233 185
R119 drain_right.n179 drain_right.n178 185
R120 drain_right.n228 drain_right.n227 185
R121 drain_right.n226 drain_right.n225 185
R122 drain_right.n183 drain_right.n182 185
R123 drain_right.n220 drain_right.n219 185
R124 drain_right.n218 drain_right.n185 185
R125 drain_right.n217 drain_right.n216 185
R126 drain_right.n188 drain_right.n186 185
R127 drain_right.n211 drain_right.n210 185
R128 drain_right.n209 drain_right.n208 185
R129 drain_right.n192 drain_right.n191 185
R130 drain_right.n203 drain_right.n202 185
R131 drain_right.n201 drain_right.n200 185
R132 drain_right.n196 drain_right.n195 185
R133 drain_right.n45 drain_right.t2 149.524
R134 drain_right.n197 drain_right.t5 149.524
R135 drain_right.n49 drain_right.n43 104.615
R136 drain_right.n50 drain_right.n49 104.615
R137 drain_right.n50 drain_right.n39 104.615
R138 drain_right.n57 drain_right.n39 104.615
R139 drain_right.n58 drain_right.n57 104.615
R140 drain_right.n58 drain_right.n35 104.615
R141 drain_right.n66 drain_right.n35 104.615
R142 drain_right.n67 drain_right.n66 104.615
R143 drain_right.n68 drain_right.n67 104.615
R144 drain_right.n68 drain_right.n31 104.615
R145 drain_right.n75 drain_right.n31 104.615
R146 drain_right.n76 drain_right.n75 104.615
R147 drain_right.n76 drain_right.n27 104.615
R148 drain_right.n83 drain_right.n27 104.615
R149 drain_right.n84 drain_right.n83 104.615
R150 drain_right.n84 drain_right.n23 104.615
R151 drain_right.n91 drain_right.n23 104.615
R152 drain_right.n92 drain_right.n91 104.615
R153 drain_right.n92 drain_right.n19 104.615
R154 drain_right.n99 drain_right.n19 104.615
R155 drain_right.n100 drain_right.n99 104.615
R156 drain_right.n100 drain_right.n15 104.615
R157 drain_right.n107 drain_right.n15 104.615
R158 drain_right.n109 drain_right.n107 104.615
R159 drain_right.n109 drain_right.n108 104.615
R160 drain_right.n108 drain_right.n11 104.615
R161 drain_right.n117 drain_right.n11 104.615
R162 drain_right.n118 drain_right.n117 104.615
R163 drain_right.n118 drain_right.n7 104.615
R164 drain_right.n125 drain_right.n7 104.615
R165 drain_right.n126 drain_right.n125 104.615
R166 drain_right.n126 drain_right.n3 104.615
R167 drain_right.n133 drain_right.n3 104.615
R168 drain_right.n134 drain_right.n133 104.615
R169 drain_right.n284 drain_right.n283 104.615
R170 drain_right.n283 drain_right.n153 104.615
R171 drain_right.n276 drain_right.n153 104.615
R172 drain_right.n276 drain_right.n275 104.615
R173 drain_right.n275 drain_right.n157 104.615
R174 drain_right.n268 drain_right.n157 104.615
R175 drain_right.n268 drain_right.n267 104.615
R176 drain_right.n267 drain_right.n161 104.615
R177 drain_right.n165 drain_right.n161 104.615
R178 drain_right.n259 drain_right.n165 104.615
R179 drain_right.n259 drain_right.n258 104.615
R180 drain_right.n258 drain_right.n166 104.615
R181 drain_right.n251 drain_right.n166 104.615
R182 drain_right.n251 drain_right.n250 104.615
R183 drain_right.n250 drain_right.n170 104.615
R184 drain_right.n243 drain_right.n170 104.615
R185 drain_right.n243 drain_right.n242 104.615
R186 drain_right.n242 drain_right.n174 104.615
R187 drain_right.n235 drain_right.n174 104.615
R188 drain_right.n235 drain_right.n234 104.615
R189 drain_right.n234 drain_right.n178 104.615
R190 drain_right.n227 drain_right.n178 104.615
R191 drain_right.n227 drain_right.n226 104.615
R192 drain_right.n226 drain_right.n182 104.615
R193 drain_right.n219 drain_right.n182 104.615
R194 drain_right.n219 drain_right.n218 104.615
R195 drain_right.n218 drain_right.n217 104.615
R196 drain_right.n217 drain_right.n186 104.615
R197 drain_right.n210 drain_right.n186 104.615
R198 drain_right.n210 drain_right.n209 104.615
R199 drain_right.n209 drain_right.n191 104.615
R200 drain_right.n202 drain_right.n191 104.615
R201 drain_right.n202 drain_right.n201 104.615
R202 drain_right.n201 drain_right.n195 104.615
R203 drain_right.n143 drain_right.n141 59.2585
R204 drain_right.n147 drain_right.n145 59.2584
R205 drain_right.n143 drain_right.n142 58.7154
R206 drain_right.n140 drain_right.n139 58.7154
R207 drain_right.n147 drain_right.n146 58.7154
R208 drain_right.n149 drain_right.n148 58.7154
R209 drain_right.t2 drain_right.n43 52.3082
R210 drain_right.t5 drain_right.n195 52.3082
R211 drain_right.n140 drain_right.n138 47.8557
R212 drain_right.n289 drain_right.n288 47.3126
R213 drain_right drain_right.n144 39.7852
R214 drain_right.n69 drain_right.n34 13.1884
R215 drain_right.n116 drain_right.n115 13.1884
R216 drain_right.n266 drain_right.n265 13.1884
R217 drain_right.n220 drain_right.n185 13.1884
R218 drain_right.n65 drain_right.n64 12.8005
R219 drain_right.n70 drain_right.n32 12.8005
R220 drain_right.n114 drain_right.n12 12.8005
R221 drain_right.n119 drain_right.n10 12.8005
R222 drain_right.n269 drain_right.n160 12.8005
R223 drain_right.n264 drain_right.n162 12.8005
R224 drain_right.n221 drain_right.n183 12.8005
R225 drain_right.n216 drain_right.n187 12.8005
R226 drain_right.n63 drain_right.n36 12.0247
R227 drain_right.n74 drain_right.n73 12.0247
R228 drain_right.n111 drain_right.n110 12.0247
R229 drain_right.n120 drain_right.n8 12.0247
R230 drain_right.n270 drain_right.n158 12.0247
R231 drain_right.n261 drain_right.n260 12.0247
R232 drain_right.n225 drain_right.n224 12.0247
R233 drain_right.n215 drain_right.n188 12.0247
R234 drain_right.n60 drain_right.n59 11.249
R235 drain_right.n77 drain_right.n30 11.249
R236 drain_right.n106 drain_right.n14 11.249
R237 drain_right.n124 drain_right.n123 11.249
R238 drain_right.n274 drain_right.n273 11.249
R239 drain_right.n257 drain_right.n164 11.249
R240 drain_right.n228 drain_right.n181 11.249
R241 drain_right.n212 drain_right.n211 11.249
R242 drain_right.n56 drain_right.n38 10.4732
R243 drain_right.n78 drain_right.n28 10.4732
R244 drain_right.n105 drain_right.n16 10.4732
R245 drain_right.n127 drain_right.n6 10.4732
R246 drain_right.n277 drain_right.n156 10.4732
R247 drain_right.n256 drain_right.n167 10.4732
R248 drain_right.n229 drain_right.n179 10.4732
R249 drain_right.n208 drain_right.n190 10.4732
R250 drain_right.n45 drain_right.n44 10.2747
R251 drain_right.n197 drain_right.n196 10.2747
R252 drain_right.n55 drain_right.n40 9.69747
R253 drain_right.n82 drain_right.n81 9.69747
R254 drain_right.n102 drain_right.n101 9.69747
R255 drain_right.n128 drain_right.n4 9.69747
R256 drain_right.n278 drain_right.n154 9.69747
R257 drain_right.n253 drain_right.n252 9.69747
R258 drain_right.n233 drain_right.n232 9.69747
R259 drain_right.n207 drain_right.n192 9.69747
R260 drain_right.n138 drain_right.n137 9.45567
R261 drain_right.n288 drain_right.n287 9.45567
R262 drain_right.n2 drain_right.n1 9.3005
R263 drain_right.n131 drain_right.n130 9.3005
R264 drain_right.n129 drain_right.n128 9.3005
R265 drain_right.n6 drain_right.n5 9.3005
R266 drain_right.n123 drain_right.n122 9.3005
R267 drain_right.n121 drain_right.n120 9.3005
R268 drain_right.n10 drain_right.n9 9.3005
R269 drain_right.n89 drain_right.n88 9.3005
R270 drain_right.n87 drain_right.n86 9.3005
R271 drain_right.n26 drain_right.n25 9.3005
R272 drain_right.n81 drain_right.n80 9.3005
R273 drain_right.n79 drain_right.n78 9.3005
R274 drain_right.n30 drain_right.n29 9.3005
R275 drain_right.n73 drain_right.n72 9.3005
R276 drain_right.n71 drain_right.n70 9.3005
R277 drain_right.n47 drain_right.n46 9.3005
R278 drain_right.n42 drain_right.n41 9.3005
R279 drain_right.n53 drain_right.n52 9.3005
R280 drain_right.n55 drain_right.n54 9.3005
R281 drain_right.n38 drain_right.n37 9.3005
R282 drain_right.n61 drain_right.n60 9.3005
R283 drain_right.n63 drain_right.n62 9.3005
R284 drain_right.n64 drain_right.n33 9.3005
R285 drain_right.n22 drain_right.n21 9.3005
R286 drain_right.n95 drain_right.n94 9.3005
R287 drain_right.n97 drain_right.n96 9.3005
R288 drain_right.n18 drain_right.n17 9.3005
R289 drain_right.n103 drain_right.n102 9.3005
R290 drain_right.n105 drain_right.n104 9.3005
R291 drain_right.n14 drain_right.n13 9.3005
R292 drain_right.n112 drain_right.n111 9.3005
R293 drain_right.n114 drain_right.n113 9.3005
R294 drain_right.n137 drain_right.n136 9.3005
R295 drain_right.n199 drain_right.n198 9.3005
R296 drain_right.n194 drain_right.n193 9.3005
R297 drain_right.n205 drain_right.n204 9.3005
R298 drain_right.n207 drain_right.n206 9.3005
R299 drain_right.n190 drain_right.n189 9.3005
R300 drain_right.n213 drain_right.n212 9.3005
R301 drain_right.n215 drain_right.n214 9.3005
R302 drain_right.n187 drain_right.n184 9.3005
R303 drain_right.n246 drain_right.n245 9.3005
R304 drain_right.n248 drain_right.n247 9.3005
R305 drain_right.n169 drain_right.n168 9.3005
R306 drain_right.n254 drain_right.n253 9.3005
R307 drain_right.n256 drain_right.n255 9.3005
R308 drain_right.n164 drain_right.n163 9.3005
R309 drain_right.n262 drain_right.n261 9.3005
R310 drain_right.n264 drain_right.n263 9.3005
R311 drain_right.n287 drain_right.n286 9.3005
R312 drain_right.n152 drain_right.n151 9.3005
R313 drain_right.n281 drain_right.n280 9.3005
R314 drain_right.n279 drain_right.n278 9.3005
R315 drain_right.n156 drain_right.n155 9.3005
R316 drain_right.n273 drain_right.n272 9.3005
R317 drain_right.n271 drain_right.n270 9.3005
R318 drain_right.n160 drain_right.n159 9.3005
R319 drain_right.n173 drain_right.n172 9.3005
R320 drain_right.n240 drain_right.n239 9.3005
R321 drain_right.n238 drain_right.n237 9.3005
R322 drain_right.n177 drain_right.n176 9.3005
R323 drain_right.n232 drain_right.n231 9.3005
R324 drain_right.n230 drain_right.n229 9.3005
R325 drain_right.n181 drain_right.n180 9.3005
R326 drain_right.n224 drain_right.n223 9.3005
R327 drain_right.n222 drain_right.n221 9.3005
R328 drain_right.n52 drain_right.n51 8.92171
R329 drain_right.n85 drain_right.n26 8.92171
R330 drain_right.n98 drain_right.n18 8.92171
R331 drain_right.n132 drain_right.n131 8.92171
R332 drain_right.n282 drain_right.n281 8.92171
R333 drain_right.n249 drain_right.n169 8.92171
R334 drain_right.n236 drain_right.n177 8.92171
R335 drain_right.n204 drain_right.n203 8.92171
R336 drain_right.n48 drain_right.n42 8.14595
R337 drain_right.n86 drain_right.n24 8.14595
R338 drain_right.n97 drain_right.n20 8.14595
R339 drain_right.n135 drain_right.n2 8.14595
R340 drain_right.n285 drain_right.n152 8.14595
R341 drain_right.n248 drain_right.n171 8.14595
R342 drain_right.n237 drain_right.n175 8.14595
R343 drain_right.n200 drain_right.n194 8.14595
R344 drain_right.n47 drain_right.n44 7.3702
R345 drain_right.n90 drain_right.n89 7.3702
R346 drain_right.n94 drain_right.n93 7.3702
R347 drain_right.n136 drain_right.n0 7.3702
R348 drain_right.n286 drain_right.n150 7.3702
R349 drain_right.n245 drain_right.n244 7.3702
R350 drain_right.n241 drain_right.n240 7.3702
R351 drain_right.n199 drain_right.n196 7.3702
R352 drain_right.n90 drain_right.n22 6.59444
R353 drain_right.n93 drain_right.n22 6.59444
R354 drain_right.n138 drain_right.n0 6.59444
R355 drain_right.n288 drain_right.n150 6.59444
R356 drain_right.n244 drain_right.n173 6.59444
R357 drain_right.n241 drain_right.n173 6.59444
R358 drain_right drain_right.n289 5.92477
R359 drain_right.n48 drain_right.n47 5.81868
R360 drain_right.n89 drain_right.n24 5.81868
R361 drain_right.n94 drain_right.n20 5.81868
R362 drain_right.n136 drain_right.n135 5.81868
R363 drain_right.n286 drain_right.n285 5.81868
R364 drain_right.n245 drain_right.n171 5.81868
R365 drain_right.n240 drain_right.n175 5.81868
R366 drain_right.n200 drain_right.n199 5.81868
R367 drain_right.n51 drain_right.n42 5.04292
R368 drain_right.n86 drain_right.n85 5.04292
R369 drain_right.n98 drain_right.n97 5.04292
R370 drain_right.n132 drain_right.n2 5.04292
R371 drain_right.n282 drain_right.n152 5.04292
R372 drain_right.n249 drain_right.n248 5.04292
R373 drain_right.n237 drain_right.n236 5.04292
R374 drain_right.n203 drain_right.n194 5.04292
R375 drain_right.n52 drain_right.n40 4.26717
R376 drain_right.n82 drain_right.n26 4.26717
R377 drain_right.n101 drain_right.n18 4.26717
R378 drain_right.n131 drain_right.n4 4.26717
R379 drain_right.n281 drain_right.n154 4.26717
R380 drain_right.n252 drain_right.n169 4.26717
R381 drain_right.n233 drain_right.n177 4.26717
R382 drain_right.n204 drain_right.n192 4.26717
R383 drain_right.n56 drain_right.n55 3.49141
R384 drain_right.n81 drain_right.n28 3.49141
R385 drain_right.n102 drain_right.n16 3.49141
R386 drain_right.n128 drain_right.n127 3.49141
R387 drain_right.n278 drain_right.n277 3.49141
R388 drain_right.n253 drain_right.n167 3.49141
R389 drain_right.n232 drain_right.n179 3.49141
R390 drain_right.n208 drain_right.n207 3.49141
R391 drain_right.n198 drain_right.n197 2.84303
R392 drain_right.n46 drain_right.n45 2.84303
R393 drain_right.n59 drain_right.n38 2.71565
R394 drain_right.n78 drain_right.n77 2.71565
R395 drain_right.n106 drain_right.n105 2.71565
R396 drain_right.n124 drain_right.n6 2.71565
R397 drain_right.n274 drain_right.n156 2.71565
R398 drain_right.n257 drain_right.n256 2.71565
R399 drain_right.n229 drain_right.n228 2.71565
R400 drain_right.n211 drain_right.n190 2.71565
R401 drain_right.n60 drain_right.n36 1.93989
R402 drain_right.n74 drain_right.n30 1.93989
R403 drain_right.n110 drain_right.n14 1.93989
R404 drain_right.n123 drain_right.n8 1.93989
R405 drain_right.n273 drain_right.n158 1.93989
R406 drain_right.n260 drain_right.n164 1.93989
R407 drain_right.n225 drain_right.n181 1.93989
R408 drain_right.n212 drain_right.n188 1.93989
R409 drain_right.n65 drain_right.n63 1.16414
R410 drain_right.n73 drain_right.n32 1.16414
R411 drain_right.n111 drain_right.n12 1.16414
R412 drain_right.n120 drain_right.n119 1.16414
R413 drain_right.n270 drain_right.n269 1.16414
R414 drain_right.n261 drain_right.n162 1.16414
R415 drain_right.n224 drain_right.n183 1.16414
R416 drain_right.n216 drain_right.n215 1.16414
R417 drain_right.n141 drain_right.t12 0.7925
R418 drain_right.n141 drain_right.t4 0.7925
R419 drain_right.n142 drain_right.t8 0.7925
R420 drain_right.n142 drain_right.t11 0.7925
R421 drain_right.n139 drain_right.t7 0.7925
R422 drain_right.n139 drain_right.t3 0.7925
R423 drain_right.n145 drain_right.t13 0.7925
R424 drain_right.n145 drain_right.t9 0.7925
R425 drain_right.n146 drain_right.t10 0.7925
R426 drain_right.n146 drain_right.t0 0.7925
R427 drain_right.n148 drain_right.t1 0.7925
R428 drain_right.n148 drain_right.t6 0.7925
R429 drain_right.n289 drain_right.n149 0.543603
R430 drain_right.n149 drain_right.n147 0.543603
R431 drain_right.n64 drain_right.n34 0.388379
R432 drain_right.n70 drain_right.n69 0.388379
R433 drain_right.n115 drain_right.n114 0.388379
R434 drain_right.n116 drain_right.n10 0.388379
R435 drain_right.n266 drain_right.n160 0.388379
R436 drain_right.n265 drain_right.n264 0.388379
R437 drain_right.n221 drain_right.n220 0.388379
R438 drain_right.n187 drain_right.n185 0.388379
R439 drain_right.n144 drain_right.n140 0.352482
R440 drain_right.n46 drain_right.n41 0.155672
R441 drain_right.n53 drain_right.n41 0.155672
R442 drain_right.n54 drain_right.n53 0.155672
R443 drain_right.n54 drain_right.n37 0.155672
R444 drain_right.n61 drain_right.n37 0.155672
R445 drain_right.n62 drain_right.n61 0.155672
R446 drain_right.n62 drain_right.n33 0.155672
R447 drain_right.n71 drain_right.n33 0.155672
R448 drain_right.n72 drain_right.n71 0.155672
R449 drain_right.n72 drain_right.n29 0.155672
R450 drain_right.n79 drain_right.n29 0.155672
R451 drain_right.n80 drain_right.n79 0.155672
R452 drain_right.n80 drain_right.n25 0.155672
R453 drain_right.n87 drain_right.n25 0.155672
R454 drain_right.n88 drain_right.n87 0.155672
R455 drain_right.n88 drain_right.n21 0.155672
R456 drain_right.n95 drain_right.n21 0.155672
R457 drain_right.n96 drain_right.n95 0.155672
R458 drain_right.n96 drain_right.n17 0.155672
R459 drain_right.n103 drain_right.n17 0.155672
R460 drain_right.n104 drain_right.n103 0.155672
R461 drain_right.n104 drain_right.n13 0.155672
R462 drain_right.n112 drain_right.n13 0.155672
R463 drain_right.n113 drain_right.n112 0.155672
R464 drain_right.n113 drain_right.n9 0.155672
R465 drain_right.n121 drain_right.n9 0.155672
R466 drain_right.n122 drain_right.n121 0.155672
R467 drain_right.n122 drain_right.n5 0.155672
R468 drain_right.n129 drain_right.n5 0.155672
R469 drain_right.n130 drain_right.n129 0.155672
R470 drain_right.n130 drain_right.n1 0.155672
R471 drain_right.n137 drain_right.n1 0.155672
R472 drain_right.n287 drain_right.n151 0.155672
R473 drain_right.n280 drain_right.n151 0.155672
R474 drain_right.n280 drain_right.n279 0.155672
R475 drain_right.n279 drain_right.n155 0.155672
R476 drain_right.n272 drain_right.n155 0.155672
R477 drain_right.n272 drain_right.n271 0.155672
R478 drain_right.n271 drain_right.n159 0.155672
R479 drain_right.n263 drain_right.n159 0.155672
R480 drain_right.n263 drain_right.n262 0.155672
R481 drain_right.n262 drain_right.n163 0.155672
R482 drain_right.n255 drain_right.n163 0.155672
R483 drain_right.n255 drain_right.n254 0.155672
R484 drain_right.n254 drain_right.n168 0.155672
R485 drain_right.n247 drain_right.n168 0.155672
R486 drain_right.n247 drain_right.n246 0.155672
R487 drain_right.n246 drain_right.n172 0.155672
R488 drain_right.n239 drain_right.n172 0.155672
R489 drain_right.n239 drain_right.n238 0.155672
R490 drain_right.n238 drain_right.n176 0.155672
R491 drain_right.n231 drain_right.n176 0.155672
R492 drain_right.n231 drain_right.n230 0.155672
R493 drain_right.n230 drain_right.n180 0.155672
R494 drain_right.n223 drain_right.n180 0.155672
R495 drain_right.n223 drain_right.n222 0.155672
R496 drain_right.n222 drain_right.n184 0.155672
R497 drain_right.n214 drain_right.n184 0.155672
R498 drain_right.n214 drain_right.n213 0.155672
R499 drain_right.n213 drain_right.n189 0.155672
R500 drain_right.n206 drain_right.n189 0.155672
R501 drain_right.n206 drain_right.n205 0.155672
R502 drain_right.n205 drain_right.n193 0.155672
R503 drain_right.n198 drain_right.n193 0.155672
R504 drain_right.n144 drain_right.n143 0.0809298
R505 source.n578 source.n444 289.615
R506 source.n432 source.n298 289.615
R507 source.n134 source.n0 289.615
R508 source.n280 source.n146 289.615
R509 source.n488 source.n487 185
R510 source.n493 source.n492 185
R511 source.n495 source.n494 185
R512 source.n484 source.n483 185
R513 source.n501 source.n500 185
R514 source.n503 source.n502 185
R515 source.n480 source.n479 185
R516 source.n510 source.n509 185
R517 source.n511 source.n478 185
R518 source.n513 source.n512 185
R519 source.n476 source.n475 185
R520 source.n519 source.n518 185
R521 source.n521 source.n520 185
R522 source.n472 source.n471 185
R523 source.n527 source.n526 185
R524 source.n529 source.n528 185
R525 source.n468 source.n467 185
R526 source.n535 source.n534 185
R527 source.n537 source.n536 185
R528 source.n464 source.n463 185
R529 source.n543 source.n542 185
R530 source.n545 source.n544 185
R531 source.n460 source.n459 185
R532 source.n551 source.n550 185
R533 source.n554 source.n553 185
R534 source.n552 source.n456 185
R535 source.n559 source.n455 185
R536 source.n561 source.n560 185
R537 source.n563 source.n562 185
R538 source.n452 source.n451 185
R539 source.n569 source.n568 185
R540 source.n571 source.n570 185
R541 source.n448 source.n447 185
R542 source.n577 source.n576 185
R543 source.n579 source.n578 185
R544 source.n342 source.n341 185
R545 source.n347 source.n346 185
R546 source.n349 source.n348 185
R547 source.n338 source.n337 185
R548 source.n355 source.n354 185
R549 source.n357 source.n356 185
R550 source.n334 source.n333 185
R551 source.n364 source.n363 185
R552 source.n365 source.n332 185
R553 source.n367 source.n366 185
R554 source.n330 source.n329 185
R555 source.n373 source.n372 185
R556 source.n375 source.n374 185
R557 source.n326 source.n325 185
R558 source.n381 source.n380 185
R559 source.n383 source.n382 185
R560 source.n322 source.n321 185
R561 source.n389 source.n388 185
R562 source.n391 source.n390 185
R563 source.n318 source.n317 185
R564 source.n397 source.n396 185
R565 source.n399 source.n398 185
R566 source.n314 source.n313 185
R567 source.n405 source.n404 185
R568 source.n408 source.n407 185
R569 source.n406 source.n310 185
R570 source.n413 source.n309 185
R571 source.n415 source.n414 185
R572 source.n417 source.n416 185
R573 source.n306 source.n305 185
R574 source.n423 source.n422 185
R575 source.n425 source.n424 185
R576 source.n302 source.n301 185
R577 source.n431 source.n430 185
R578 source.n433 source.n432 185
R579 source.n135 source.n134 185
R580 source.n133 source.n132 185
R581 source.n4 source.n3 185
R582 source.n127 source.n126 185
R583 source.n125 source.n124 185
R584 source.n8 source.n7 185
R585 source.n119 source.n118 185
R586 source.n117 source.n116 185
R587 source.n115 source.n11 185
R588 source.n15 source.n12 185
R589 source.n110 source.n109 185
R590 source.n108 source.n107 185
R591 source.n17 source.n16 185
R592 source.n102 source.n101 185
R593 source.n100 source.n99 185
R594 source.n21 source.n20 185
R595 source.n94 source.n93 185
R596 source.n92 source.n91 185
R597 source.n25 source.n24 185
R598 source.n86 source.n85 185
R599 source.n84 source.n83 185
R600 source.n29 source.n28 185
R601 source.n78 source.n77 185
R602 source.n76 source.n75 185
R603 source.n33 source.n32 185
R604 source.n70 source.n69 185
R605 source.n68 source.n35 185
R606 source.n67 source.n66 185
R607 source.n38 source.n36 185
R608 source.n61 source.n60 185
R609 source.n59 source.n58 185
R610 source.n42 source.n41 185
R611 source.n53 source.n52 185
R612 source.n51 source.n50 185
R613 source.n46 source.n45 185
R614 source.n281 source.n280 185
R615 source.n279 source.n278 185
R616 source.n150 source.n149 185
R617 source.n273 source.n272 185
R618 source.n271 source.n270 185
R619 source.n154 source.n153 185
R620 source.n265 source.n264 185
R621 source.n263 source.n262 185
R622 source.n261 source.n157 185
R623 source.n161 source.n158 185
R624 source.n256 source.n255 185
R625 source.n254 source.n253 185
R626 source.n163 source.n162 185
R627 source.n248 source.n247 185
R628 source.n246 source.n245 185
R629 source.n167 source.n166 185
R630 source.n240 source.n239 185
R631 source.n238 source.n237 185
R632 source.n171 source.n170 185
R633 source.n232 source.n231 185
R634 source.n230 source.n229 185
R635 source.n175 source.n174 185
R636 source.n224 source.n223 185
R637 source.n222 source.n221 185
R638 source.n179 source.n178 185
R639 source.n216 source.n215 185
R640 source.n214 source.n181 185
R641 source.n213 source.n212 185
R642 source.n184 source.n182 185
R643 source.n207 source.n206 185
R644 source.n205 source.n204 185
R645 source.n188 source.n187 185
R646 source.n199 source.n198 185
R647 source.n197 source.n196 185
R648 source.n192 source.n191 185
R649 source.n489 source.t22 149.524
R650 source.n343 source.t3 149.524
R651 source.n47 source.t8 149.524
R652 source.n193 source.t19 149.524
R653 source.n493 source.n487 104.615
R654 source.n494 source.n493 104.615
R655 source.n494 source.n483 104.615
R656 source.n501 source.n483 104.615
R657 source.n502 source.n501 104.615
R658 source.n502 source.n479 104.615
R659 source.n510 source.n479 104.615
R660 source.n511 source.n510 104.615
R661 source.n512 source.n511 104.615
R662 source.n512 source.n475 104.615
R663 source.n519 source.n475 104.615
R664 source.n520 source.n519 104.615
R665 source.n520 source.n471 104.615
R666 source.n527 source.n471 104.615
R667 source.n528 source.n527 104.615
R668 source.n528 source.n467 104.615
R669 source.n535 source.n467 104.615
R670 source.n536 source.n535 104.615
R671 source.n536 source.n463 104.615
R672 source.n543 source.n463 104.615
R673 source.n544 source.n543 104.615
R674 source.n544 source.n459 104.615
R675 source.n551 source.n459 104.615
R676 source.n553 source.n551 104.615
R677 source.n553 source.n552 104.615
R678 source.n552 source.n455 104.615
R679 source.n561 source.n455 104.615
R680 source.n562 source.n561 104.615
R681 source.n562 source.n451 104.615
R682 source.n569 source.n451 104.615
R683 source.n570 source.n569 104.615
R684 source.n570 source.n447 104.615
R685 source.n577 source.n447 104.615
R686 source.n578 source.n577 104.615
R687 source.n347 source.n341 104.615
R688 source.n348 source.n347 104.615
R689 source.n348 source.n337 104.615
R690 source.n355 source.n337 104.615
R691 source.n356 source.n355 104.615
R692 source.n356 source.n333 104.615
R693 source.n364 source.n333 104.615
R694 source.n365 source.n364 104.615
R695 source.n366 source.n365 104.615
R696 source.n366 source.n329 104.615
R697 source.n373 source.n329 104.615
R698 source.n374 source.n373 104.615
R699 source.n374 source.n325 104.615
R700 source.n381 source.n325 104.615
R701 source.n382 source.n381 104.615
R702 source.n382 source.n321 104.615
R703 source.n389 source.n321 104.615
R704 source.n390 source.n389 104.615
R705 source.n390 source.n317 104.615
R706 source.n397 source.n317 104.615
R707 source.n398 source.n397 104.615
R708 source.n398 source.n313 104.615
R709 source.n405 source.n313 104.615
R710 source.n407 source.n405 104.615
R711 source.n407 source.n406 104.615
R712 source.n406 source.n309 104.615
R713 source.n415 source.n309 104.615
R714 source.n416 source.n415 104.615
R715 source.n416 source.n305 104.615
R716 source.n423 source.n305 104.615
R717 source.n424 source.n423 104.615
R718 source.n424 source.n301 104.615
R719 source.n431 source.n301 104.615
R720 source.n432 source.n431 104.615
R721 source.n134 source.n133 104.615
R722 source.n133 source.n3 104.615
R723 source.n126 source.n3 104.615
R724 source.n126 source.n125 104.615
R725 source.n125 source.n7 104.615
R726 source.n118 source.n7 104.615
R727 source.n118 source.n117 104.615
R728 source.n117 source.n11 104.615
R729 source.n15 source.n11 104.615
R730 source.n109 source.n15 104.615
R731 source.n109 source.n108 104.615
R732 source.n108 source.n16 104.615
R733 source.n101 source.n16 104.615
R734 source.n101 source.n100 104.615
R735 source.n100 source.n20 104.615
R736 source.n93 source.n20 104.615
R737 source.n93 source.n92 104.615
R738 source.n92 source.n24 104.615
R739 source.n85 source.n24 104.615
R740 source.n85 source.n84 104.615
R741 source.n84 source.n28 104.615
R742 source.n77 source.n28 104.615
R743 source.n77 source.n76 104.615
R744 source.n76 source.n32 104.615
R745 source.n69 source.n32 104.615
R746 source.n69 source.n68 104.615
R747 source.n68 source.n67 104.615
R748 source.n67 source.n36 104.615
R749 source.n60 source.n36 104.615
R750 source.n60 source.n59 104.615
R751 source.n59 source.n41 104.615
R752 source.n52 source.n41 104.615
R753 source.n52 source.n51 104.615
R754 source.n51 source.n45 104.615
R755 source.n280 source.n279 104.615
R756 source.n279 source.n149 104.615
R757 source.n272 source.n149 104.615
R758 source.n272 source.n271 104.615
R759 source.n271 source.n153 104.615
R760 source.n264 source.n153 104.615
R761 source.n264 source.n263 104.615
R762 source.n263 source.n157 104.615
R763 source.n161 source.n157 104.615
R764 source.n255 source.n161 104.615
R765 source.n255 source.n254 104.615
R766 source.n254 source.n162 104.615
R767 source.n247 source.n162 104.615
R768 source.n247 source.n246 104.615
R769 source.n246 source.n166 104.615
R770 source.n239 source.n166 104.615
R771 source.n239 source.n238 104.615
R772 source.n238 source.n170 104.615
R773 source.n231 source.n170 104.615
R774 source.n231 source.n230 104.615
R775 source.n230 source.n174 104.615
R776 source.n223 source.n174 104.615
R777 source.n223 source.n222 104.615
R778 source.n222 source.n178 104.615
R779 source.n215 source.n178 104.615
R780 source.n215 source.n214 104.615
R781 source.n214 source.n213 104.615
R782 source.n213 source.n182 104.615
R783 source.n206 source.n182 104.615
R784 source.n206 source.n205 104.615
R785 source.n205 source.n187 104.615
R786 source.n198 source.n187 104.615
R787 source.n198 source.n197 104.615
R788 source.n197 source.n191 104.615
R789 source.t22 source.n487 52.3082
R790 source.t3 source.n341 52.3082
R791 source.t8 source.n45 52.3082
R792 source.t19 source.n191 52.3082
R793 source.n443 source.n442 42.0366
R794 source.n441 source.n440 42.0366
R795 source.n439 source.n438 42.0366
R796 source.n297 source.n296 42.0366
R797 source.n295 source.n294 42.0366
R798 source.n293 source.n292 42.0366
R799 source.n141 source.n140 42.0366
R800 source.n143 source.n142 42.0366
R801 source.n145 source.n144 42.0366
R802 source.n287 source.n286 42.0366
R803 source.n289 source.n288 42.0366
R804 source.n291 source.n290 42.0366
R805 source.n293 source.n291 32.2224
R806 source.n583 source.n582 30.6338
R807 source.n437 source.n436 30.6338
R808 source.n139 source.n138 30.6338
R809 source.n285 source.n284 30.6338
R810 source.n584 source.n139 26.1448
R811 source.n513 source.n478 13.1884
R812 source.n560 source.n559 13.1884
R813 source.n367 source.n332 13.1884
R814 source.n414 source.n413 13.1884
R815 source.n116 source.n115 13.1884
R816 source.n70 source.n35 13.1884
R817 source.n262 source.n261 13.1884
R818 source.n216 source.n181 13.1884
R819 source.n509 source.n508 12.8005
R820 source.n514 source.n476 12.8005
R821 source.n558 source.n456 12.8005
R822 source.n563 source.n454 12.8005
R823 source.n363 source.n362 12.8005
R824 source.n368 source.n330 12.8005
R825 source.n412 source.n310 12.8005
R826 source.n417 source.n308 12.8005
R827 source.n119 source.n10 12.8005
R828 source.n114 source.n12 12.8005
R829 source.n71 source.n33 12.8005
R830 source.n66 source.n37 12.8005
R831 source.n265 source.n156 12.8005
R832 source.n260 source.n158 12.8005
R833 source.n217 source.n179 12.8005
R834 source.n212 source.n183 12.8005
R835 source.n507 source.n480 12.0247
R836 source.n518 source.n517 12.0247
R837 source.n555 source.n554 12.0247
R838 source.n564 source.n452 12.0247
R839 source.n361 source.n334 12.0247
R840 source.n372 source.n371 12.0247
R841 source.n409 source.n408 12.0247
R842 source.n418 source.n306 12.0247
R843 source.n120 source.n8 12.0247
R844 source.n111 source.n110 12.0247
R845 source.n75 source.n74 12.0247
R846 source.n65 source.n38 12.0247
R847 source.n266 source.n154 12.0247
R848 source.n257 source.n256 12.0247
R849 source.n221 source.n220 12.0247
R850 source.n211 source.n184 12.0247
R851 source.n504 source.n503 11.249
R852 source.n521 source.n474 11.249
R853 source.n550 source.n458 11.249
R854 source.n568 source.n567 11.249
R855 source.n358 source.n357 11.249
R856 source.n375 source.n328 11.249
R857 source.n404 source.n312 11.249
R858 source.n422 source.n421 11.249
R859 source.n124 source.n123 11.249
R860 source.n107 source.n14 11.249
R861 source.n78 source.n31 11.249
R862 source.n62 source.n61 11.249
R863 source.n270 source.n269 11.249
R864 source.n253 source.n160 11.249
R865 source.n224 source.n177 11.249
R866 source.n208 source.n207 11.249
R867 source.n500 source.n482 10.4732
R868 source.n522 source.n472 10.4732
R869 source.n549 source.n460 10.4732
R870 source.n571 source.n450 10.4732
R871 source.n354 source.n336 10.4732
R872 source.n376 source.n326 10.4732
R873 source.n403 source.n314 10.4732
R874 source.n425 source.n304 10.4732
R875 source.n127 source.n6 10.4732
R876 source.n106 source.n17 10.4732
R877 source.n79 source.n29 10.4732
R878 source.n58 source.n40 10.4732
R879 source.n273 source.n152 10.4732
R880 source.n252 source.n163 10.4732
R881 source.n225 source.n175 10.4732
R882 source.n204 source.n186 10.4732
R883 source.n489 source.n488 10.2747
R884 source.n343 source.n342 10.2747
R885 source.n47 source.n46 10.2747
R886 source.n193 source.n192 10.2747
R887 source.n499 source.n484 9.69747
R888 source.n526 source.n525 9.69747
R889 source.n546 source.n545 9.69747
R890 source.n572 source.n448 9.69747
R891 source.n353 source.n338 9.69747
R892 source.n380 source.n379 9.69747
R893 source.n400 source.n399 9.69747
R894 source.n426 source.n302 9.69747
R895 source.n128 source.n4 9.69747
R896 source.n103 source.n102 9.69747
R897 source.n83 source.n82 9.69747
R898 source.n57 source.n42 9.69747
R899 source.n274 source.n150 9.69747
R900 source.n249 source.n248 9.69747
R901 source.n229 source.n228 9.69747
R902 source.n203 source.n188 9.69747
R903 source.n582 source.n581 9.45567
R904 source.n436 source.n435 9.45567
R905 source.n138 source.n137 9.45567
R906 source.n284 source.n283 9.45567
R907 source.n446 source.n445 9.3005
R908 source.n575 source.n574 9.3005
R909 source.n573 source.n572 9.3005
R910 source.n450 source.n449 9.3005
R911 source.n567 source.n566 9.3005
R912 source.n565 source.n564 9.3005
R913 source.n454 source.n453 9.3005
R914 source.n533 source.n532 9.3005
R915 source.n531 source.n530 9.3005
R916 source.n470 source.n469 9.3005
R917 source.n525 source.n524 9.3005
R918 source.n523 source.n522 9.3005
R919 source.n474 source.n473 9.3005
R920 source.n517 source.n516 9.3005
R921 source.n515 source.n514 9.3005
R922 source.n491 source.n490 9.3005
R923 source.n486 source.n485 9.3005
R924 source.n497 source.n496 9.3005
R925 source.n499 source.n498 9.3005
R926 source.n482 source.n481 9.3005
R927 source.n505 source.n504 9.3005
R928 source.n507 source.n506 9.3005
R929 source.n508 source.n477 9.3005
R930 source.n466 source.n465 9.3005
R931 source.n539 source.n538 9.3005
R932 source.n541 source.n540 9.3005
R933 source.n462 source.n461 9.3005
R934 source.n547 source.n546 9.3005
R935 source.n549 source.n548 9.3005
R936 source.n458 source.n457 9.3005
R937 source.n556 source.n555 9.3005
R938 source.n558 source.n557 9.3005
R939 source.n581 source.n580 9.3005
R940 source.n300 source.n299 9.3005
R941 source.n429 source.n428 9.3005
R942 source.n427 source.n426 9.3005
R943 source.n304 source.n303 9.3005
R944 source.n421 source.n420 9.3005
R945 source.n419 source.n418 9.3005
R946 source.n308 source.n307 9.3005
R947 source.n387 source.n386 9.3005
R948 source.n385 source.n384 9.3005
R949 source.n324 source.n323 9.3005
R950 source.n379 source.n378 9.3005
R951 source.n377 source.n376 9.3005
R952 source.n328 source.n327 9.3005
R953 source.n371 source.n370 9.3005
R954 source.n369 source.n368 9.3005
R955 source.n345 source.n344 9.3005
R956 source.n340 source.n339 9.3005
R957 source.n351 source.n350 9.3005
R958 source.n353 source.n352 9.3005
R959 source.n336 source.n335 9.3005
R960 source.n359 source.n358 9.3005
R961 source.n361 source.n360 9.3005
R962 source.n362 source.n331 9.3005
R963 source.n320 source.n319 9.3005
R964 source.n393 source.n392 9.3005
R965 source.n395 source.n394 9.3005
R966 source.n316 source.n315 9.3005
R967 source.n401 source.n400 9.3005
R968 source.n403 source.n402 9.3005
R969 source.n312 source.n311 9.3005
R970 source.n410 source.n409 9.3005
R971 source.n412 source.n411 9.3005
R972 source.n435 source.n434 9.3005
R973 source.n49 source.n48 9.3005
R974 source.n44 source.n43 9.3005
R975 source.n55 source.n54 9.3005
R976 source.n57 source.n56 9.3005
R977 source.n40 source.n39 9.3005
R978 source.n63 source.n62 9.3005
R979 source.n65 source.n64 9.3005
R980 source.n37 source.n34 9.3005
R981 source.n96 source.n95 9.3005
R982 source.n98 source.n97 9.3005
R983 source.n19 source.n18 9.3005
R984 source.n104 source.n103 9.3005
R985 source.n106 source.n105 9.3005
R986 source.n14 source.n13 9.3005
R987 source.n112 source.n111 9.3005
R988 source.n114 source.n113 9.3005
R989 source.n137 source.n136 9.3005
R990 source.n2 source.n1 9.3005
R991 source.n131 source.n130 9.3005
R992 source.n129 source.n128 9.3005
R993 source.n6 source.n5 9.3005
R994 source.n123 source.n122 9.3005
R995 source.n121 source.n120 9.3005
R996 source.n10 source.n9 9.3005
R997 source.n23 source.n22 9.3005
R998 source.n90 source.n89 9.3005
R999 source.n88 source.n87 9.3005
R1000 source.n27 source.n26 9.3005
R1001 source.n82 source.n81 9.3005
R1002 source.n80 source.n79 9.3005
R1003 source.n31 source.n30 9.3005
R1004 source.n74 source.n73 9.3005
R1005 source.n72 source.n71 9.3005
R1006 source.n195 source.n194 9.3005
R1007 source.n190 source.n189 9.3005
R1008 source.n201 source.n200 9.3005
R1009 source.n203 source.n202 9.3005
R1010 source.n186 source.n185 9.3005
R1011 source.n209 source.n208 9.3005
R1012 source.n211 source.n210 9.3005
R1013 source.n183 source.n180 9.3005
R1014 source.n242 source.n241 9.3005
R1015 source.n244 source.n243 9.3005
R1016 source.n165 source.n164 9.3005
R1017 source.n250 source.n249 9.3005
R1018 source.n252 source.n251 9.3005
R1019 source.n160 source.n159 9.3005
R1020 source.n258 source.n257 9.3005
R1021 source.n260 source.n259 9.3005
R1022 source.n283 source.n282 9.3005
R1023 source.n148 source.n147 9.3005
R1024 source.n277 source.n276 9.3005
R1025 source.n275 source.n274 9.3005
R1026 source.n152 source.n151 9.3005
R1027 source.n269 source.n268 9.3005
R1028 source.n267 source.n266 9.3005
R1029 source.n156 source.n155 9.3005
R1030 source.n169 source.n168 9.3005
R1031 source.n236 source.n235 9.3005
R1032 source.n234 source.n233 9.3005
R1033 source.n173 source.n172 9.3005
R1034 source.n228 source.n227 9.3005
R1035 source.n226 source.n225 9.3005
R1036 source.n177 source.n176 9.3005
R1037 source.n220 source.n219 9.3005
R1038 source.n218 source.n217 9.3005
R1039 source.n496 source.n495 8.92171
R1040 source.n529 source.n470 8.92171
R1041 source.n542 source.n462 8.92171
R1042 source.n576 source.n575 8.92171
R1043 source.n350 source.n349 8.92171
R1044 source.n383 source.n324 8.92171
R1045 source.n396 source.n316 8.92171
R1046 source.n430 source.n429 8.92171
R1047 source.n132 source.n131 8.92171
R1048 source.n99 source.n19 8.92171
R1049 source.n86 source.n27 8.92171
R1050 source.n54 source.n53 8.92171
R1051 source.n278 source.n277 8.92171
R1052 source.n245 source.n165 8.92171
R1053 source.n232 source.n173 8.92171
R1054 source.n200 source.n199 8.92171
R1055 source.n492 source.n486 8.14595
R1056 source.n530 source.n468 8.14595
R1057 source.n541 source.n464 8.14595
R1058 source.n579 source.n446 8.14595
R1059 source.n346 source.n340 8.14595
R1060 source.n384 source.n322 8.14595
R1061 source.n395 source.n318 8.14595
R1062 source.n433 source.n300 8.14595
R1063 source.n135 source.n2 8.14595
R1064 source.n98 source.n21 8.14595
R1065 source.n87 source.n25 8.14595
R1066 source.n50 source.n44 8.14595
R1067 source.n281 source.n148 8.14595
R1068 source.n244 source.n167 8.14595
R1069 source.n233 source.n171 8.14595
R1070 source.n196 source.n190 8.14595
R1071 source.n491 source.n488 7.3702
R1072 source.n534 source.n533 7.3702
R1073 source.n538 source.n537 7.3702
R1074 source.n580 source.n444 7.3702
R1075 source.n345 source.n342 7.3702
R1076 source.n388 source.n387 7.3702
R1077 source.n392 source.n391 7.3702
R1078 source.n434 source.n298 7.3702
R1079 source.n136 source.n0 7.3702
R1080 source.n95 source.n94 7.3702
R1081 source.n91 source.n90 7.3702
R1082 source.n49 source.n46 7.3702
R1083 source.n282 source.n146 7.3702
R1084 source.n241 source.n240 7.3702
R1085 source.n237 source.n236 7.3702
R1086 source.n195 source.n192 7.3702
R1087 source.n534 source.n466 6.59444
R1088 source.n537 source.n466 6.59444
R1089 source.n582 source.n444 6.59444
R1090 source.n388 source.n320 6.59444
R1091 source.n391 source.n320 6.59444
R1092 source.n436 source.n298 6.59444
R1093 source.n138 source.n0 6.59444
R1094 source.n94 source.n23 6.59444
R1095 source.n91 source.n23 6.59444
R1096 source.n284 source.n146 6.59444
R1097 source.n240 source.n169 6.59444
R1098 source.n237 source.n169 6.59444
R1099 source.n492 source.n491 5.81868
R1100 source.n533 source.n468 5.81868
R1101 source.n538 source.n464 5.81868
R1102 source.n580 source.n579 5.81868
R1103 source.n346 source.n345 5.81868
R1104 source.n387 source.n322 5.81868
R1105 source.n392 source.n318 5.81868
R1106 source.n434 source.n433 5.81868
R1107 source.n136 source.n135 5.81868
R1108 source.n95 source.n21 5.81868
R1109 source.n90 source.n25 5.81868
R1110 source.n50 source.n49 5.81868
R1111 source.n282 source.n281 5.81868
R1112 source.n241 source.n167 5.81868
R1113 source.n236 source.n171 5.81868
R1114 source.n196 source.n195 5.81868
R1115 source.n584 source.n583 5.53498
R1116 source.n495 source.n486 5.04292
R1117 source.n530 source.n529 5.04292
R1118 source.n542 source.n541 5.04292
R1119 source.n576 source.n446 5.04292
R1120 source.n349 source.n340 5.04292
R1121 source.n384 source.n383 5.04292
R1122 source.n396 source.n395 5.04292
R1123 source.n430 source.n300 5.04292
R1124 source.n132 source.n2 5.04292
R1125 source.n99 source.n98 5.04292
R1126 source.n87 source.n86 5.04292
R1127 source.n53 source.n44 5.04292
R1128 source.n278 source.n148 5.04292
R1129 source.n245 source.n244 5.04292
R1130 source.n233 source.n232 5.04292
R1131 source.n199 source.n190 5.04292
R1132 source.n496 source.n484 4.26717
R1133 source.n526 source.n470 4.26717
R1134 source.n545 source.n462 4.26717
R1135 source.n575 source.n448 4.26717
R1136 source.n350 source.n338 4.26717
R1137 source.n380 source.n324 4.26717
R1138 source.n399 source.n316 4.26717
R1139 source.n429 source.n302 4.26717
R1140 source.n131 source.n4 4.26717
R1141 source.n102 source.n19 4.26717
R1142 source.n83 source.n27 4.26717
R1143 source.n54 source.n42 4.26717
R1144 source.n277 source.n150 4.26717
R1145 source.n248 source.n165 4.26717
R1146 source.n229 source.n173 4.26717
R1147 source.n200 source.n188 4.26717
R1148 source.n500 source.n499 3.49141
R1149 source.n525 source.n472 3.49141
R1150 source.n546 source.n460 3.49141
R1151 source.n572 source.n571 3.49141
R1152 source.n354 source.n353 3.49141
R1153 source.n379 source.n326 3.49141
R1154 source.n400 source.n314 3.49141
R1155 source.n426 source.n425 3.49141
R1156 source.n128 source.n127 3.49141
R1157 source.n103 source.n17 3.49141
R1158 source.n82 source.n29 3.49141
R1159 source.n58 source.n57 3.49141
R1160 source.n274 source.n273 3.49141
R1161 source.n249 source.n163 3.49141
R1162 source.n228 source.n175 3.49141
R1163 source.n204 source.n203 3.49141
R1164 source.n48 source.n47 2.84303
R1165 source.n194 source.n193 2.84303
R1166 source.n490 source.n489 2.84303
R1167 source.n344 source.n343 2.84303
R1168 source.n503 source.n482 2.71565
R1169 source.n522 source.n521 2.71565
R1170 source.n550 source.n549 2.71565
R1171 source.n568 source.n450 2.71565
R1172 source.n357 source.n336 2.71565
R1173 source.n376 source.n375 2.71565
R1174 source.n404 source.n403 2.71565
R1175 source.n422 source.n304 2.71565
R1176 source.n124 source.n6 2.71565
R1177 source.n107 source.n106 2.71565
R1178 source.n79 source.n78 2.71565
R1179 source.n61 source.n40 2.71565
R1180 source.n270 source.n152 2.71565
R1181 source.n253 source.n252 2.71565
R1182 source.n225 source.n224 2.71565
R1183 source.n207 source.n186 2.71565
R1184 source.n504 source.n480 1.93989
R1185 source.n518 source.n474 1.93989
R1186 source.n554 source.n458 1.93989
R1187 source.n567 source.n452 1.93989
R1188 source.n358 source.n334 1.93989
R1189 source.n372 source.n328 1.93989
R1190 source.n408 source.n312 1.93989
R1191 source.n421 source.n306 1.93989
R1192 source.n123 source.n8 1.93989
R1193 source.n110 source.n14 1.93989
R1194 source.n75 source.n31 1.93989
R1195 source.n62 source.n38 1.93989
R1196 source.n269 source.n154 1.93989
R1197 source.n256 source.n160 1.93989
R1198 source.n221 source.n177 1.93989
R1199 source.n208 source.n184 1.93989
R1200 source.n509 source.n507 1.16414
R1201 source.n517 source.n476 1.16414
R1202 source.n555 source.n456 1.16414
R1203 source.n564 source.n563 1.16414
R1204 source.n363 source.n361 1.16414
R1205 source.n371 source.n330 1.16414
R1206 source.n409 source.n310 1.16414
R1207 source.n418 source.n417 1.16414
R1208 source.n120 source.n119 1.16414
R1209 source.n111 source.n12 1.16414
R1210 source.n74 source.n33 1.16414
R1211 source.n66 source.n65 1.16414
R1212 source.n266 source.n265 1.16414
R1213 source.n257 source.n158 1.16414
R1214 source.n220 source.n179 1.16414
R1215 source.n212 source.n211 1.16414
R1216 source.n442 source.t21 0.7925
R1217 source.n442 source.t14 0.7925
R1218 source.n440 source.t25 0.7925
R1219 source.n440 source.t18 0.7925
R1220 source.n438 source.t24 0.7925
R1221 source.n438 source.t17 0.7925
R1222 source.n296 source.t9 0.7925
R1223 source.n296 source.t10 0.7925
R1224 source.n294 source.t2 0.7925
R1225 source.n294 source.t12 0.7925
R1226 source.n292 source.t0 0.7925
R1227 source.n292 source.t5 0.7925
R1228 source.n140 source.t1 0.7925
R1229 source.n140 source.t6 0.7925
R1230 source.n142 source.t13 0.7925
R1231 source.n142 source.t11 0.7925
R1232 source.n144 source.t7 0.7925
R1233 source.n144 source.t4 0.7925
R1234 source.n286 source.t26 0.7925
R1235 source.n286 source.t15 0.7925
R1236 source.n288 source.t16 0.7925
R1237 source.n288 source.t20 0.7925
R1238 source.n290 source.t23 0.7925
R1239 source.n290 source.t27 0.7925
R1240 source.n285 source.n145 0.741879
R1241 source.n439 source.n437 0.741879
R1242 source.n291 source.n289 0.543603
R1243 source.n289 source.n287 0.543603
R1244 source.n287 source.n285 0.543603
R1245 source.n145 source.n143 0.543603
R1246 source.n143 source.n141 0.543603
R1247 source.n141 source.n139 0.543603
R1248 source.n295 source.n293 0.543603
R1249 source.n297 source.n295 0.543603
R1250 source.n437 source.n297 0.543603
R1251 source.n441 source.n439 0.543603
R1252 source.n443 source.n441 0.543603
R1253 source.n583 source.n443 0.543603
R1254 source.n508 source.n478 0.388379
R1255 source.n514 source.n513 0.388379
R1256 source.n559 source.n558 0.388379
R1257 source.n560 source.n454 0.388379
R1258 source.n362 source.n332 0.388379
R1259 source.n368 source.n367 0.388379
R1260 source.n413 source.n412 0.388379
R1261 source.n414 source.n308 0.388379
R1262 source.n116 source.n10 0.388379
R1263 source.n115 source.n114 0.388379
R1264 source.n71 source.n70 0.388379
R1265 source.n37 source.n35 0.388379
R1266 source.n262 source.n156 0.388379
R1267 source.n261 source.n260 0.388379
R1268 source.n217 source.n216 0.388379
R1269 source.n183 source.n181 0.388379
R1270 source source.n584 0.188
R1271 source.n490 source.n485 0.155672
R1272 source.n497 source.n485 0.155672
R1273 source.n498 source.n497 0.155672
R1274 source.n498 source.n481 0.155672
R1275 source.n505 source.n481 0.155672
R1276 source.n506 source.n505 0.155672
R1277 source.n506 source.n477 0.155672
R1278 source.n515 source.n477 0.155672
R1279 source.n516 source.n515 0.155672
R1280 source.n516 source.n473 0.155672
R1281 source.n523 source.n473 0.155672
R1282 source.n524 source.n523 0.155672
R1283 source.n524 source.n469 0.155672
R1284 source.n531 source.n469 0.155672
R1285 source.n532 source.n531 0.155672
R1286 source.n532 source.n465 0.155672
R1287 source.n539 source.n465 0.155672
R1288 source.n540 source.n539 0.155672
R1289 source.n540 source.n461 0.155672
R1290 source.n547 source.n461 0.155672
R1291 source.n548 source.n547 0.155672
R1292 source.n548 source.n457 0.155672
R1293 source.n556 source.n457 0.155672
R1294 source.n557 source.n556 0.155672
R1295 source.n557 source.n453 0.155672
R1296 source.n565 source.n453 0.155672
R1297 source.n566 source.n565 0.155672
R1298 source.n566 source.n449 0.155672
R1299 source.n573 source.n449 0.155672
R1300 source.n574 source.n573 0.155672
R1301 source.n574 source.n445 0.155672
R1302 source.n581 source.n445 0.155672
R1303 source.n344 source.n339 0.155672
R1304 source.n351 source.n339 0.155672
R1305 source.n352 source.n351 0.155672
R1306 source.n352 source.n335 0.155672
R1307 source.n359 source.n335 0.155672
R1308 source.n360 source.n359 0.155672
R1309 source.n360 source.n331 0.155672
R1310 source.n369 source.n331 0.155672
R1311 source.n370 source.n369 0.155672
R1312 source.n370 source.n327 0.155672
R1313 source.n377 source.n327 0.155672
R1314 source.n378 source.n377 0.155672
R1315 source.n378 source.n323 0.155672
R1316 source.n385 source.n323 0.155672
R1317 source.n386 source.n385 0.155672
R1318 source.n386 source.n319 0.155672
R1319 source.n393 source.n319 0.155672
R1320 source.n394 source.n393 0.155672
R1321 source.n394 source.n315 0.155672
R1322 source.n401 source.n315 0.155672
R1323 source.n402 source.n401 0.155672
R1324 source.n402 source.n311 0.155672
R1325 source.n410 source.n311 0.155672
R1326 source.n411 source.n410 0.155672
R1327 source.n411 source.n307 0.155672
R1328 source.n419 source.n307 0.155672
R1329 source.n420 source.n419 0.155672
R1330 source.n420 source.n303 0.155672
R1331 source.n427 source.n303 0.155672
R1332 source.n428 source.n427 0.155672
R1333 source.n428 source.n299 0.155672
R1334 source.n435 source.n299 0.155672
R1335 source.n137 source.n1 0.155672
R1336 source.n130 source.n1 0.155672
R1337 source.n130 source.n129 0.155672
R1338 source.n129 source.n5 0.155672
R1339 source.n122 source.n5 0.155672
R1340 source.n122 source.n121 0.155672
R1341 source.n121 source.n9 0.155672
R1342 source.n113 source.n9 0.155672
R1343 source.n113 source.n112 0.155672
R1344 source.n112 source.n13 0.155672
R1345 source.n105 source.n13 0.155672
R1346 source.n105 source.n104 0.155672
R1347 source.n104 source.n18 0.155672
R1348 source.n97 source.n18 0.155672
R1349 source.n97 source.n96 0.155672
R1350 source.n96 source.n22 0.155672
R1351 source.n89 source.n22 0.155672
R1352 source.n89 source.n88 0.155672
R1353 source.n88 source.n26 0.155672
R1354 source.n81 source.n26 0.155672
R1355 source.n81 source.n80 0.155672
R1356 source.n80 source.n30 0.155672
R1357 source.n73 source.n30 0.155672
R1358 source.n73 source.n72 0.155672
R1359 source.n72 source.n34 0.155672
R1360 source.n64 source.n34 0.155672
R1361 source.n64 source.n63 0.155672
R1362 source.n63 source.n39 0.155672
R1363 source.n56 source.n39 0.155672
R1364 source.n56 source.n55 0.155672
R1365 source.n55 source.n43 0.155672
R1366 source.n48 source.n43 0.155672
R1367 source.n283 source.n147 0.155672
R1368 source.n276 source.n147 0.155672
R1369 source.n276 source.n275 0.155672
R1370 source.n275 source.n151 0.155672
R1371 source.n268 source.n151 0.155672
R1372 source.n268 source.n267 0.155672
R1373 source.n267 source.n155 0.155672
R1374 source.n259 source.n155 0.155672
R1375 source.n259 source.n258 0.155672
R1376 source.n258 source.n159 0.155672
R1377 source.n251 source.n159 0.155672
R1378 source.n251 source.n250 0.155672
R1379 source.n250 source.n164 0.155672
R1380 source.n243 source.n164 0.155672
R1381 source.n243 source.n242 0.155672
R1382 source.n242 source.n168 0.155672
R1383 source.n235 source.n168 0.155672
R1384 source.n235 source.n234 0.155672
R1385 source.n234 source.n172 0.155672
R1386 source.n227 source.n172 0.155672
R1387 source.n227 source.n226 0.155672
R1388 source.n226 source.n176 0.155672
R1389 source.n219 source.n176 0.155672
R1390 source.n219 source.n218 0.155672
R1391 source.n218 source.n180 0.155672
R1392 source.n210 source.n180 0.155672
R1393 source.n210 source.n209 0.155672
R1394 source.n209 source.n185 0.155672
R1395 source.n202 source.n185 0.155672
R1396 source.n202 source.n201 0.155672
R1397 source.n201 source.n189 0.155672
R1398 source.n194 source.n189 0.155672
R1399 plus.n3 plus.t0 2169.73
R1400 plus.n15 plus.t10 2169.73
R1401 plus.n20 plus.t12 2169.73
R1402 plus.n32 plus.t2 2169.73
R1403 plus.n1 plus.t11 2112.77
R1404 plus.n4 plus.t4 2112.77
R1405 plus.n6 plus.t8 2112.77
R1406 plus.n12 plus.t3 2112.77
R1407 plus.n14 plus.t6 2112.77
R1408 plus.n18 plus.t7 2112.77
R1409 plus.n21 plus.t5 2112.77
R1410 plus.n23 plus.t13 2112.77
R1411 plus.n29 plus.t1 2112.77
R1412 plus.n31 plus.t9 2112.77
R1413 plus.n3 plus.n2 161.489
R1414 plus.n20 plus.n19 161.489
R1415 plus.n5 plus.n2 161.3
R1416 plus.n8 plus.n7 161.3
R1417 plus.n9 plus.n1 161.3
R1418 plus.n11 plus.n10 161.3
R1419 plus.n13 plus.n0 161.3
R1420 plus.n16 plus.n15 161.3
R1421 plus.n22 plus.n19 161.3
R1422 plus.n25 plus.n24 161.3
R1423 plus.n26 plus.n18 161.3
R1424 plus.n28 plus.n27 161.3
R1425 plus.n30 plus.n17 161.3
R1426 plus.n33 plus.n32 161.3
R1427 plus.n7 plus.n1 73.0308
R1428 plus.n11 plus.n1 73.0308
R1429 plus.n28 plus.n18 73.0308
R1430 plus.n24 plus.n18 73.0308
R1431 plus.n6 plus.n5 54.0429
R1432 plus.n13 plus.n12 54.0429
R1433 plus.n30 plus.n29 54.0429
R1434 plus.n23 plus.n22 54.0429
R1435 plus.n5 plus.n4 37.9763
R1436 plus.n14 plus.n13 37.9763
R1437 plus.n31 plus.n30 37.9763
R1438 plus.n22 plus.n21 37.9763
R1439 plus.n4 plus.n3 35.055
R1440 plus.n15 plus.n14 35.055
R1441 plus.n32 plus.n31 35.055
R1442 plus.n21 plus.n20 35.055
R1443 plus plus.n33 34.4933
R1444 plus.n7 plus.n6 18.9884
R1445 plus.n12 plus.n11 18.9884
R1446 plus.n29 plus.n28 18.9884
R1447 plus.n24 plus.n23 18.9884
R1448 plus plus.n16 17.1047
R1449 plus.n8 plus.n2 0.189894
R1450 plus.n9 plus.n8 0.189894
R1451 plus.n10 plus.n9 0.189894
R1452 plus.n10 plus.n0 0.189894
R1453 plus.n16 plus.n0 0.189894
R1454 plus.n33 plus.n17 0.189894
R1455 plus.n27 plus.n17 0.189894
R1456 plus.n27 plus.n26 0.189894
R1457 plus.n26 plus.n25 0.189894
R1458 plus.n25 plus.n19 0.189894
R1459 drain_left.n134 drain_left.n0 289.615
R1460 drain_left.n279 drain_left.n145 289.615
R1461 drain_left.n44 drain_left.n43 185
R1462 drain_left.n49 drain_left.n48 185
R1463 drain_left.n51 drain_left.n50 185
R1464 drain_left.n40 drain_left.n39 185
R1465 drain_left.n57 drain_left.n56 185
R1466 drain_left.n59 drain_left.n58 185
R1467 drain_left.n36 drain_left.n35 185
R1468 drain_left.n66 drain_left.n65 185
R1469 drain_left.n67 drain_left.n34 185
R1470 drain_left.n69 drain_left.n68 185
R1471 drain_left.n32 drain_left.n31 185
R1472 drain_left.n75 drain_left.n74 185
R1473 drain_left.n77 drain_left.n76 185
R1474 drain_left.n28 drain_left.n27 185
R1475 drain_left.n83 drain_left.n82 185
R1476 drain_left.n85 drain_left.n84 185
R1477 drain_left.n24 drain_left.n23 185
R1478 drain_left.n91 drain_left.n90 185
R1479 drain_left.n93 drain_left.n92 185
R1480 drain_left.n20 drain_left.n19 185
R1481 drain_left.n99 drain_left.n98 185
R1482 drain_left.n101 drain_left.n100 185
R1483 drain_left.n16 drain_left.n15 185
R1484 drain_left.n107 drain_left.n106 185
R1485 drain_left.n110 drain_left.n109 185
R1486 drain_left.n108 drain_left.n12 185
R1487 drain_left.n115 drain_left.n11 185
R1488 drain_left.n117 drain_left.n116 185
R1489 drain_left.n119 drain_left.n118 185
R1490 drain_left.n8 drain_left.n7 185
R1491 drain_left.n125 drain_left.n124 185
R1492 drain_left.n127 drain_left.n126 185
R1493 drain_left.n4 drain_left.n3 185
R1494 drain_left.n133 drain_left.n132 185
R1495 drain_left.n135 drain_left.n134 185
R1496 drain_left.n280 drain_left.n279 185
R1497 drain_left.n278 drain_left.n277 185
R1498 drain_left.n149 drain_left.n148 185
R1499 drain_left.n272 drain_left.n271 185
R1500 drain_left.n270 drain_left.n269 185
R1501 drain_left.n153 drain_left.n152 185
R1502 drain_left.n264 drain_left.n263 185
R1503 drain_left.n262 drain_left.n261 185
R1504 drain_left.n260 drain_left.n156 185
R1505 drain_left.n160 drain_left.n157 185
R1506 drain_left.n255 drain_left.n254 185
R1507 drain_left.n253 drain_left.n252 185
R1508 drain_left.n162 drain_left.n161 185
R1509 drain_left.n247 drain_left.n246 185
R1510 drain_left.n245 drain_left.n244 185
R1511 drain_left.n166 drain_left.n165 185
R1512 drain_left.n239 drain_left.n238 185
R1513 drain_left.n237 drain_left.n236 185
R1514 drain_left.n170 drain_left.n169 185
R1515 drain_left.n231 drain_left.n230 185
R1516 drain_left.n229 drain_left.n228 185
R1517 drain_left.n174 drain_left.n173 185
R1518 drain_left.n223 drain_left.n222 185
R1519 drain_left.n221 drain_left.n220 185
R1520 drain_left.n178 drain_left.n177 185
R1521 drain_left.n215 drain_left.n214 185
R1522 drain_left.n213 drain_left.n180 185
R1523 drain_left.n212 drain_left.n211 185
R1524 drain_left.n183 drain_left.n181 185
R1525 drain_left.n206 drain_left.n205 185
R1526 drain_left.n204 drain_left.n203 185
R1527 drain_left.n187 drain_left.n186 185
R1528 drain_left.n198 drain_left.n197 185
R1529 drain_left.n196 drain_left.n195 185
R1530 drain_left.n191 drain_left.n190 185
R1531 drain_left.n45 drain_left.t11 149.524
R1532 drain_left.n192 drain_left.t13 149.524
R1533 drain_left.n49 drain_left.n43 104.615
R1534 drain_left.n50 drain_left.n49 104.615
R1535 drain_left.n50 drain_left.n39 104.615
R1536 drain_left.n57 drain_left.n39 104.615
R1537 drain_left.n58 drain_left.n57 104.615
R1538 drain_left.n58 drain_left.n35 104.615
R1539 drain_left.n66 drain_left.n35 104.615
R1540 drain_left.n67 drain_left.n66 104.615
R1541 drain_left.n68 drain_left.n67 104.615
R1542 drain_left.n68 drain_left.n31 104.615
R1543 drain_left.n75 drain_left.n31 104.615
R1544 drain_left.n76 drain_left.n75 104.615
R1545 drain_left.n76 drain_left.n27 104.615
R1546 drain_left.n83 drain_left.n27 104.615
R1547 drain_left.n84 drain_left.n83 104.615
R1548 drain_left.n84 drain_left.n23 104.615
R1549 drain_left.n91 drain_left.n23 104.615
R1550 drain_left.n92 drain_left.n91 104.615
R1551 drain_left.n92 drain_left.n19 104.615
R1552 drain_left.n99 drain_left.n19 104.615
R1553 drain_left.n100 drain_left.n99 104.615
R1554 drain_left.n100 drain_left.n15 104.615
R1555 drain_left.n107 drain_left.n15 104.615
R1556 drain_left.n109 drain_left.n107 104.615
R1557 drain_left.n109 drain_left.n108 104.615
R1558 drain_left.n108 drain_left.n11 104.615
R1559 drain_left.n117 drain_left.n11 104.615
R1560 drain_left.n118 drain_left.n117 104.615
R1561 drain_left.n118 drain_left.n7 104.615
R1562 drain_left.n125 drain_left.n7 104.615
R1563 drain_left.n126 drain_left.n125 104.615
R1564 drain_left.n126 drain_left.n3 104.615
R1565 drain_left.n133 drain_left.n3 104.615
R1566 drain_left.n134 drain_left.n133 104.615
R1567 drain_left.n279 drain_left.n278 104.615
R1568 drain_left.n278 drain_left.n148 104.615
R1569 drain_left.n271 drain_left.n148 104.615
R1570 drain_left.n271 drain_left.n270 104.615
R1571 drain_left.n270 drain_left.n152 104.615
R1572 drain_left.n263 drain_left.n152 104.615
R1573 drain_left.n263 drain_left.n262 104.615
R1574 drain_left.n262 drain_left.n156 104.615
R1575 drain_left.n160 drain_left.n156 104.615
R1576 drain_left.n254 drain_left.n160 104.615
R1577 drain_left.n254 drain_left.n253 104.615
R1578 drain_left.n253 drain_left.n161 104.615
R1579 drain_left.n246 drain_left.n161 104.615
R1580 drain_left.n246 drain_left.n245 104.615
R1581 drain_left.n245 drain_left.n165 104.615
R1582 drain_left.n238 drain_left.n165 104.615
R1583 drain_left.n238 drain_left.n237 104.615
R1584 drain_left.n237 drain_left.n169 104.615
R1585 drain_left.n230 drain_left.n169 104.615
R1586 drain_left.n230 drain_left.n229 104.615
R1587 drain_left.n229 drain_left.n173 104.615
R1588 drain_left.n222 drain_left.n173 104.615
R1589 drain_left.n222 drain_left.n221 104.615
R1590 drain_left.n221 drain_left.n177 104.615
R1591 drain_left.n214 drain_left.n177 104.615
R1592 drain_left.n214 drain_left.n213 104.615
R1593 drain_left.n213 drain_left.n212 104.615
R1594 drain_left.n212 drain_left.n181 104.615
R1595 drain_left.n205 drain_left.n181 104.615
R1596 drain_left.n205 drain_left.n204 104.615
R1597 drain_left.n204 drain_left.n186 104.615
R1598 drain_left.n197 drain_left.n186 104.615
R1599 drain_left.n197 drain_left.n196 104.615
R1600 drain_left.n196 drain_left.n190 104.615
R1601 drain_left.n143 drain_left.n141 59.2585
R1602 drain_left.n143 drain_left.n142 58.7154
R1603 drain_left.n140 drain_left.n139 58.7154
R1604 drain_left.n287 drain_left.n286 58.7154
R1605 drain_left.n285 drain_left.n284 58.7154
R1606 drain_left.n289 drain_left.n288 58.7153
R1607 drain_left.t11 drain_left.n43 52.3082
R1608 drain_left.t13 drain_left.n190 52.3082
R1609 drain_left.n140 drain_left.n138 47.8557
R1610 drain_left.n285 drain_left.n283 47.8557
R1611 drain_left drain_left.n144 40.3384
R1612 drain_left.n69 drain_left.n34 13.1884
R1613 drain_left.n116 drain_left.n115 13.1884
R1614 drain_left.n261 drain_left.n260 13.1884
R1615 drain_left.n215 drain_left.n180 13.1884
R1616 drain_left.n65 drain_left.n64 12.8005
R1617 drain_left.n70 drain_left.n32 12.8005
R1618 drain_left.n114 drain_left.n12 12.8005
R1619 drain_left.n119 drain_left.n10 12.8005
R1620 drain_left.n264 drain_left.n155 12.8005
R1621 drain_left.n259 drain_left.n157 12.8005
R1622 drain_left.n216 drain_left.n178 12.8005
R1623 drain_left.n211 drain_left.n182 12.8005
R1624 drain_left.n63 drain_left.n36 12.0247
R1625 drain_left.n74 drain_left.n73 12.0247
R1626 drain_left.n111 drain_left.n110 12.0247
R1627 drain_left.n120 drain_left.n8 12.0247
R1628 drain_left.n265 drain_left.n153 12.0247
R1629 drain_left.n256 drain_left.n255 12.0247
R1630 drain_left.n220 drain_left.n219 12.0247
R1631 drain_left.n210 drain_left.n183 12.0247
R1632 drain_left.n60 drain_left.n59 11.249
R1633 drain_left.n77 drain_left.n30 11.249
R1634 drain_left.n106 drain_left.n14 11.249
R1635 drain_left.n124 drain_left.n123 11.249
R1636 drain_left.n269 drain_left.n268 11.249
R1637 drain_left.n252 drain_left.n159 11.249
R1638 drain_left.n223 drain_left.n176 11.249
R1639 drain_left.n207 drain_left.n206 11.249
R1640 drain_left.n56 drain_left.n38 10.4732
R1641 drain_left.n78 drain_left.n28 10.4732
R1642 drain_left.n105 drain_left.n16 10.4732
R1643 drain_left.n127 drain_left.n6 10.4732
R1644 drain_left.n272 drain_left.n151 10.4732
R1645 drain_left.n251 drain_left.n162 10.4732
R1646 drain_left.n224 drain_left.n174 10.4732
R1647 drain_left.n203 drain_left.n185 10.4732
R1648 drain_left.n45 drain_left.n44 10.2747
R1649 drain_left.n192 drain_left.n191 10.2747
R1650 drain_left.n55 drain_left.n40 9.69747
R1651 drain_left.n82 drain_left.n81 9.69747
R1652 drain_left.n102 drain_left.n101 9.69747
R1653 drain_left.n128 drain_left.n4 9.69747
R1654 drain_left.n273 drain_left.n149 9.69747
R1655 drain_left.n248 drain_left.n247 9.69747
R1656 drain_left.n228 drain_left.n227 9.69747
R1657 drain_left.n202 drain_left.n187 9.69747
R1658 drain_left.n138 drain_left.n137 9.45567
R1659 drain_left.n283 drain_left.n282 9.45567
R1660 drain_left.n2 drain_left.n1 9.3005
R1661 drain_left.n131 drain_left.n130 9.3005
R1662 drain_left.n129 drain_left.n128 9.3005
R1663 drain_left.n6 drain_left.n5 9.3005
R1664 drain_left.n123 drain_left.n122 9.3005
R1665 drain_left.n121 drain_left.n120 9.3005
R1666 drain_left.n10 drain_left.n9 9.3005
R1667 drain_left.n89 drain_left.n88 9.3005
R1668 drain_left.n87 drain_left.n86 9.3005
R1669 drain_left.n26 drain_left.n25 9.3005
R1670 drain_left.n81 drain_left.n80 9.3005
R1671 drain_left.n79 drain_left.n78 9.3005
R1672 drain_left.n30 drain_left.n29 9.3005
R1673 drain_left.n73 drain_left.n72 9.3005
R1674 drain_left.n71 drain_left.n70 9.3005
R1675 drain_left.n47 drain_left.n46 9.3005
R1676 drain_left.n42 drain_left.n41 9.3005
R1677 drain_left.n53 drain_left.n52 9.3005
R1678 drain_left.n55 drain_left.n54 9.3005
R1679 drain_left.n38 drain_left.n37 9.3005
R1680 drain_left.n61 drain_left.n60 9.3005
R1681 drain_left.n63 drain_left.n62 9.3005
R1682 drain_left.n64 drain_left.n33 9.3005
R1683 drain_left.n22 drain_left.n21 9.3005
R1684 drain_left.n95 drain_left.n94 9.3005
R1685 drain_left.n97 drain_left.n96 9.3005
R1686 drain_left.n18 drain_left.n17 9.3005
R1687 drain_left.n103 drain_left.n102 9.3005
R1688 drain_left.n105 drain_left.n104 9.3005
R1689 drain_left.n14 drain_left.n13 9.3005
R1690 drain_left.n112 drain_left.n111 9.3005
R1691 drain_left.n114 drain_left.n113 9.3005
R1692 drain_left.n137 drain_left.n136 9.3005
R1693 drain_left.n194 drain_left.n193 9.3005
R1694 drain_left.n189 drain_left.n188 9.3005
R1695 drain_left.n200 drain_left.n199 9.3005
R1696 drain_left.n202 drain_left.n201 9.3005
R1697 drain_left.n185 drain_left.n184 9.3005
R1698 drain_left.n208 drain_left.n207 9.3005
R1699 drain_left.n210 drain_left.n209 9.3005
R1700 drain_left.n182 drain_left.n179 9.3005
R1701 drain_left.n241 drain_left.n240 9.3005
R1702 drain_left.n243 drain_left.n242 9.3005
R1703 drain_left.n164 drain_left.n163 9.3005
R1704 drain_left.n249 drain_left.n248 9.3005
R1705 drain_left.n251 drain_left.n250 9.3005
R1706 drain_left.n159 drain_left.n158 9.3005
R1707 drain_left.n257 drain_left.n256 9.3005
R1708 drain_left.n259 drain_left.n258 9.3005
R1709 drain_left.n282 drain_left.n281 9.3005
R1710 drain_left.n147 drain_left.n146 9.3005
R1711 drain_left.n276 drain_left.n275 9.3005
R1712 drain_left.n274 drain_left.n273 9.3005
R1713 drain_left.n151 drain_left.n150 9.3005
R1714 drain_left.n268 drain_left.n267 9.3005
R1715 drain_left.n266 drain_left.n265 9.3005
R1716 drain_left.n155 drain_left.n154 9.3005
R1717 drain_left.n168 drain_left.n167 9.3005
R1718 drain_left.n235 drain_left.n234 9.3005
R1719 drain_left.n233 drain_left.n232 9.3005
R1720 drain_left.n172 drain_left.n171 9.3005
R1721 drain_left.n227 drain_left.n226 9.3005
R1722 drain_left.n225 drain_left.n224 9.3005
R1723 drain_left.n176 drain_left.n175 9.3005
R1724 drain_left.n219 drain_left.n218 9.3005
R1725 drain_left.n217 drain_left.n216 9.3005
R1726 drain_left.n52 drain_left.n51 8.92171
R1727 drain_left.n85 drain_left.n26 8.92171
R1728 drain_left.n98 drain_left.n18 8.92171
R1729 drain_left.n132 drain_left.n131 8.92171
R1730 drain_left.n277 drain_left.n276 8.92171
R1731 drain_left.n244 drain_left.n164 8.92171
R1732 drain_left.n231 drain_left.n172 8.92171
R1733 drain_left.n199 drain_left.n198 8.92171
R1734 drain_left.n48 drain_left.n42 8.14595
R1735 drain_left.n86 drain_left.n24 8.14595
R1736 drain_left.n97 drain_left.n20 8.14595
R1737 drain_left.n135 drain_left.n2 8.14595
R1738 drain_left.n280 drain_left.n147 8.14595
R1739 drain_left.n243 drain_left.n166 8.14595
R1740 drain_left.n232 drain_left.n170 8.14595
R1741 drain_left.n195 drain_left.n189 8.14595
R1742 drain_left.n47 drain_left.n44 7.3702
R1743 drain_left.n90 drain_left.n89 7.3702
R1744 drain_left.n94 drain_left.n93 7.3702
R1745 drain_left.n136 drain_left.n0 7.3702
R1746 drain_left.n281 drain_left.n145 7.3702
R1747 drain_left.n240 drain_left.n239 7.3702
R1748 drain_left.n236 drain_left.n235 7.3702
R1749 drain_left.n194 drain_left.n191 7.3702
R1750 drain_left.n90 drain_left.n22 6.59444
R1751 drain_left.n93 drain_left.n22 6.59444
R1752 drain_left.n138 drain_left.n0 6.59444
R1753 drain_left.n283 drain_left.n145 6.59444
R1754 drain_left.n239 drain_left.n168 6.59444
R1755 drain_left.n236 drain_left.n168 6.59444
R1756 drain_left drain_left.n289 6.19632
R1757 drain_left.n48 drain_left.n47 5.81868
R1758 drain_left.n89 drain_left.n24 5.81868
R1759 drain_left.n94 drain_left.n20 5.81868
R1760 drain_left.n136 drain_left.n135 5.81868
R1761 drain_left.n281 drain_left.n280 5.81868
R1762 drain_left.n240 drain_left.n166 5.81868
R1763 drain_left.n235 drain_left.n170 5.81868
R1764 drain_left.n195 drain_left.n194 5.81868
R1765 drain_left.n51 drain_left.n42 5.04292
R1766 drain_left.n86 drain_left.n85 5.04292
R1767 drain_left.n98 drain_left.n97 5.04292
R1768 drain_left.n132 drain_left.n2 5.04292
R1769 drain_left.n277 drain_left.n147 5.04292
R1770 drain_left.n244 drain_left.n243 5.04292
R1771 drain_left.n232 drain_left.n231 5.04292
R1772 drain_left.n198 drain_left.n189 5.04292
R1773 drain_left.n52 drain_left.n40 4.26717
R1774 drain_left.n82 drain_left.n26 4.26717
R1775 drain_left.n101 drain_left.n18 4.26717
R1776 drain_left.n131 drain_left.n4 4.26717
R1777 drain_left.n276 drain_left.n149 4.26717
R1778 drain_left.n247 drain_left.n164 4.26717
R1779 drain_left.n228 drain_left.n172 4.26717
R1780 drain_left.n199 drain_left.n187 4.26717
R1781 drain_left.n56 drain_left.n55 3.49141
R1782 drain_left.n81 drain_left.n28 3.49141
R1783 drain_left.n102 drain_left.n16 3.49141
R1784 drain_left.n128 drain_left.n127 3.49141
R1785 drain_left.n273 drain_left.n272 3.49141
R1786 drain_left.n248 drain_left.n162 3.49141
R1787 drain_left.n227 drain_left.n174 3.49141
R1788 drain_left.n203 drain_left.n202 3.49141
R1789 drain_left.n193 drain_left.n192 2.84303
R1790 drain_left.n46 drain_left.n45 2.84303
R1791 drain_left.n59 drain_left.n38 2.71565
R1792 drain_left.n78 drain_left.n77 2.71565
R1793 drain_left.n106 drain_left.n105 2.71565
R1794 drain_left.n124 drain_left.n6 2.71565
R1795 drain_left.n269 drain_left.n151 2.71565
R1796 drain_left.n252 drain_left.n251 2.71565
R1797 drain_left.n224 drain_left.n223 2.71565
R1798 drain_left.n206 drain_left.n185 2.71565
R1799 drain_left.n60 drain_left.n36 1.93989
R1800 drain_left.n74 drain_left.n30 1.93989
R1801 drain_left.n110 drain_left.n14 1.93989
R1802 drain_left.n123 drain_left.n8 1.93989
R1803 drain_left.n268 drain_left.n153 1.93989
R1804 drain_left.n255 drain_left.n159 1.93989
R1805 drain_left.n220 drain_left.n176 1.93989
R1806 drain_left.n207 drain_left.n183 1.93989
R1807 drain_left.n65 drain_left.n63 1.16414
R1808 drain_left.n73 drain_left.n32 1.16414
R1809 drain_left.n111 drain_left.n12 1.16414
R1810 drain_left.n120 drain_left.n119 1.16414
R1811 drain_left.n265 drain_left.n264 1.16414
R1812 drain_left.n256 drain_left.n157 1.16414
R1813 drain_left.n219 drain_left.n178 1.16414
R1814 drain_left.n211 drain_left.n210 1.16414
R1815 drain_left.n141 drain_left.t8 0.7925
R1816 drain_left.n141 drain_left.t1 0.7925
R1817 drain_left.n142 drain_left.t6 0.7925
R1818 drain_left.n142 drain_left.t0 0.7925
R1819 drain_left.n139 drain_left.t4 0.7925
R1820 drain_left.n139 drain_left.t12 0.7925
R1821 drain_left.n288 drain_left.t7 0.7925
R1822 drain_left.n288 drain_left.t3 0.7925
R1823 drain_left.n286 drain_left.t2 0.7925
R1824 drain_left.n286 drain_left.t10 0.7925
R1825 drain_left.n284 drain_left.t9 0.7925
R1826 drain_left.n284 drain_left.t5 0.7925
R1827 drain_left.n287 drain_left.n285 0.543603
R1828 drain_left.n289 drain_left.n287 0.543603
R1829 drain_left.n64 drain_left.n34 0.388379
R1830 drain_left.n70 drain_left.n69 0.388379
R1831 drain_left.n115 drain_left.n114 0.388379
R1832 drain_left.n116 drain_left.n10 0.388379
R1833 drain_left.n261 drain_left.n155 0.388379
R1834 drain_left.n260 drain_left.n259 0.388379
R1835 drain_left.n216 drain_left.n215 0.388379
R1836 drain_left.n182 drain_left.n180 0.388379
R1837 drain_left.n144 drain_left.n140 0.352482
R1838 drain_left.n46 drain_left.n41 0.155672
R1839 drain_left.n53 drain_left.n41 0.155672
R1840 drain_left.n54 drain_left.n53 0.155672
R1841 drain_left.n54 drain_left.n37 0.155672
R1842 drain_left.n61 drain_left.n37 0.155672
R1843 drain_left.n62 drain_left.n61 0.155672
R1844 drain_left.n62 drain_left.n33 0.155672
R1845 drain_left.n71 drain_left.n33 0.155672
R1846 drain_left.n72 drain_left.n71 0.155672
R1847 drain_left.n72 drain_left.n29 0.155672
R1848 drain_left.n79 drain_left.n29 0.155672
R1849 drain_left.n80 drain_left.n79 0.155672
R1850 drain_left.n80 drain_left.n25 0.155672
R1851 drain_left.n87 drain_left.n25 0.155672
R1852 drain_left.n88 drain_left.n87 0.155672
R1853 drain_left.n88 drain_left.n21 0.155672
R1854 drain_left.n95 drain_left.n21 0.155672
R1855 drain_left.n96 drain_left.n95 0.155672
R1856 drain_left.n96 drain_left.n17 0.155672
R1857 drain_left.n103 drain_left.n17 0.155672
R1858 drain_left.n104 drain_left.n103 0.155672
R1859 drain_left.n104 drain_left.n13 0.155672
R1860 drain_left.n112 drain_left.n13 0.155672
R1861 drain_left.n113 drain_left.n112 0.155672
R1862 drain_left.n113 drain_left.n9 0.155672
R1863 drain_left.n121 drain_left.n9 0.155672
R1864 drain_left.n122 drain_left.n121 0.155672
R1865 drain_left.n122 drain_left.n5 0.155672
R1866 drain_left.n129 drain_left.n5 0.155672
R1867 drain_left.n130 drain_left.n129 0.155672
R1868 drain_left.n130 drain_left.n1 0.155672
R1869 drain_left.n137 drain_left.n1 0.155672
R1870 drain_left.n282 drain_left.n146 0.155672
R1871 drain_left.n275 drain_left.n146 0.155672
R1872 drain_left.n275 drain_left.n274 0.155672
R1873 drain_left.n274 drain_left.n150 0.155672
R1874 drain_left.n267 drain_left.n150 0.155672
R1875 drain_left.n267 drain_left.n266 0.155672
R1876 drain_left.n266 drain_left.n154 0.155672
R1877 drain_left.n258 drain_left.n154 0.155672
R1878 drain_left.n258 drain_left.n257 0.155672
R1879 drain_left.n257 drain_left.n158 0.155672
R1880 drain_left.n250 drain_left.n158 0.155672
R1881 drain_left.n250 drain_left.n249 0.155672
R1882 drain_left.n249 drain_left.n163 0.155672
R1883 drain_left.n242 drain_left.n163 0.155672
R1884 drain_left.n242 drain_left.n241 0.155672
R1885 drain_left.n241 drain_left.n167 0.155672
R1886 drain_left.n234 drain_left.n167 0.155672
R1887 drain_left.n234 drain_left.n233 0.155672
R1888 drain_left.n233 drain_left.n171 0.155672
R1889 drain_left.n226 drain_left.n171 0.155672
R1890 drain_left.n226 drain_left.n225 0.155672
R1891 drain_left.n225 drain_left.n175 0.155672
R1892 drain_left.n218 drain_left.n175 0.155672
R1893 drain_left.n218 drain_left.n217 0.155672
R1894 drain_left.n217 drain_left.n179 0.155672
R1895 drain_left.n209 drain_left.n179 0.155672
R1896 drain_left.n209 drain_left.n208 0.155672
R1897 drain_left.n208 drain_left.n184 0.155672
R1898 drain_left.n201 drain_left.n184 0.155672
R1899 drain_left.n201 drain_left.n200 0.155672
R1900 drain_left.n200 drain_left.n188 0.155672
R1901 drain_left.n193 drain_left.n188 0.155672
R1902 drain_left.n144 drain_left.n143 0.0809298
C0 plus minus 7.70658f
C1 minus source 9.57778f
C2 drain_right drain_left 0.889001f
C3 plus source 9.59318f
C4 minus drain_right 10.4678f
C5 minus drain_left 0.171678f
C6 plus drain_right 0.325724f
C7 source drain_right 55.4743f
C8 plus drain_left 10.6286f
C9 source drain_left 55.4954f
C10 drain_right a_n1724_n5888# 11.24571f
C11 drain_left a_n1724_n5888# 11.519239f
C12 source a_n1724_n5888# 10.681088f
C13 minus a_n1724_n5888# 7.58053f
C14 plus a_n1724_n5888# 10.41975f
C15 drain_left.n0 a_n1724_n5888# 0.042815f
C16 drain_left.n1 a_n1724_n5888# 0.031057f
C17 drain_left.n2 a_n1724_n5888# 0.016689f
C18 drain_left.n3 a_n1724_n5888# 0.039446f
C19 drain_left.n4 a_n1724_n5888# 0.01767f
C20 drain_left.n5 a_n1724_n5888# 0.031057f
C21 drain_left.n6 a_n1724_n5888# 0.016689f
C22 drain_left.n7 a_n1724_n5888# 0.039446f
C23 drain_left.n8 a_n1724_n5888# 0.01767f
C24 drain_left.n9 a_n1724_n5888# 0.031057f
C25 drain_left.n10 a_n1724_n5888# 0.016689f
C26 drain_left.n11 a_n1724_n5888# 0.039446f
C27 drain_left.n12 a_n1724_n5888# 0.01767f
C28 drain_left.n13 a_n1724_n5888# 0.031057f
C29 drain_left.n14 a_n1724_n5888# 0.016689f
C30 drain_left.n15 a_n1724_n5888# 0.039446f
C31 drain_left.n16 a_n1724_n5888# 0.01767f
C32 drain_left.n17 a_n1724_n5888# 0.031057f
C33 drain_left.n18 a_n1724_n5888# 0.016689f
C34 drain_left.n19 a_n1724_n5888# 0.039446f
C35 drain_left.n20 a_n1724_n5888# 0.01767f
C36 drain_left.n21 a_n1724_n5888# 0.031057f
C37 drain_left.n22 a_n1724_n5888# 0.016689f
C38 drain_left.n23 a_n1724_n5888# 0.039446f
C39 drain_left.n24 a_n1724_n5888# 0.01767f
C40 drain_left.n25 a_n1724_n5888# 0.031057f
C41 drain_left.n26 a_n1724_n5888# 0.016689f
C42 drain_left.n27 a_n1724_n5888# 0.039446f
C43 drain_left.n28 a_n1724_n5888# 0.01767f
C44 drain_left.n29 a_n1724_n5888# 0.031057f
C45 drain_left.n30 a_n1724_n5888# 0.016689f
C46 drain_left.n31 a_n1724_n5888# 0.039446f
C47 drain_left.n32 a_n1724_n5888# 0.01767f
C48 drain_left.n33 a_n1724_n5888# 0.031057f
C49 drain_left.n34 a_n1724_n5888# 0.017179f
C50 drain_left.n35 a_n1724_n5888# 0.039446f
C51 drain_left.n36 a_n1724_n5888# 0.01767f
C52 drain_left.n37 a_n1724_n5888# 0.031057f
C53 drain_left.n38 a_n1724_n5888# 0.016689f
C54 drain_left.n39 a_n1724_n5888# 0.039446f
C55 drain_left.n40 a_n1724_n5888# 0.01767f
C56 drain_left.n41 a_n1724_n5888# 0.031057f
C57 drain_left.n42 a_n1724_n5888# 0.016689f
C58 drain_left.n43 a_n1724_n5888# 0.029584f
C59 drain_left.n44 a_n1724_n5888# 0.027885f
C60 drain_left.t11 a_n1724_n5888# 0.068796f
C61 drain_left.n45 a_n1724_n5888# 0.37892f
C62 drain_left.n46 a_n1724_n5888# 3.36254f
C63 drain_left.n47 a_n1724_n5888# 0.016689f
C64 drain_left.n48 a_n1724_n5888# 0.01767f
C65 drain_left.n49 a_n1724_n5888# 0.039446f
C66 drain_left.n50 a_n1724_n5888# 0.039446f
C67 drain_left.n51 a_n1724_n5888# 0.01767f
C68 drain_left.n52 a_n1724_n5888# 0.016689f
C69 drain_left.n53 a_n1724_n5888# 0.031057f
C70 drain_left.n54 a_n1724_n5888# 0.031057f
C71 drain_left.n55 a_n1724_n5888# 0.016689f
C72 drain_left.n56 a_n1724_n5888# 0.01767f
C73 drain_left.n57 a_n1724_n5888# 0.039446f
C74 drain_left.n58 a_n1724_n5888# 0.039446f
C75 drain_left.n59 a_n1724_n5888# 0.01767f
C76 drain_left.n60 a_n1724_n5888# 0.016689f
C77 drain_left.n61 a_n1724_n5888# 0.031057f
C78 drain_left.n62 a_n1724_n5888# 0.031057f
C79 drain_left.n63 a_n1724_n5888# 0.016689f
C80 drain_left.n64 a_n1724_n5888# 0.016689f
C81 drain_left.n65 a_n1724_n5888# 0.01767f
C82 drain_left.n66 a_n1724_n5888# 0.039446f
C83 drain_left.n67 a_n1724_n5888# 0.039446f
C84 drain_left.n68 a_n1724_n5888# 0.039446f
C85 drain_left.n69 a_n1724_n5888# 0.017179f
C86 drain_left.n70 a_n1724_n5888# 0.016689f
C87 drain_left.n71 a_n1724_n5888# 0.031057f
C88 drain_left.n72 a_n1724_n5888# 0.031057f
C89 drain_left.n73 a_n1724_n5888# 0.016689f
C90 drain_left.n74 a_n1724_n5888# 0.01767f
C91 drain_left.n75 a_n1724_n5888# 0.039446f
C92 drain_left.n76 a_n1724_n5888# 0.039446f
C93 drain_left.n77 a_n1724_n5888# 0.01767f
C94 drain_left.n78 a_n1724_n5888# 0.016689f
C95 drain_left.n79 a_n1724_n5888# 0.031057f
C96 drain_left.n80 a_n1724_n5888# 0.031057f
C97 drain_left.n81 a_n1724_n5888# 0.016689f
C98 drain_left.n82 a_n1724_n5888# 0.01767f
C99 drain_left.n83 a_n1724_n5888# 0.039446f
C100 drain_left.n84 a_n1724_n5888# 0.039446f
C101 drain_left.n85 a_n1724_n5888# 0.01767f
C102 drain_left.n86 a_n1724_n5888# 0.016689f
C103 drain_left.n87 a_n1724_n5888# 0.031057f
C104 drain_left.n88 a_n1724_n5888# 0.031057f
C105 drain_left.n89 a_n1724_n5888# 0.016689f
C106 drain_left.n90 a_n1724_n5888# 0.01767f
C107 drain_left.n91 a_n1724_n5888# 0.039446f
C108 drain_left.n92 a_n1724_n5888# 0.039446f
C109 drain_left.n93 a_n1724_n5888# 0.01767f
C110 drain_left.n94 a_n1724_n5888# 0.016689f
C111 drain_left.n95 a_n1724_n5888# 0.031057f
C112 drain_left.n96 a_n1724_n5888# 0.031057f
C113 drain_left.n97 a_n1724_n5888# 0.016689f
C114 drain_left.n98 a_n1724_n5888# 0.01767f
C115 drain_left.n99 a_n1724_n5888# 0.039446f
C116 drain_left.n100 a_n1724_n5888# 0.039446f
C117 drain_left.n101 a_n1724_n5888# 0.01767f
C118 drain_left.n102 a_n1724_n5888# 0.016689f
C119 drain_left.n103 a_n1724_n5888# 0.031057f
C120 drain_left.n104 a_n1724_n5888# 0.031057f
C121 drain_left.n105 a_n1724_n5888# 0.016689f
C122 drain_left.n106 a_n1724_n5888# 0.01767f
C123 drain_left.n107 a_n1724_n5888# 0.039446f
C124 drain_left.n108 a_n1724_n5888# 0.039446f
C125 drain_left.n109 a_n1724_n5888# 0.039446f
C126 drain_left.n110 a_n1724_n5888# 0.01767f
C127 drain_left.n111 a_n1724_n5888# 0.016689f
C128 drain_left.n112 a_n1724_n5888# 0.031057f
C129 drain_left.n113 a_n1724_n5888# 0.031057f
C130 drain_left.n114 a_n1724_n5888# 0.016689f
C131 drain_left.n115 a_n1724_n5888# 0.017179f
C132 drain_left.n116 a_n1724_n5888# 0.017179f
C133 drain_left.n117 a_n1724_n5888# 0.039446f
C134 drain_left.n118 a_n1724_n5888# 0.039446f
C135 drain_left.n119 a_n1724_n5888# 0.01767f
C136 drain_left.n120 a_n1724_n5888# 0.016689f
C137 drain_left.n121 a_n1724_n5888# 0.031057f
C138 drain_left.n122 a_n1724_n5888# 0.031057f
C139 drain_left.n123 a_n1724_n5888# 0.016689f
C140 drain_left.n124 a_n1724_n5888# 0.01767f
C141 drain_left.n125 a_n1724_n5888# 0.039446f
C142 drain_left.n126 a_n1724_n5888# 0.039446f
C143 drain_left.n127 a_n1724_n5888# 0.01767f
C144 drain_left.n128 a_n1724_n5888# 0.016689f
C145 drain_left.n129 a_n1724_n5888# 0.031057f
C146 drain_left.n130 a_n1724_n5888# 0.031057f
C147 drain_left.n131 a_n1724_n5888# 0.016689f
C148 drain_left.n132 a_n1724_n5888# 0.01767f
C149 drain_left.n133 a_n1724_n5888# 0.039446f
C150 drain_left.n134 a_n1724_n5888# 0.083911f
C151 drain_left.n135 a_n1724_n5888# 0.01767f
C152 drain_left.n136 a_n1724_n5888# 0.016689f
C153 drain_left.n137 a_n1724_n5888# 0.068392f
C154 drain_left.n138 a_n1724_n5888# 0.069439f
C155 drain_left.t4 a_n1724_n5888# 0.613552f
C156 drain_left.t12 a_n1724_n5888# 0.613552f
C157 drain_left.n139 a_n1724_n5888# 5.65454f
C158 drain_left.n140 a_n1724_n5888# 0.465076f
C159 drain_left.t8 a_n1724_n5888# 0.613552f
C160 drain_left.t1 a_n1724_n5888# 0.613552f
C161 drain_left.n141 a_n1724_n5888# 5.65806f
C162 drain_left.t6 a_n1724_n5888# 0.613552f
C163 drain_left.t0 a_n1724_n5888# 0.613552f
C164 drain_left.n142 a_n1724_n5888# 5.65454f
C165 drain_left.n143 a_n1724_n5888# 0.714083f
C166 drain_left.n144 a_n1724_n5888# 2.49578f
C167 drain_left.n145 a_n1724_n5888# 0.042815f
C168 drain_left.n146 a_n1724_n5888# 0.031057f
C169 drain_left.n147 a_n1724_n5888# 0.016689f
C170 drain_left.n148 a_n1724_n5888# 0.039446f
C171 drain_left.n149 a_n1724_n5888# 0.01767f
C172 drain_left.n150 a_n1724_n5888# 0.031057f
C173 drain_left.n151 a_n1724_n5888# 0.016689f
C174 drain_left.n152 a_n1724_n5888# 0.039446f
C175 drain_left.n153 a_n1724_n5888# 0.01767f
C176 drain_left.n154 a_n1724_n5888# 0.031057f
C177 drain_left.n155 a_n1724_n5888# 0.016689f
C178 drain_left.n156 a_n1724_n5888# 0.039446f
C179 drain_left.n157 a_n1724_n5888# 0.01767f
C180 drain_left.n158 a_n1724_n5888# 0.031057f
C181 drain_left.n159 a_n1724_n5888# 0.016689f
C182 drain_left.n160 a_n1724_n5888# 0.039446f
C183 drain_left.n161 a_n1724_n5888# 0.039446f
C184 drain_left.n162 a_n1724_n5888# 0.01767f
C185 drain_left.n163 a_n1724_n5888# 0.031057f
C186 drain_left.n164 a_n1724_n5888# 0.016689f
C187 drain_left.n165 a_n1724_n5888# 0.039446f
C188 drain_left.n166 a_n1724_n5888# 0.01767f
C189 drain_left.n167 a_n1724_n5888# 0.031057f
C190 drain_left.n168 a_n1724_n5888# 0.016689f
C191 drain_left.n169 a_n1724_n5888# 0.039446f
C192 drain_left.n170 a_n1724_n5888# 0.01767f
C193 drain_left.n171 a_n1724_n5888# 0.031057f
C194 drain_left.n172 a_n1724_n5888# 0.016689f
C195 drain_left.n173 a_n1724_n5888# 0.039446f
C196 drain_left.n174 a_n1724_n5888# 0.01767f
C197 drain_left.n175 a_n1724_n5888# 0.031057f
C198 drain_left.n176 a_n1724_n5888# 0.016689f
C199 drain_left.n177 a_n1724_n5888# 0.039446f
C200 drain_left.n178 a_n1724_n5888# 0.01767f
C201 drain_left.n179 a_n1724_n5888# 0.031057f
C202 drain_left.n180 a_n1724_n5888# 0.017179f
C203 drain_left.n181 a_n1724_n5888# 0.039446f
C204 drain_left.n182 a_n1724_n5888# 0.016689f
C205 drain_left.n183 a_n1724_n5888# 0.01767f
C206 drain_left.n184 a_n1724_n5888# 0.031057f
C207 drain_left.n185 a_n1724_n5888# 0.016689f
C208 drain_left.n186 a_n1724_n5888# 0.039446f
C209 drain_left.n187 a_n1724_n5888# 0.01767f
C210 drain_left.n188 a_n1724_n5888# 0.031057f
C211 drain_left.n189 a_n1724_n5888# 0.016689f
C212 drain_left.n190 a_n1724_n5888# 0.029584f
C213 drain_left.n191 a_n1724_n5888# 0.027885f
C214 drain_left.t13 a_n1724_n5888# 0.068796f
C215 drain_left.n192 a_n1724_n5888# 0.37892f
C216 drain_left.n193 a_n1724_n5888# 3.36254f
C217 drain_left.n194 a_n1724_n5888# 0.016689f
C218 drain_left.n195 a_n1724_n5888# 0.01767f
C219 drain_left.n196 a_n1724_n5888# 0.039446f
C220 drain_left.n197 a_n1724_n5888# 0.039446f
C221 drain_left.n198 a_n1724_n5888# 0.01767f
C222 drain_left.n199 a_n1724_n5888# 0.016689f
C223 drain_left.n200 a_n1724_n5888# 0.031057f
C224 drain_left.n201 a_n1724_n5888# 0.031057f
C225 drain_left.n202 a_n1724_n5888# 0.016689f
C226 drain_left.n203 a_n1724_n5888# 0.01767f
C227 drain_left.n204 a_n1724_n5888# 0.039446f
C228 drain_left.n205 a_n1724_n5888# 0.039446f
C229 drain_left.n206 a_n1724_n5888# 0.01767f
C230 drain_left.n207 a_n1724_n5888# 0.016689f
C231 drain_left.n208 a_n1724_n5888# 0.031057f
C232 drain_left.n209 a_n1724_n5888# 0.031057f
C233 drain_left.n210 a_n1724_n5888# 0.016689f
C234 drain_left.n211 a_n1724_n5888# 0.01767f
C235 drain_left.n212 a_n1724_n5888# 0.039446f
C236 drain_left.n213 a_n1724_n5888# 0.039446f
C237 drain_left.n214 a_n1724_n5888# 0.039446f
C238 drain_left.n215 a_n1724_n5888# 0.017179f
C239 drain_left.n216 a_n1724_n5888# 0.016689f
C240 drain_left.n217 a_n1724_n5888# 0.031057f
C241 drain_left.n218 a_n1724_n5888# 0.031057f
C242 drain_left.n219 a_n1724_n5888# 0.016689f
C243 drain_left.n220 a_n1724_n5888# 0.01767f
C244 drain_left.n221 a_n1724_n5888# 0.039446f
C245 drain_left.n222 a_n1724_n5888# 0.039446f
C246 drain_left.n223 a_n1724_n5888# 0.01767f
C247 drain_left.n224 a_n1724_n5888# 0.016689f
C248 drain_left.n225 a_n1724_n5888# 0.031057f
C249 drain_left.n226 a_n1724_n5888# 0.031057f
C250 drain_left.n227 a_n1724_n5888# 0.016689f
C251 drain_left.n228 a_n1724_n5888# 0.01767f
C252 drain_left.n229 a_n1724_n5888# 0.039446f
C253 drain_left.n230 a_n1724_n5888# 0.039446f
C254 drain_left.n231 a_n1724_n5888# 0.01767f
C255 drain_left.n232 a_n1724_n5888# 0.016689f
C256 drain_left.n233 a_n1724_n5888# 0.031057f
C257 drain_left.n234 a_n1724_n5888# 0.031057f
C258 drain_left.n235 a_n1724_n5888# 0.016689f
C259 drain_left.n236 a_n1724_n5888# 0.01767f
C260 drain_left.n237 a_n1724_n5888# 0.039446f
C261 drain_left.n238 a_n1724_n5888# 0.039446f
C262 drain_left.n239 a_n1724_n5888# 0.01767f
C263 drain_left.n240 a_n1724_n5888# 0.016689f
C264 drain_left.n241 a_n1724_n5888# 0.031057f
C265 drain_left.n242 a_n1724_n5888# 0.031057f
C266 drain_left.n243 a_n1724_n5888# 0.016689f
C267 drain_left.n244 a_n1724_n5888# 0.01767f
C268 drain_left.n245 a_n1724_n5888# 0.039446f
C269 drain_left.n246 a_n1724_n5888# 0.039446f
C270 drain_left.n247 a_n1724_n5888# 0.01767f
C271 drain_left.n248 a_n1724_n5888# 0.016689f
C272 drain_left.n249 a_n1724_n5888# 0.031057f
C273 drain_left.n250 a_n1724_n5888# 0.031057f
C274 drain_left.n251 a_n1724_n5888# 0.016689f
C275 drain_left.n252 a_n1724_n5888# 0.01767f
C276 drain_left.n253 a_n1724_n5888# 0.039446f
C277 drain_left.n254 a_n1724_n5888# 0.039446f
C278 drain_left.n255 a_n1724_n5888# 0.01767f
C279 drain_left.n256 a_n1724_n5888# 0.016689f
C280 drain_left.n257 a_n1724_n5888# 0.031057f
C281 drain_left.n258 a_n1724_n5888# 0.031057f
C282 drain_left.n259 a_n1724_n5888# 0.016689f
C283 drain_left.n260 a_n1724_n5888# 0.017179f
C284 drain_left.n261 a_n1724_n5888# 0.017179f
C285 drain_left.n262 a_n1724_n5888# 0.039446f
C286 drain_left.n263 a_n1724_n5888# 0.039446f
C287 drain_left.n264 a_n1724_n5888# 0.01767f
C288 drain_left.n265 a_n1724_n5888# 0.016689f
C289 drain_left.n266 a_n1724_n5888# 0.031057f
C290 drain_left.n267 a_n1724_n5888# 0.031057f
C291 drain_left.n268 a_n1724_n5888# 0.016689f
C292 drain_left.n269 a_n1724_n5888# 0.01767f
C293 drain_left.n270 a_n1724_n5888# 0.039446f
C294 drain_left.n271 a_n1724_n5888# 0.039446f
C295 drain_left.n272 a_n1724_n5888# 0.01767f
C296 drain_left.n273 a_n1724_n5888# 0.016689f
C297 drain_left.n274 a_n1724_n5888# 0.031057f
C298 drain_left.n275 a_n1724_n5888# 0.031057f
C299 drain_left.n276 a_n1724_n5888# 0.016689f
C300 drain_left.n277 a_n1724_n5888# 0.01767f
C301 drain_left.n278 a_n1724_n5888# 0.039446f
C302 drain_left.n279 a_n1724_n5888# 0.083911f
C303 drain_left.n280 a_n1724_n5888# 0.01767f
C304 drain_left.n281 a_n1724_n5888# 0.016689f
C305 drain_left.n282 a_n1724_n5888# 0.068392f
C306 drain_left.n283 a_n1724_n5888# 0.069439f
C307 drain_left.t9 a_n1724_n5888# 0.613552f
C308 drain_left.t5 a_n1724_n5888# 0.613552f
C309 drain_left.n284 a_n1724_n5888# 5.65454f
C310 drain_left.n285 a_n1724_n5888# 0.482154f
C311 drain_left.t2 a_n1724_n5888# 0.613552f
C312 drain_left.t10 a_n1724_n5888# 0.613552f
C313 drain_left.n286 a_n1724_n5888# 5.65454f
C314 drain_left.n287 a_n1724_n5888# 0.371218f
C315 drain_left.t7 a_n1724_n5888# 0.613552f
C316 drain_left.t3 a_n1724_n5888# 0.613552f
C317 drain_left.n288 a_n1724_n5888# 5.65453f
C318 drain_left.n289 a_n1724_n5888# 0.629737f
C319 plus.n0 a_n1724_n5888# 0.052081f
C320 plus.t6 a_n1724_n5888# 1.09904f
C321 plus.t3 a_n1724_n5888# 1.09904f
C322 plus.t11 a_n1724_n5888# 1.09904f
C323 plus.n1 a_n1724_n5888# 0.417195f
C324 plus.n2 a_n1724_n5888# 0.122703f
C325 plus.t8 a_n1724_n5888# 1.09904f
C326 plus.t4 a_n1724_n5888# 1.09904f
C327 plus.t0 a_n1724_n5888# 1.1097f
C328 plus.n3 a_n1724_n5888# 0.416893f
C329 plus.n4 a_n1724_n5888# 0.399918f
C330 plus.n5 a_n1724_n5888# 0.021451f
C331 plus.n6 a_n1724_n5888# 0.399918f
C332 plus.n7 a_n1724_n5888# 0.021451f
C333 plus.n8 a_n1724_n5888# 0.052081f
C334 plus.n9 a_n1724_n5888# 0.052081f
C335 plus.n10 a_n1724_n5888# 0.052081f
C336 plus.n11 a_n1724_n5888# 0.021451f
C337 plus.n12 a_n1724_n5888# 0.399918f
C338 plus.n13 a_n1724_n5888# 0.021451f
C339 plus.n14 a_n1724_n5888# 0.399918f
C340 plus.t10 a_n1724_n5888# 1.1097f
C341 plus.n15 a_n1724_n5888# 0.416811f
C342 plus.n16 a_n1724_n5888# 0.93395f
C343 plus.n17 a_n1724_n5888# 0.052081f
C344 plus.t2 a_n1724_n5888# 1.1097f
C345 plus.t9 a_n1724_n5888# 1.09904f
C346 plus.t1 a_n1724_n5888# 1.09904f
C347 plus.t7 a_n1724_n5888# 1.09904f
C348 plus.n18 a_n1724_n5888# 0.417195f
C349 plus.n19 a_n1724_n5888# 0.122703f
C350 plus.t13 a_n1724_n5888# 1.09904f
C351 plus.t5 a_n1724_n5888# 1.09904f
C352 plus.t12 a_n1724_n5888# 1.1097f
C353 plus.n20 a_n1724_n5888# 0.416893f
C354 plus.n21 a_n1724_n5888# 0.399918f
C355 plus.n22 a_n1724_n5888# 0.021451f
C356 plus.n23 a_n1724_n5888# 0.399918f
C357 plus.n24 a_n1724_n5888# 0.021451f
C358 plus.n25 a_n1724_n5888# 0.052081f
C359 plus.n26 a_n1724_n5888# 0.052081f
C360 plus.n27 a_n1724_n5888# 0.052081f
C361 plus.n28 a_n1724_n5888# 0.021451f
C362 plus.n29 a_n1724_n5888# 0.399918f
C363 plus.n30 a_n1724_n5888# 0.021451f
C364 plus.n31 a_n1724_n5888# 0.399918f
C365 plus.n32 a_n1724_n5888# 0.416811f
C366 plus.n33 a_n1724_n5888# 1.98206f
C367 source.n0 a_n1724_n5888# 0.043231f
C368 source.n1 a_n1724_n5888# 0.031359f
C369 source.n2 a_n1724_n5888# 0.016851f
C370 source.n3 a_n1724_n5888# 0.039829f
C371 source.n4 a_n1724_n5888# 0.017842f
C372 source.n5 a_n1724_n5888# 0.031359f
C373 source.n6 a_n1724_n5888# 0.016851f
C374 source.n7 a_n1724_n5888# 0.039829f
C375 source.n8 a_n1724_n5888# 0.017842f
C376 source.n9 a_n1724_n5888# 0.031359f
C377 source.n10 a_n1724_n5888# 0.016851f
C378 source.n11 a_n1724_n5888# 0.039829f
C379 source.n12 a_n1724_n5888# 0.017842f
C380 source.n13 a_n1724_n5888# 0.031359f
C381 source.n14 a_n1724_n5888# 0.016851f
C382 source.n15 a_n1724_n5888# 0.039829f
C383 source.n16 a_n1724_n5888# 0.039829f
C384 source.n17 a_n1724_n5888# 0.017842f
C385 source.n18 a_n1724_n5888# 0.031359f
C386 source.n19 a_n1724_n5888# 0.016851f
C387 source.n20 a_n1724_n5888# 0.039829f
C388 source.n21 a_n1724_n5888# 0.017842f
C389 source.n22 a_n1724_n5888# 0.031359f
C390 source.n23 a_n1724_n5888# 0.016851f
C391 source.n24 a_n1724_n5888# 0.039829f
C392 source.n25 a_n1724_n5888# 0.017842f
C393 source.n26 a_n1724_n5888# 0.031359f
C394 source.n27 a_n1724_n5888# 0.016851f
C395 source.n28 a_n1724_n5888# 0.039829f
C396 source.n29 a_n1724_n5888# 0.017842f
C397 source.n30 a_n1724_n5888# 0.031359f
C398 source.n31 a_n1724_n5888# 0.016851f
C399 source.n32 a_n1724_n5888# 0.039829f
C400 source.n33 a_n1724_n5888# 0.017842f
C401 source.n34 a_n1724_n5888# 0.031359f
C402 source.n35 a_n1724_n5888# 0.017346f
C403 source.n36 a_n1724_n5888# 0.039829f
C404 source.n37 a_n1724_n5888# 0.016851f
C405 source.n38 a_n1724_n5888# 0.017842f
C406 source.n39 a_n1724_n5888# 0.031359f
C407 source.n40 a_n1724_n5888# 0.016851f
C408 source.n41 a_n1724_n5888# 0.039829f
C409 source.n42 a_n1724_n5888# 0.017842f
C410 source.n43 a_n1724_n5888# 0.031359f
C411 source.n44 a_n1724_n5888# 0.016851f
C412 source.n45 a_n1724_n5888# 0.029872f
C413 source.n46 a_n1724_n5888# 0.028156f
C414 source.t8 a_n1724_n5888# 0.069465f
C415 source.n47 a_n1724_n5888# 0.382605f
C416 source.n48 a_n1724_n5888# 3.39524f
C417 source.n49 a_n1724_n5888# 0.016851f
C418 source.n50 a_n1724_n5888# 0.017842f
C419 source.n51 a_n1724_n5888# 0.039829f
C420 source.n52 a_n1724_n5888# 0.039829f
C421 source.n53 a_n1724_n5888# 0.017842f
C422 source.n54 a_n1724_n5888# 0.016851f
C423 source.n55 a_n1724_n5888# 0.031359f
C424 source.n56 a_n1724_n5888# 0.031359f
C425 source.n57 a_n1724_n5888# 0.016851f
C426 source.n58 a_n1724_n5888# 0.017842f
C427 source.n59 a_n1724_n5888# 0.039829f
C428 source.n60 a_n1724_n5888# 0.039829f
C429 source.n61 a_n1724_n5888# 0.017842f
C430 source.n62 a_n1724_n5888# 0.016851f
C431 source.n63 a_n1724_n5888# 0.031359f
C432 source.n64 a_n1724_n5888# 0.031359f
C433 source.n65 a_n1724_n5888# 0.016851f
C434 source.n66 a_n1724_n5888# 0.017842f
C435 source.n67 a_n1724_n5888# 0.039829f
C436 source.n68 a_n1724_n5888# 0.039829f
C437 source.n69 a_n1724_n5888# 0.039829f
C438 source.n70 a_n1724_n5888# 0.017346f
C439 source.n71 a_n1724_n5888# 0.016851f
C440 source.n72 a_n1724_n5888# 0.031359f
C441 source.n73 a_n1724_n5888# 0.031359f
C442 source.n74 a_n1724_n5888# 0.016851f
C443 source.n75 a_n1724_n5888# 0.017842f
C444 source.n76 a_n1724_n5888# 0.039829f
C445 source.n77 a_n1724_n5888# 0.039829f
C446 source.n78 a_n1724_n5888# 0.017842f
C447 source.n79 a_n1724_n5888# 0.016851f
C448 source.n80 a_n1724_n5888# 0.031359f
C449 source.n81 a_n1724_n5888# 0.031359f
C450 source.n82 a_n1724_n5888# 0.016851f
C451 source.n83 a_n1724_n5888# 0.017842f
C452 source.n84 a_n1724_n5888# 0.039829f
C453 source.n85 a_n1724_n5888# 0.039829f
C454 source.n86 a_n1724_n5888# 0.017842f
C455 source.n87 a_n1724_n5888# 0.016851f
C456 source.n88 a_n1724_n5888# 0.031359f
C457 source.n89 a_n1724_n5888# 0.031359f
C458 source.n90 a_n1724_n5888# 0.016851f
C459 source.n91 a_n1724_n5888# 0.017842f
C460 source.n92 a_n1724_n5888# 0.039829f
C461 source.n93 a_n1724_n5888# 0.039829f
C462 source.n94 a_n1724_n5888# 0.017842f
C463 source.n95 a_n1724_n5888# 0.016851f
C464 source.n96 a_n1724_n5888# 0.031359f
C465 source.n97 a_n1724_n5888# 0.031359f
C466 source.n98 a_n1724_n5888# 0.016851f
C467 source.n99 a_n1724_n5888# 0.017842f
C468 source.n100 a_n1724_n5888# 0.039829f
C469 source.n101 a_n1724_n5888# 0.039829f
C470 source.n102 a_n1724_n5888# 0.017842f
C471 source.n103 a_n1724_n5888# 0.016851f
C472 source.n104 a_n1724_n5888# 0.031359f
C473 source.n105 a_n1724_n5888# 0.031359f
C474 source.n106 a_n1724_n5888# 0.016851f
C475 source.n107 a_n1724_n5888# 0.017842f
C476 source.n108 a_n1724_n5888# 0.039829f
C477 source.n109 a_n1724_n5888# 0.039829f
C478 source.n110 a_n1724_n5888# 0.017842f
C479 source.n111 a_n1724_n5888# 0.016851f
C480 source.n112 a_n1724_n5888# 0.031359f
C481 source.n113 a_n1724_n5888# 0.031359f
C482 source.n114 a_n1724_n5888# 0.016851f
C483 source.n115 a_n1724_n5888# 0.017346f
C484 source.n116 a_n1724_n5888# 0.017346f
C485 source.n117 a_n1724_n5888# 0.039829f
C486 source.n118 a_n1724_n5888# 0.039829f
C487 source.n119 a_n1724_n5888# 0.017842f
C488 source.n120 a_n1724_n5888# 0.016851f
C489 source.n121 a_n1724_n5888# 0.031359f
C490 source.n122 a_n1724_n5888# 0.031359f
C491 source.n123 a_n1724_n5888# 0.016851f
C492 source.n124 a_n1724_n5888# 0.017842f
C493 source.n125 a_n1724_n5888# 0.039829f
C494 source.n126 a_n1724_n5888# 0.039829f
C495 source.n127 a_n1724_n5888# 0.017842f
C496 source.n128 a_n1724_n5888# 0.016851f
C497 source.n129 a_n1724_n5888# 0.031359f
C498 source.n130 a_n1724_n5888# 0.031359f
C499 source.n131 a_n1724_n5888# 0.016851f
C500 source.n132 a_n1724_n5888# 0.017842f
C501 source.n133 a_n1724_n5888# 0.039829f
C502 source.n134 a_n1724_n5888# 0.084727f
C503 source.n135 a_n1724_n5888# 0.017842f
C504 source.n136 a_n1724_n5888# 0.016851f
C505 source.n137 a_n1724_n5888# 0.069057f
C506 source.n138 a_n1724_n5888# 0.047147f
C507 source.n139 a_n1724_n5888# 2.46456f
C508 source.t1 a_n1724_n5888# 0.619518f
C509 source.t6 a_n1724_n5888# 0.619518f
C510 source.n140 a_n1724_n5888# 5.60673f
C511 source.n141 a_n1724_n5888# 0.43501f
C512 source.t13 a_n1724_n5888# 0.619518f
C513 source.t11 a_n1724_n5888# 0.619518f
C514 source.n142 a_n1724_n5888# 5.60673f
C515 source.n143 a_n1724_n5888# 0.43501f
C516 source.t7 a_n1724_n5888# 0.619518f
C517 source.t4 a_n1724_n5888# 0.619518f
C518 source.n144 a_n1724_n5888# 5.60673f
C519 source.n145 a_n1724_n5888# 0.455045f
C520 source.n146 a_n1724_n5888# 0.043231f
C521 source.n147 a_n1724_n5888# 0.031359f
C522 source.n148 a_n1724_n5888# 0.016851f
C523 source.n149 a_n1724_n5888# 0.039829f
C524 source.n150 a_n1724_n5888# 0.017842f
C525 source.n151 a_n1724_n5888# 0.031359f
C526 source.n152 a_n1724_n5888# 0.016851f
C527 source.n153 a_n1724_n5888# 0.039829f
C528 source.n154 a_n1724_n5888# 0.017842f
C529 source.n155 a_n1724_n5888# 0.031359f
C530 source.n156 a_n1724_n5888# 0.016851f
C531 source.n157 a_n1724_n5888# 0.039829f
C532 source.n158 a_n1724_n5888# 0.017842f
C533 source.n159 a_n1724_n5888# 0.031359f
C534 source.n160 a_n1724_n5888# 0.016851f
C535 source.n161 a_n1724_n5888# 0.039829f
C536 source.n162 a_n1724_n5888# 0.039829f
C537 source.n163 a_n1724_n5888# 0.017842f
C538 source.n164 a_n1724_n5888# 0.031359f
C539 source.n165 a_n1724_n5888# 0.016851f
C540 source.n166 a_n1724_n5888# 0.039829f
C541 source.n167 a_n1724_n5888# 0.017842f
C542 source.n168 a_n1724_n5888# 0.031359f
C543 source.n169 a_n1724_n5888# 0.016851f
C544 source.n170 a_n1724_n5888# 0.039829f
C545 source.n171 a_n1724_n5888# 0.017842f
C546 source.n172 a_n1724_n5888# 0.031359f
C547 source.n173 a_n1724_n5888# 0.016851f
C548 source.n174 a_n1724_n5888# 0.039829f
C549 source.n175 a_n1724_n5888# 0.017842f
C550 source.n176 a_n1724_n5888# 0.031359f
C551 source.n177 a_n1724_n5888# 0.016851f
C552 source.n178 a_n1724_n5888# 0.039829f
C553 source.n179 a_n1724_n5888# 0.017842f
C554 source.n180 a_n1724_n5888# 0.031359f
C555 source.n181 a_n1724_n5888# 0.017346f
C556 source.n182 a_n1724_n5888# 0.039829f
C557 source.n183 a_n1724_n5888# 0.016851f
C558 source.n184 a_n1724_n5888# 0.017842f
C559 source.n185 a_n1724_n5888# 0.031359f
C560 source.n186 a_n1724_n5888# 0.016851f
C561 source.n187 a_n1724_n5888# 0.039829f
C562 source.n188 a_n1724_n5888# 0.017842f
C563 source.n189 a_n1724_n5888# 0.031359f
C564 source.n190 a_n1724_n5888# 0.016851f
C565 source.n191 a_n1724_n5888# 0.029872f
C566 source.n192 a_n1724_n5888# 0.028156f
C567 source.t19 a_n1724_n5888# 0.069465f
C568 source.n193 a_n1724_n5888# 0.382605f
C569 source.n194 a_n1724_n5888# 3.39524f
C570 source.n195 a_n1724_n5888# 0.016851f
C571 source.n196 a_n1724_n5888# 0.017842f
C572 source.n197 a_n1724_n5888# 0.039829f
C573 source.n198 a_n1724_n5888# 0.039829f
C574 source.n199 a_n1724_n5888# 0.017842f
C575 source.n200 a_n1724_n5888# 0.016851f
C576 source.n201 a_n1724_n5888# 0.031359f
C577 source.n202 a_n1724_n5888# 0.031359f
C578 source.n203 a_n1724_n5888# 0.016851f
C579 source.n204 a_n1724_n5888# 0.017842f
C580 source.n205 a_n1724_n5888# 0.039829f
C581 source.n206 a_n1724_n5888# 0.039829f
C582 source.n207 a_n1724_n5888# 0.017842f
C583 source.n208 a_n1724_n5888# 0.016851f
C584 source.n209 a_n1724_n5888# 0.031359f
C585 source.n210 a_n1724_n5888# 0.031359f
C586 source.n211 a_n1724_n5888# 0.016851f
C587 source.n212 a_n1724_n5888# 0.017842f
C588 source.n213 a_n1724_n5888# 0.039829f
C589 source.n214 a_n1724_n5888# 0.039829f
C590 source.n215 a_n1724_n5888# 0.039829f
C591 source.n216 a_n1724_n5888# 0.017346f
C592 source.n217 a_n1724_n5888# 0.016851f
C593 source.n218 a_n1724_n5888# 0.031359f
C594 source.n219 a_n1724_n5888# 0.031359f
C595 source.n220 a_n1724_n5888# 0.016851f
C596 source.n221 a_n1724_n5888# 0.017842f
C597 source.n222 a_n1724_n5888# 0.039829f
C598 source.n223 a_n1724_n5888# 0.039829f
C599 source.n224 a_n1724_n5888# 0.017842f
C600 source.n225 a_n1724_n5888# 0.016851f
C601 source.n226 a_n1724_n5888# 0.031359f
C602 source.n227 a_n1724_n5888# 0.031359f
C603 source.n228 a_n1724_n5888# 0.016851f
C604 source.n229 a_n1724_n5888# 0.017842f
C605 source.n230 a_n1724_n5888# 0.039829f
C606 source.n231 a_n1724_n5888# 0.039829f
C607 source.n232 a_n1724_n5888# 0.017842f
C608 source.n233 a_n1724_n5888# 0.016851f
C609 source.n234 a_n1724_n5888# 0.031359f
C610 source.n235 a_n1724_n5888# 0.031359f
C611 source.n236 a_n1724_n5888# 0.016851f
C612 source.n237 a_n1724_n5888# 0.017842f
C613 source.n238 a_n1724_n5888# 0.039829f
C614 source.n239 a_n1724_n5888# 0.039829f
C615 source.n240 a_n1724_n5888# 0.017842f
C616 source.n241 a_n1724_n5888# 0.016851f
C617 source.n242 a_n1724_n5888# 0.031359f
C618 source.n243 a_n1724_n5888# 0.031359f
C619 source.n244 a_n1724_n5888# 0.016851f
C620 source.n245 a_n1724_n5888# 0.017842f
C621 source.n246 a_n1724_n5888# 0.039829f
C622 source.n247 a_n1724_n5888# 0.039829f
C623 source.n248 a_n1724_n5888# 0.017842f
C624 source.n249 a_n1724_n5888# 0.016851f
C625 source.n250 a_n1724_n5888# 0.031359f
C626 source.n251 a_n1724_n5888# 0.031359f
C627 source.n252 a_n1724_n5888# 0.016851f
C628 source.n253 a_n1724_n5888# 0.017842f
C629 source.n254 a_n1724_n5888# 0.039829f
C630 source.n255 a_n1724_n5888# 0.039829f
C631 source.n256 a_n1724_n5888# 0.017842f
C632 source.n257 a_n1724_n5888# 0.016851f
C633 source.n258 a_n1724_n5888# 0.031359f
C634 source.n259 a_n1724_n5888# 0.031359f
C635 source.n260 a_n1724_n5888# 0.016851f
C636 source.n261 a_n1724_n5888# 0.017346f
C637 source.n262 a_n1724_n5888# 0.017346f
C638 source.n263 a_n1724_n5888# 0.039829f
C639 source.n264 a_n1724_n5888# 0.039829f
C640 source.n265 a_n1724_n5888# 0.017842f
C641 source.n266 a_n1724_n5888# 0.016851f
C642 source.n267 a_n1724_n5888# 0.031359f
C643 source.n268 a_n1724_n5888# 0.031359f
C644 source.n269 a_n1724_n5888# 0.016851f
C645 source.n270 a_n1724_n5888# 0.017842f
C646 source.n271 a_n1724_n5888# 0.039829f
C647 source.n272 a_n1724_n5888# 0.039829f
C648 source.n273 a_n1724_n5888# 0.017842f
C649 source.n274 a_n1724_n5888# 0.016851f
C650 source.n275 a_n1724_n5888# 0.031359f
C651 source.n276 a_n1724_n5888# 0.031359f
C652 source.n277 a_n1724_n5888# 0.016851f
C653 source.n278 a_n1724_n5888# 0.017842f
C654 source.n279 a_n1724_n5888# 0.039829f
C655 source.n280 a_n1724_n5888# 0.084727f
C656 source.n281 a_n1724_n5888# 0.017842f
C657 source.n282 a_n1724_n5888# 0.016851f
C658 source.n283 a_n1724_n5888# 0.069057f
C659 source.n284 a_n1724_n5888# 0.047147f
C660 source.n285 a_n1724_n5888# 0.154642f
C661 source.t26 a_n1724_n5888# 0.619518f
C662 source.t15 a_n1724_n5888# 0.619518f
C663 source.n286 a_n1724_n5888# 5.60673f
C664 source.n287 a_n1724_n5888# 0.43501f
C665 source.t16 a_n1724_n5888# 0.619518f
C666 source.t20 a_n1724_n5888# 0.619518f
C667 source.n288 a_n1724_n5888# 5.60673f
C668 source.n289 a_n1724_n5888# 0.43501f
C669 source.t23 a_n1724_n5888# 0.619518f
C670 source.t27 a_n1724_n5888# 0.619518f
C671 source.n290 a_n1724_n5888# 5.60673f
C672 source.n291 a_n1724_n5888# 3.39997f
C673 source.t0 a_n1724_n5888# 0.619518f
C674 source.t5 a_n1724_n5888# 0.619518f
C675 source.n292 a_n1724_n5888# 5.60673f
C676 source.n293 a_n1724_n5888# 3.39997f
C677 source.t2 a_n1724_n5888# 0.619518f
C678 source.t12 a_n1724_n5888# 0.619518f
C679 source.n294 a_n1724_n5888# 5.60673f
C680 source.n295 a_n1724_n5888# 0.435012f
C681 source.t9 a_n1724_n5888# 0.619518f
C682 source.t10 a_n1724_n5888# 0.619518f
C683 source.n296 a_n1724_n5888# 5.60673f
C684 source.n297 a_n1724_n5888# 0.435012f
C685 source.n298 a_n1724_n5888# 0.043231f
C686 source.n299 a_n1724_n5888# 0.031359f
C687 source.n300 a_n1724_n5888# 0.016851f
C688 source.n301 a_n1724_n5888# 0.039829f
C689 source.n302 a_n1724_n5888# 0.017842f
C690 source.n303 a_n1724_n5888# 0.031359f
C691 source.n304 a_n1724_n5888# 0.016851f
C692 source.n305 a_n1724_n5888# 0.039829f
C693 source.n306 a_n1724_n5888# 0.017842f
C694 source.n307 a_n1724_n5888# 0.031359f
C695 source.n308 a_n1724_n5888# 0.016851f
C696 source.n309 a_n1724_n5888# 0.039829f
C697 source.n310 a_n1724_n5888# 0.017842f
C698 source.n311 a_n1724_n5888# 0.031359f
C699 source.n312 a_n1724_n5888# 0.016851f
C700 source.n313 a_n1724_n5888# 0.039829f
C701 source.n314 a_n1724_n5888# 0.017842f
C702 source.n315 a_n1724_n5888# 0.031359f
C703 source.n316 a_n1724_n5888# 0.016851f
C704 source.n317 a_n1724_n5888# 0.039829f
C705 source.n318 a_n1724_n5888# 0.017842f
C706 source.n319 a_n1724_n5888# 0.031359f
C707 source.n320 a_n1724_n5888# 0.016851f
C708 source.n321 a_n1724_n5888# 0.039829f
C709 source.n322 a_n1724_n5888# 0.017842f
C710 source.n323 a_n1724_n5888# 0.031359f
C711 source.n324 a_n1724_n5888# 0.016851f
C712 source.n325 a_n1724_n5888# 0.039829f
C713 source.n326 a_n1724_n5888# 0.017842f
C714 source.n327 a_n1724_n5888# 0.031359f
C715 source.n328 a_n1724_n5888# 0.016851f
C716 source.n329 a_n1724_n5888# 0.039829f
C717 source.n330 a_n1724_n5888# 0.017842f
C718 source.n331 a_n1724_n5888# 0.031359f
C719 source.n332 a_n1724_n5888# 0.017346f
C720 source.n333 a_n1724_n5888# 0.039829f
C721 source.n334 a_n1724_n5888# 0.017842f
C722 source.n335 a_n1724_n5888# 0.031359f
C723 source.n336 a_n1724_n5888# 0.016851f
C724 source.n337 a_n1724_n5888# 0.039829f
C725 source.n338 a_n1724_n5888# 0.017842f
C726 source.n339 a_n1724_n5888# 0.031359f
C727 source.n340 a_n1724_n5888# 0.016851f
C728 source.n341 a_n1724_n5888# 0.029872f
C729 source.n342 a_n1724_n5888# 0.028156f
C730 source.t3 a_n1724_n5888# 0.069465f
C731 source.n343 a_n1724_n5888# 0.382605f
C732 source.n344 a_n1724_n5888# 3.39524f
C733 source.n345 a_n1724_n5888# 0.016851f
C734 source.n346 a_n1724_n5888# 0.017842f
C735 source.n347 a_n1724_n5888# 0.039829f
C736 source.n348 a_n1724_n5888# 0.039829f
C737 source.n349 a_n1724_n5888# 0.017842f
C738 source.n350 a_n1724_n5888# 0.016851f
C739 source.n351 a_n1724_n5888# 0.031359f
C740 source.n352 a_n1724_n5888# 0.031359f
C741 source.n353 a_n1724_n5888# 0.016851f
C742 source.n354 a_n1724_n5888# 0.017842f
C743 source.n355 a_n1724_n5888# 0.039829f
C744 source.n356 a_n1724_n5888# 0.039829f
C745 source.n357 a_n1724_n5888# 0.017842f
C746 source.n358 a_n1724_n5888# 0.016851f
C747 source.n359 a_n1724_n5888# 0.031359f
C748 source.n360 a_n1724_n5888# 0.031359f
C749 source.n361 a_n1724_n5888# 0.016851f
C750 source.n362 a_n1724_n5888# 0.016851f
C751 source.n363 a_n1724_n5888# 0.017842f
C752 source.n364 a_n1724_n5888# 0.039829f
C753 source.n365 a_n1724_n5888# 0.039829f
C754 source.n366 a_n1724_n5888# 0.039829f
C755 source.n367 a_n1724_n5888# 0.017346f
C756 source.n368 a_n1724_n5888# 0.016851f
C757 source.n369 a_n1724_n5888# 0.031359f
C758 source.n370 a_n1724_n5888# 0.031359f
C759 source.n371 a_n1724_n5888# 0.016851f
C760 source.n372 a_n1724_n5888# 0.017842f
C761 source.n373 a_n1724_n5888# 0.039829f
C762 source.n374 a_n1724_n5888# 0.039829f
C763 source.n375 a_n1724_n5888# 0.017842f
C764 source.n376 a_n1724_n5888# 0.016851f
C765 source.n377 a_n1724_n5888# 0.031359f
C766 source.n378 a_n1724_n5888# 0.031359f
C767 source.n379 a_n1724_n5888# 0.016851f
C768 source.n380 a_n1724_n5888# 0.017842f
C769 source.n381 a_n1724_n5888# 0.039829f
C770 source.n382 a_n1724_n5888# 0.039829f
C771 source.n383 a_n1724_n5888# 0.017842f
C772 source.n384 a_n1724_n5888# 0.016851f
C773 source.n385 a_n1724_n5888# 0.031359f
C774 source.n386 a_n1724_n5888# 0.031359f
C775 source.n387 a_n1724_n5888# 0.016851f
C776 source.n388 a_n1724_n5888# 0.017842f
C777 source.n389 a_n1724_n5888# 0.039829f
C778 source.n390 a_n1724_n5888# 0.039829f
C779 source.n391 a_n1724_n5888# 0.017842f
C780 source.n392 a_n1724_n5888# 0.016851f
C781 source.n393 a_n1724_n5888# 0.031359f
C782 source.n394 a_n1724_n5888# 0.031359f
C783 source.n395 a_n1724_n5888# 0.016851f
C784 source.n396 a_n1724_n5888# 0.017842f
C785 source.n397 a_n1724_n5888# 0.039829f
C786 source.n398 a_n1724_n5888# 0.039829f
C787 source.n399 a_n1724_n5888# 0.017842f
C788 source.n400 a_n1724_n5888# 0.016851f
C789 source.n401 a_n1724_n5888# 0.031359f
C790 source.n402 a_n1724_n5888# 0.031359f
C791 source.n403 a_n1724_n5888# 0.016851f
C792 source.n404 a_n1724_n5888# 0.017842f
C793 source.n405 a_n1724_n5888# 0.039829f
C794 source.n406 a_n1724_n5888# 0.039829f
C795 source.n407 a_n1724_n5888# 0.039829f
C796 source.n408 a_n1724_n5888# 0.017842f
C797 source.n409 a_n1724_n5888# 0.016851f
C798 source.n410 a_n1724_n5888# 0.031359f
C799 source.n411 a_n1724_n5888# 0.031359f
C800 source.n412 a_n1724_n5888# 0.016851f
C801 source.n413 a_n1724_n5888# 0.017346f
C802 source.n414 a_n1724_n5888# 0.017346f
C803 source.n415 a_n1724_n5888# 0.039829f
C804 source.n416 a_n1724_n5888# 0.039829f
C805 source.n417 a_n1724_n5888# 0.017842f
C806 source.n418 a_n1724_n5888# 0.016851f
C807 source.n419 a_n1724_n5888# 0.031359f
C808 source.n420 a_n1724_n5888# 0.031359f
C809 source.n421 a_n1724_n5888# 0.016851f
C810 source.n422 a_n1724_n5888# 0.017842f
C811 source.n423 a_n1724_n5888# 0.039829f
C812 source.n424 a_n1724_n5888# 0.039829f
C813 source.n425 a_n1724_n5888# 0.017842f
C814 source.n426 a_n1724_n5888# 0.016851f
C815 source.n427 a_n1724_n5888# 0.031359f
C816 source.n428 a_n1724_n5888# 0.031359f
C817 source.n429 a_n1724_n5888# 0.016851f
C818 source.n430 a_n1724_n5888# 0.017842f
C819 source.n431 a_n1724_n5888# 0.039829f
C820 source.n432 a_n1724_n5888# 0.084727f
C821 source.n433 a_n1724_n5888# 0.017842f
C822 source.n434 a_n1724_n5888# 0.016851f
C823 source.n435 a_n1724_n5888# 0.069057f
C824 source.n436 a_n1724_n5888# 0.047147f
C825 source.n437 a_n1724_n5888# 0.154642f
C826 source.t24 a_n1724_n5888# 0.619518f
C827 source.t17 a_n1724_n5888# 0.619518f
C828 source.n438 a_n1724_n5888# 5.60673f
C829 source.n439 a_n1724_n5888# 0.455047f
C830 source.t25 a_n1724_n5888# 0.619518f
C831 source.t18 a_n1724_n5888# 0.619518f
C832 source.n440 a_n1724_n5888# 5.60673f
C833 source.n441 a_n1724_n5888# 0.435012f
C834 source.t21 a_n1724_n5888# 0.619518f
C835 source.t14 a_n1724_n5888# 0.619518f
C836 source.n442 a_n1724_n5888# 5.60673f
C837 source.n443 a_n1724_n5888# 0.435012f
C838 source.n444 a_n1724_n5888# 0.043231f
C839 source.n445 a_n1724_n5888# 0.031359f
C840 source.n446 a_n1724_n5888# 0.016851f
C841 source.n447 a_n1724_n5888# 0.039829f
C842 source.n448 a_n1724_n5888# 0.017842f
C843 source.n449 a_n1724_n5888# 0.031359f
C844 source.n450 a_n1724_n5888# 0.016851f
C845 source.n451 a_n1724_n5888# 0.039829f
C846 source.n452 a_n1724_n5888# 0.017842f
C847 source.n453 a_n1724_n5888# 0.031359f
C848 source.n454 a_n1724_n5888# 0.016851f
C849 source.n455 a_n1724_n5888# 0.039829f
C850 source.n456 a_n1724_n5888# 0.017842f
C851 source.n457 a_n1724_n5888# 0.031359f
C852 source.n458 a_n1724_n5888# 0.016851f
C853 source.n459 a_n1724_n5888# 0.039829f
C854 source.n460 a_n1724_n5888# 0.017842f
C855 source.n461 a_n1724_n5888# 0.031359f
C856 source.n462 a_n1724_n5888# 0.016851f
C857 source.n463 a_n1724_n5888# 0.039829f
C858 source.n464 a_n1724_n5888# 0.017842f
C859 source.n465 a_n1724_n5888# 0.031359f
C860 source.n466 a_n1724_n5888# 0.016851f
C861 source.n467 a_n1724_n5888# 0.039829f
C862 source.n468 a_n1724_n5888# 0.017842f
C863 source.n469 a_n1724_n5888# 0.031359f
C864 source.n470 a_n1724_n5888# 0.016851f
C865 source.n471 a_n1724_n5888# 0.039829f
C866 source.n472 a_n1724_n5888# 0.017842f
C867 source.n473 a_n1724_n5888# 0.031359f
C868 source.n474 a_n1724_n5888# 0.016851f
C869 source.n475 a_n1724_n5888# 0.039829f
C870 source.n476 a_n1724_n5888# 0.017842f
C871 source.n477 a_n1724_n5888# 0.031359f
C872 source.n478 a_n1724_n5888# 0.017346f
C873 source.n479 a_n1724_n5888# 0.039829f
C874 source.n480 a_n1724_n5888# 0.017842f
C875 source.n481 a_n1724_n5888# 0.031359f
C876 source.n482 a_n1724_n5888# 0.016851f
C877 source.n483 a_n1724_n5888# 0.039829f
C878 source.n484 a_n1724_n5888# 0.017842f
C879 source.n485 a_n1724_n5888# 0.031359f
C880 source.n486 a_n1724_n5888# 0.016851f
C881 source.n487 a_n1724_n5888# 0.029872f
C882 source.n488 a_n1724_n5888# 0.028156f
C883 source.t22 a_n1724_n5888# 0.069465f
C884 source.n489 a_n1724_n5888# 0.382605f
C885 source.n490 a_n1724_n5888# 3.39524f
C886 source.n491 a_n1724_n5888# 0.016851f
C887 source.n492 a_n1724_n5888# 0.017842f
C888 source.n493 a_n1724_n5888# 0.039829f
C889 source.n494 a_n1724_n5888# 0.039829f
C890 source.n495 a_n1724_n5888# 0.017842f
C891 source.n496 a_n1724_n5888# 0.016851f
C892 source.n497 a_n1724_n5888# 0.031359f
C893 source.n498 a_n1724_n5888# 0.031359f
C894 source.n499 a_n1724_n5888# 0.016851f
C895 source.n500 a_n1724_n5888# 0.017842f
C896 source.n501 a_n1724_n5888# 0.039829f
C897 source.n502 a_n1724_n5888# 0.039829f
C898 source.n503 a_n1724_n5888# 0.017842f
C899 source.n504 a_n1724_n5888# 0.016851f
C900 source.n505 a_n1724_n5888# 0.031359f
C901 source.n506 a_n1724_n5888# 0.031359f
C902 source.n507 a_n1724_n5888# 0.016851f
C903 source.n508 a_n1724_n5888# 0.016851f
C904 source.n509 a_n1724_n5888# 0.017842f
C905 source.n510 a_n1724_n5888# 0.039829f
C906 source.n511 a_n1724_n5888# 0.039829f
C907 source.n512 a_n1724_n5888# 0.039829f
C908 source.n513 a_n1724_n5888# 0.017346f
C909 source.n514 a_n1724_n5888# 0.016851f
C910 source.n515 a_n1724_n5888# 0.031359f
C911 source.n516 a_n1724_n5888# 0.031359f
C912 source.n517 a_n1724_n5888# 0.016851f
C913 source.n518 a_n1724_n5888# 0.017842f
C914 source.n519 a_n1724_n5888# 0.039829f
C915 source.n520 a_n1724_n5888# 0.039829f
C916 source.n521 a_n1724_n5888# 0.017842f
C917 source.n522 a_n1724_n5888# 0.016851f
C918 source.n523 a_n1724_n5888# 0.031359f
C919 source.n524 a_n1724_n5888# 0.031359f
C920 source.n525 a_n1724_n5888# 0.016851f
C921 source.n526 a_n1724_n5888# 0.017842f
C922 source.n527 a_n1724_n5888# 0.039829f
C923 source.n528 a_n1724_n5888# 0.039829f
C924 source.n529 a_n1724_n5888# 0.017842f
C925 source.n530 a_n1724_n5888# 0.016851f
C926 source.n531 a_n1724_n5888# 0.031359f
C927 source.n532 a_n1724_n5888# 0.031359f
C928 source.n533 a_n1724_n5888# 0.016851f
C929 source.n534 a_n1724_n5888# 0.017842f
C930 source.n535 a_n1724_n5888# 0.039829f
C931 source.n536 a_n1724_n5888# 0.039829f
C932 source.n537 a_n1724_n5888# 0.017842f
C933 source.n538 a_n1724_n5888# 0.016851f
C934 source.n539 a_n1724_n5888# 0.031359f
C935 source.n540 a_n1724_n5888# 0.031359f
C936 source.n541 a_n1724_n5888# 0.016851f
C937 source.n542 a_n1724_n5888# 0.017842f
C938 source.n543 a_n1724_n5888# 0.039829f
C939 source.n544 a_n1724_n5888# 0.039829f
C940 source.n545 a_n1724_n5888# 0.017842f
C941 source.n546 a_n1724_n5888# 0.016851f
C942 source.n547 a_n1724_n5888# 0.031359f
C943 source.n548 a_n1724_n5888# 0.031359f
C944 source.n549 a_n1724_n5888# 0.016851f
C945 source.n550 a_n1724_n5888# 0.017842f
C946 source.n551 a_n1724_n5888# 0.039829f
C947 source.n552 a_n1724_n5888# 0.039829f
C948 source.n553 a_n1724_n5888# 0.039829f
C949 source.n554 a_n1724_n5888# 0.017842f
C950 source.n555 a_n1724_n5888# 0.016851f
C951 source.n556 a_n1724_n5888# 0.031359f
C952 source.n557 a_n1724_n5888# 0.031359f
C953 source.n558 a_n1724_n5888# 0.016851f
C954 source.n559 a_n1724_n5888# 0.017346f
C955 source.n560 a_n1724_n5888# 0.017346f
C956 source.n561 a_n1724_n5888# 0.039829f
C957 source.n562 a_n1724_n5888# 0.039829f
C958 source.n563 a_n1724_n5888# 0.017842f
C959 source.n564 a_n1724_n5888# 0.016851f
C960 source.n565 a_n1724_n5888# 0.031359f
C961 source.n566 a_n1724_n5888# 0.031359f
C962 source.n567 a_n1724_n5888# 0.016851f
C963 source.n568 a_n1724_n5888# 0.017842f
C964 source.n569 a_n1724_n5888# 0.039829f
C965 source.n570 a_n1724_n5888# 0.039829f
C966 source.n571 a_n1724_n5888# 0.017842f
C967 source.n572 a_n1724_n5888# 0.016851f
C968 source.n573 a_n1724_n5888# 0.031359f
C969 source.n574 a_n1724_n5888# 0.031359f
C970 source.n575 a_n1724_n5888# 0.016851f
C971 source.n576 a_n1724_n5888# 0.017842f
C972 source.n577 a_n1724_n5888# 0.039829f
C973 source.n578 a_n1724_n5888# 0.084727f
C974 source.n579 a_n1724_n5888# 0.017842f
C975 source.n580 a_n1724_n5888# 0.016851f
C976 source.n581 a_n1724_n5888# 0.069057f
C977 source.n582 a_n1724_n5888# 0.047147f
C978 source.n583 a_n1724_n5888# 0.304223f
C979 source.n584 a_n1724_n5888# 3.3429f
C980 drain_right.n0 a_n1724_n5888# 0.042829f
C981 drain_right.n1 a_n1724_n5888# 0.031067f
C982 drain_right.n2 a_n1724_n5888# 0.016694f
C983 drain_right.n3 a_n1724_n5888# 0.039459f
C984 drain_right.n4 a_n1724_n5888# 0.017676f
C985 drain_right.n5 a_n1724_n5888# 0.031067f
C986 drain_right.n6 a_n1724_n5888# 0.016694f
C987 drain_right.n7 a_n1724_n5888# 0.039459f
C988 drain_right.n8 a_n1724_n5888# 0.017676f
C989 drain_right.n9 a_n1724_n5888# 0.031067f
C990 drain_right.n10 a_n1724_n5888# 0.016694f
C991 drain_right.n11 a_n1724_n5888# 0.039459f
C992 drain_right.n12 a_n1724_n5888# 0.017676f
C993 drain_right.n13 a_n1724_n5888# 0.031067f
C994 drain_right.n14 a_n1724_n5888# 0.016694f
C995 drain_right.n15 a_n1724_n5888# 0.039459f
C996 drain_right.n16 a_n1724_n5888# 0.017676f
C997 drain_right.n17 a_n1724_n5888# 0.031067f
C998 drain_right.n18 a_n1724_n5888# 0.016694f
C999 drain_right.n19 a_n1724_n5888# 0.039459f
C1000 drain_right.n20 a_n1724_n5888# 0.017676f
C1001 drain_right.n21 a_n1724_n5888# 0.031067f
C1002 drain_right.n22 a_n1724_n5888# 0.016694f
C1003 drain_right.n23 a_n1724_n5888# 0.039459f
C1004 drain_right.n24 a_n1724_n5888# 0.017676f
C1005 drain_right.n25 a_n1724_n5888# 0.031067f
C1006 drain_right.n26 a_n1724_n5888# 0.016694f
C1007 drain_right.n27 a_n1724_n5888# 0.039459f
C1008 drain_right.n28 a_n1724_n5888# 0.017676f
C1009 drain_right.n29 a_n1724_n5888# 0.031067f
C1010 drain_right.n30 a_n1724_n5888# 0.016694f
C1011 drain_right.n31 a_n1724_n5888# 0.039459f
C1012 drain_right.n32 a_n1724_n5888# 0.017676f
C1013 drain_right.n33 a_n1724_n5888# 0.031067f
C1014 drain_right.n34 a_n1724_n5888# 0.017185f
C1015 drain_right.n35 a_n1724_n5888# 0.039459f
C1016 drain_right.n36 a_n1724_n5888# 0.017676f
C1017 drain_right.n37 a_n1724_n5888# 0.031067f
C1018 drain_right.n38 a_n1724_n5888# 0.016694f
C1019 drain_right.n39 a_n1724_n5888# 0.039459f
C1020 drain_right.n40 a_n1724_n5888# 0.017676f
C1021 drain_right.n41 a_n1724_n5888# 0.031067f
C1022 drain_right.n42 a_n1724_n5888# 0.016694f
C1023 drain_right.n43 a_n1724_n5888# 0.029594f
C1024 drain_right.n44 a_n1724_n5888# 0.027894f
C1025 drain_right.t2 a_n1724_n5888# 0.068818f
C1026 drain_right.n45 a_n1724_n5888# 0.379043f
C1027 drain_right.n46 a_n1724_n5888# 3.36364f
C1028 drain_right.n47 a_n1724_n5888# 0.016694f
C1029 drain_right.n48 a_n1724_n5888# 0.017676f
C1030 drain_right.n49 a_n1724_n5888# 0.039459f
C1031 drain_right.n50 a_n1724_n5888# 0.039459f
C1032 drain_right.n51 a_n1724_n5888# 0.017676f
C1033 drain_right.n52 a_n1724_n5888# 0.016694f
C1034 drain_right.n53 a_n1724_n5888# 0.031067f
C1035 drain_right.n54 a_n1724_n5888# 0.031067f
C1036 drain_right.n55 a_n1724_n5888# 0.016694f
C1037 drain_right.n56 a_n1724_n5888# 0.017676f
C1038 drain_right.n57 a_n1724_n5888# 0.039459f
C1039 drain_right.n58 a_n1724_n5888# 0.039459f
C1040 drain_right.n59 a_n1724_n5888# 0.017676f
C1041 drain_right.n60 a_n1724_n5888# 0.016694f
C1042 drain_right.n61 a_n1724_n5888# 0.031067f
C1043 drain_right.n62 a_n1724_n5888# 0.031067f
C1044 drain_right.n63 a_n1724_n5888# 0.016694f
C1045 drain_right.n64 a_n1724_n5888# 0.016694f
C1046 drain_right.n65 a_n1724_n5888# 0.017676f
C1047 drain_right.n66 a_n1724_n5888# 0.039459f
C1048 drain_right.n67 a_n1724_n5888# 0.039459f
C1049 drain_right.n68 a_n1724_n5888# 0.039459f
C1050 drain_right.n69 a_n1724_n5888# 0.017185f
C1051 drain_right.n70 a_n1724_n5888# 0.016694f
C1052 drain_right.n71 a_n1724_n5888# 0.031067f
C1053 drain_right.n72 a_n1724_n5888# 0.031067f
C1054 drain_right.n73 a_n1724_n5888# 0.016694f
C1055 drain_right.n74 a_n1724_n5888# 0.017676f
C1056 drain_right.n75 a_n1724_n5888# 0.039459f
C1057 drain_right.n76 a_n1724_n5888# 0.039459f
C1058 drain_right.n77 a_n1724_n5888# 0.017676f
C1059 drain_right.n78 a_n1724_n5888# 0.016694f
C1060 drain_right.n79 a_n1724_n5888# 0.031067f
C1061 drain_right.n80 a_n1724_n5888# 0.031067f
C1062 drain_right.n81 a_n1724_n5888# 0.016694f
C1063 drain_right.n82 a_n1724_n5888# 0.017676f
C1064 drain_right.n83 a_n1724_n5888# 0.039459f
C1065 drain_right.n84 a_n1724_n5888# 0.039459f
C1066 drain_right.n85 a_n1724_n5888# 0.017676f
C1067 drain_right.n86 a_n1724_n5888# 0.016694f
C1068 drain_right.n87 a_n1724_n5888# 0.031067f
C1069 drain_right.n88 a_n1724_n5888# 0.031067f
C1070 drain_right.n89 a_n1724_n5888# 0.016694f
C1071 drain_right.n90 a_n1724_n5888# 0.017676f
C1072 drain_right.n91 a_n1724_n5888# 0.039459f
C1073 drain_right.n92 a_n1724_n5888# 0.039459f
C1074 drain_right.n93 a_n1724_n5888# 0.017676f
C1075 drain_right.n94 a_n1724_n5888# 0.016694f
C1076 drain_right.n95 a_n1724_n5888# 0.031067f
C1077 drain_right.n96 a_n1724_n5888# 0.031067f
C1078 drain_right.n97 a_n1724_n5888# 0.016694f
C1079 drain_right.n98 a_n1724_n5888# 0.017676f
C1080 drain_right.n99 a_n1724_n5888# 0.039459f
C1081 drain_right.n100 a_n1724_n5888# 0.039459f
C1082 drain_right.n101 a_n1724_n5888# 0.017676f
C1083 drain_right.n102 a_n1724_n5888# 0.016694f
C1084 drain_right.n103 a_n1724_n5888# 0.031067f
C1085 drain_right.n104 a_n1724_n5888# 0.031067f
C1086 drain_right.n105 a_n1724_n5888# 0.016694f
C1087 drain_right.n106 a_n1724_n5888# 0.017676f
C1088 drain_right.n107 a_n1724_n5888# 0.039459f
C1089 drain_right.n108 a_n1724_n5888# 0.039459f
C1090 drain_right.n109 a_n1724_n5888# 0.039459f
C1091 drain_right.n110 a_n1724_n5888# 0.017676f
C1092 drain_right.n111 a_n1724_n5888# 0.016694f
C1093 drain_right.n112 a_n1724_n5888# 0.031067f
C1094 drain_right.n113 a_n1724_n5888# 0.031067f
C1095 drain_right.n114 a_n1724_n5888# 0.016694f
C1096 drain_right.n115 a_n1724_n5888# 0.017185f
C1097 drain_right.n116 a_n1724_n5888# 0.017185f
C1098 drain_right.n117 a_n1724_n5888# 0.039459f
C1099 drain_right.n118 a_n1724_n5888# 0.039459f
C1100 drain_right.n119 a_n1724_n5888# 0.017676f
C1101 drain_right.n120 a_n1724_n5888# 0.016694f
C1102 drain_right.n121 a_n1724_n5888# 0.031067f
C1103 drain_right.n122 a_n1724_n5888# 0.031067f
C1104 drain_right.n123 a_n1724_n5888# 0.016694f
C1105 drain_right.n124 a_n1724_n5888# 0.017676f
C1106 drain_right.n125 a_n1724_n5888# 0.039459f
C1107 drain_right.n126 a_n1724_n5888# 0.039459f
C1108 drain_right.n127 a_n1724_n5888# 0.017676f
C1109 drain_right.n128 a_n1724_n5888# 0.016694f
C1110 drain_right.n129 a_n1724_n5888# 0.031067f
C1111 drain_right.n130 a_n1724_n5888# 0.031067f
C1112 drain_right.n131 a_n1724_n5888# 0.016694f
C1113 drain_right.n132 a_n1724_n5888# 0.017676f
C1114 drain_right.n133 a_n1724_n5888# 0.039459f
C1115 drain_right.n134 a_n1724_n5888# 0.083939f
C1116 drain_right.n135 a_n1724_n5888# 0.017676f
C1117 drain_right.n136 a_n1724_n5888# 0.016694f
C1118 drain_right.n137 a_n1724_n5888# 0.068415f
C1119 drain_right.n138 a_n1724_n5888# 0.069461f
C1120 drain_right.t7 a_n1724_n5888# 0.613751f
C1121 drain_right.t3 a_n1724_n5888# 0.613751f
C1122 drain_right.n139 a_n1724_n5888# 5.65638f
C1123 drain_right.n140 a_n1724_n5888# 0.465227f
C1124 drain_right.t12 a_n1724_n5888# 0.613751f
C1125 drain_right.t4 a_n1724_n5888# 0.613751f
C1126 drain_right.n141 a_n1724_n5888# 5.6599f
C1127 drain_right.t8 a_n1724_n5888# 0.613751f
C1128 drain_right.t11 a_n1724_n5888# 0.613751f
C1129 drain_right.n142 a_n1724_n5888# 5.65638f
C1130 drain_right.n143 a_n1724_n5888# 0.714315f
C1131 drain_right.n144 a_n1724_n5888# 2.43209f
C1132 drain_right.t13 a_n1724_n5888# 0.613751f
C1133 drain_right.t9 a_n1724_n5888# 0.613751f
C1134 drain_right.n145 a_n1724_n5888# 5.65989f
C1135 drain_right.t10 a_n1724_n5888# 0.613751f
C1136 drain_right.t0 a_n1724_n5888# 0.613751f
C1137 drain_right.n146 a_n1724_n5888# 5.65638f
C1138 drain_right.n147 a_n1724_n5888# 0.751687f
C1139 drain_right.t1 a_n1724_n5888# 0.613751f
C1140 drain_right.t6 a_n1724_n5888# 0.613751f
C1141 drain_right.n148 a_n1724_n5888# 5.65638f
C1142 drain_right.n149 a_n1724_n5888# 0.371339f
C1143 drain_right.n150 a_n1724_n5888# 0.042829f
C1144 drain_right.n151 a_n1724_n5888# 0.031067f
C1145 drain_right.n152 a_n1724_n5888# 0.016694f
C1146 drain_right.n153 a_n1724_n5888# 0.039459f
C1147 drain_right.n154 a_n1724_n5888# 0.017676f
C1148 drain_right.n155 a_n1724_n5888# 0.031067f
C1149 drain_right.n156 a_n1724_n5888# 0.016694f
C1150 drain_right.n157 a_n1724_n5888# 0.039459f
C1151 drain_right.n158 a_n1724_n5888# 0.017676f
C1152 drain_right.n159 a_n1724_n5888# 0.031067f
C1153 drain_right.n160 a_n1724_n5888# 0.016694f
C1154 drain_right.n161 a_n1724_n5888# 0.039459f
C1155 drain_right.n162 a_n1724_n5888# 0.017676f
C1156 drain_right.n163 a_n1724_n5888# 0.031067f
C1157 drain_right.n164 a_n1724_n5888# 0.016694f
C1158 drain_right.n165 a_n1724_n5888# 0.039459f
C1159 drain_right.n166 a_n1724_n5888# 0.039459f
C1160 drain_right.n167 a_n1724_n5888# 0.017676f
C1161 drain_right.n168 a_n1724_n5888# 0.031067f
C1162 drain_right.n169 a_n1724_n5888# 0.016694f
C1163 drain_right.n170 a_n1724_n5888# 0.039459f
C1164 drain_right.n171 a_n1724_n5888# 0.017676f
C1165 drain_right.n172 a_n1724_n5888# 0.031067f
C1166 drain_right.n173 a_n1724_n5888# 0.016694f
C1167 drain_right.n174 a_n1724_n5888# 0.039459f
C1168 drain_right.n175 a_n1724_n5888# 0.017676f
C1169 drain_right.n176 a_n1724_n5888# 0.031067f
C1170 drain_right.n177 a_n1724_n5888# 0.016694f
C1171 drain_right.n178 a_n1724_n5888# 0.039459f
C1172 drain_right.n179 a_n1724_n5888# 0.017676f
C1173 drain_right.n180 a_n1724_n5888# 0.031067f
C1174 drain_right.n181 a_n1724_n5888# 0.016694f
C1175 drain_right.n182 a_n1724_n5888# 0.039459f
C1176 drain_right.n183 a_n1724_n5888# 0.017676f
C1177 drain_right.n184 a_n1724_n5888# 0.031067f
C1178 drain_right.n185 a_n1724_n5888# 0.017185f
C1179 drain_right.n186 a_n1724_n5888# 0.039459f
C1180 drain_right.n187 a_n1724_n5888# 0.016694f
C1181 drain_right.n188 a_n1724_n5888# 0.017676f
C1182 drain_right.n189 a_n1724_n5888# 0.031067f
C1183 drain_right.n190 a_n1724_n5888# 0.016694f
C1184 drain_right.n191 a_n1724_n5888# 0.039459f
C1185 drain_right.n192 a_n1724_n5888# 0.017676f
C1186 drain_right.n193 a_n1724_n5888# 0.031067f
C1187 drain_right.n194 a_n1724_n5888# 0.016694f
C1188 drain_right.n195 a_n1724_n5888# 0.029594f
C1189 drain_right.n196 a_n1724_n5888# 0.027894f
C1190 drain_right.t5 a_n1724_n5888# 0.068818f
C1191 drain_right.n197 a_n1724_n5888# 0.379043f
C1192 drain_right.n198 a_n1724_n5888# 3.36364f
C1193 drain_right.n199 a_n1724_n5888# 0.016694f
C1194 drain_right.n200 a_n1724_n5888# 0.017676f
C1195 drain_right.n201 a_n1724_n5888# 0.039459f
C1196 drain_right.n202 a_n1724_n5888# 0.039459f
C1197 drain_right.n203 a_n1724_n5888# 0.017676f
C1198 drain_right.n204 a_n1724_n5888# 0.016694f
C1199 drain_right.n205 a_n1724_n5888# 0.031067f
C1200 drain_right.n206 a_n1724_n5888# 0.031067f
C1201 drain_right.n207 a_n1724_n5888# 0.016694f
C1202 drain_right.n208 a_n1724_n5888# 0.017676f
C1203 drain_right.n209 a_n1724_n5888# 0.039459f
C1204 drain_right.n210 a_n1724_n5888# 0.039459f
C1205 drain_right.n211 a_n1724_n5888# 0.017676f
C1206 drain_right.n212 a_n1724_n5888# 0.016694f
C1207 drain_right.n213 a_n1724_n5888# 0.031067f
C1208 drain_right.n214 a_n1724_n5888# 0.031067f
C1209 drain_right.n215 a_n1724_n5888# 0.016694f
C1210 drain_right.n216 a_n1724_n5888# 0.017676f
C1211 drain_right.n217 a_n1724_n5888# 0.039459f
C1212 drain_right.n218 a_n1724_n5888# 0.039459f
C1213 drain_right.n219 a_n1724_n5888# 0.039459f
C1214 drain_right.n220 a_n1724_n5888# 0.017185f
C1215 drain_right.n221 a_n1724_n5888# 0.016694f
C1216 drain_right.n222 a_n1724_n5888# 0.031067f
C1217 drain_right.n223 a_n1724_n5888# 0.031067f
C1218 drain_right.n224 a_n1724_n5888# 0.016694f
C1219 drain_right.n225 a_n1724_n5888# 0.017676f
C1220 drain_right.n226 a_n1724_n5888# 0.039459f
C1221 drain_right.n227 a_n1724_n5888# 0.039459f
C1222 drain_right.n228 a_n1724_n5888# 0.017676f
C1223 drain_right.n229 a_n1724_n5888# 0.016694f
C1224 drain_right.n230 a_n1724_n5888# 0.031067f
C1225 drain_right.n231 a_n1724_n5888# 0.031067f
C1226 drain_right.n232 a_n1724_n5888# 0.016694f
C1227 drain_right.n233 a_n1724_n5888# 0.017676f
C1228 drain_right.n234 a_n1724_n5888# 0.039459f
C1229 drain_right.n235 a_n1724_n5888# 0.039459f
C1230 drain_right.n236 a_n1724_n5888# 0.017676f
C1231 drain_right.n237 a_n1724_n5888# 0.016694f
C1232 drain_right.n238 a_n1724_n5888# 0.031067f
C1233 drain_right.n239 a_n1724_n5888# 0.031067f
C1234 drain_right.n240 a_n1724_n5888# 0.016694f
C1235 drain_right.n241 a_n1724_n5888# 0.017676f
C1236 drain_right.n242 a_n1724_n5888# 0.039459f
C1237 drain_right.n243 a_n1724_n5888# 0.039459f
C1238 drain_right.n244 a_n1724_n5888# 0.017676f
C1239 drain_right.n245 a_n1724_n5888# 0.016694f
C1240 drain_right.n246 a_n1724_n5888# 0.031067f
C1241 drain_right.n247 a_n1724_n5888# 0.031067f
C1242 drain_right.n248 a_n1724_n5888# 0.016694f
C1243 drain_right.n249 a_n1724_n5888# 0.017676f
C1244 drain_right.n250 a_n1724_n5888# 0.039459f
C1245 drain_right.n251 a_n1724_n5888# 0.039459f
C1246 drain_right.n252 a_n1724_n5888# 0.017676f
C1247 drain_right.n253 a_n1724_n5888# 0.016694f
C1248 drain_right.n254 a_n1724_n5888# 0.031067f
C1249 drain_right.n255 a_n1724_n5888# 0.031067f
C1250 drain_right.n256 a_n1724_n5888# 0.016694f
C1251 drain_right.n257 a_n1724_n5888# 0.017676f
C1252 drain_right.n258 a_n1724_n5888# 0.039459f
C1253 drain_right.n259 a_n1724_n5888# 0.039459f
C1254 drain_right.n260 a_n1724_n5888# 0.017676f
C1255 drain_right.n261 a_n1724_n5888# 0.016694f
C1256 drain_right.n262 a_n1724_n5888# 0.031067f
C1257 drain_right.n263 a_n1724_n5888# 0.031067f
C1258 drain_right.n264 a_n1724_n5888# 0.016694f
C1259 drain_right.n265 a_n1724_n5888# 0.017185f
C1260 drain_right.n266 a_n1724_n5888# 0.017185f
C1261 drain_right.n267 a_n1724_n5888# 0.039459f
C1262 drain_right.n268 a_n1724_n5888# 0.039459f
C1263 drain_right.n269 a_n1724_n5888# 0.017676f
C1264 drain_right.n270 a_n1724_n5888# 0.016694f
C1265 drain_right.n271 a_n1724_n5888# 0.031067f
C1266 drain_right.n272 a_n1724_n5888# 0.031067f
C1267 drain_right.n273 a_n1724_n5888# 0.016694f
C1268 drain_right.n274 a_n1724_n5888# 0.017676f
C1269 drain_right.n275 a_n1724_n5888# 0.039459f
C1270 drain_right.n276 a_n1724_n5888# 0.039459f
C1271 drain_right.n277 a_n1724_n5888# 0.017676f
C1272 drain_right.n278 a_n1724_n5888# 0.016694f
C1273 drain_right.n279 a_n1724_n5888# 0.031067f
C1274 drain_right.n280 a_n1724_n5888# 0.031067f
C1275 drain_right.n281 a_n1724_n5888# 0.016694f
C1276 drain_right.n282 a_n1724_n5888# 0.017676f
C1277 drain_right.n283 a_n1724_n5888# 0.039459f
C1278 drain_right.n284 a_n1724_n5888# 0.083939f
C1279 drain_right.n285 a_n1724_n5888# 0.017676f
C1280 drain_right.n286 a_n1724_n5888# 0.016694f
C1281 drain_right.n287 a_n1724_n5888# 0.068415f
C1282 drain_right.n288 a_n1724_n5888# 0.068188f
C1283 drain_right.n289 a_n1724_n5888# 0.371422f
C1284 minus.n0 a_n1724_n5888# 0.051699f
C1285 minus.t4 a_n1724_n5888# 1.10157f
C1286 minus.t0 a_n1724_n5888# 1.09099f
C1287 minus.t11 a_n1724_n5888# 1.09099f
C1288 minus.t7 a_n1724_n5888# 1.09099f
C1289 minus.n1 a_n1724_n5888# 0.414136f
C1290 minus.n2 a_n1724_n5888# 0.121803f
C1291 minus.t1 a_n1724_n5888# 1.09099f
C1292 minus.t12 a_n1724_n5888# 1.09099f
C1293 minus.t8 a_n1724_n5888# 1.10157f
C1294 minus.n3 a_n1724_n5888# 0.413837f
C1295 minus.n4 a_n1724_n5888# 0.396986f
C1296 minus.n5 a_n1724_n5888# 0.021294f
C1297 minus.n6 a_n1724_n5888# 0.396986f
C1298 minus.n7 a_n1724_n5888# 0.021294f
C1299 minus.n8 a_n1724_n5888# 0.051699f
C1300 minus.n9 a_n1724_n5888# 0.051699f
C1301 minus.n10 a_n1724_n5888# 0.051699f
C1302 minus.n11 a_n1724_n5888# 0.021294f
C1303 minus.n12 a_n1724_n5888# 0.396986f
C1304 minus.n13 a_n1724_n5888# 0.021294f
C1305 minus.n14 a_n1724_n5888# 0.396986f
C1306 minus.n15 a_n1724_n5888# 0.413755f
C1307 minus.n16 a_n1724_n5888# 2.57568f
C1308 minus.n17 a_n1724_n5888# 0.051699f
C1309 minus.t13 a_n1724_n5888# 1.09099f
C1310 minus.t6 a_n1724_n5888# 1.09099f
C1311 minus.t9 a_n1724_n5888# 1.09099f
C1312 minus.n18 a_n1724_n5888# 0.414136f
C1313 minus.n19 a_n1724_n5888# 0.121803f
C1314 minus.t2 a_n1724_n5888# 1.09099f
C1315 minus.t10 a_n1724_n5888# 1.09099f
C1316 minus.t3 a_n1724_n5888# 1.10157f
C1317 minus.n20 a_n1724_n5888# 0.413837f
C1318 minus.n21 a_n1724_n5888# 0.396986f
C1319 minus.n22 a_n1724_n5888# 0.021294f
C1320 minus.n23 a_n1724_n5888# 0.396986f
C1321 minus.n24 a_n1724_n5888# 0.021294f
C1322 minus.n25 a_n1724_n5888# 0.051699f
C1323 minus.n26 a_n1724_n5888# 0.051699f
C1324 minus.n27 a_n1724_n5888# 0.051699f
C1325 minus.n28 a_n1724_n5888# 0.021294f
C1326 minus.n29 a_n1724_n5888# 0.396986f
C1327 minus.n30 a_n1724_n5888# 0.021294f
C1328 minus.n31 a_n1724_n5888# 0.396986f
C1329 minus.t5 a_n1724_n5888# 1.10157f
C1330 minus.n32 a_n1724_n5888# 0.413755f
C1331 minus.n33 a_n1724_n5888# 0.342432f
C1332 minus.n34 a_n1724_n5888# 3.04491f
.ends

