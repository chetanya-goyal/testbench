* NGSPICE file created from diffpair492.ext - technology: sky130A

.subckt diffpair492 minus drain_right drain_left source plus
X0 drain_left.t5 plus.t0 source.t7 a_n1140_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X1 drain_left.t4 plus.t1 source.t8 a_n1140_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X2 a_n1140_n3888# a_n1140_n3888# a_n1140_n3888# a_n1140_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=46.8 ps=246.24 w=15 l=0.2
X3 drain_right.t5 minus.t0 source.t1 a_n1140_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X4 source.t6 plus.t2 drain_left.t3 a_n1140_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X5 source.t10 plus.t3 drain_left.t2 a_n1140_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X6 drain_right.t4 minus.t1 source.t2 a_n1140_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X7 source.t0 minus.t2 drain_right.t3 a_n1140_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X8 drain_right.t2 minus.t3 source.t5 a_n1140_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X9 a_n1140_n3888# a_n1140_n3888# a_n1140_n3888# a_n1140_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X10 drain_left.t1 plus.t4 source.t11 a_n1140_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=2.475 ps=15.33 w=15 l=0.2
X11 source.t4 minus.t4 drain_right.t1 a_n1140_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=2.475 ps=15.33 w=15 l=0.2
X12 a_n1140_n3888# a_n1140_n3888# a_n1140_n3888# a_n1140_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X13 drain_right.t0 minus.t5 source.t3 a_n1140_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
X14 a_n1140_n3888# a_n1140_n3888# a_n1140_n3888# a_n1140_n3888# sky130_fd_pr__nfet_01v8 ad=5.85 pd=30.78 as=0 ps=0 w=15 l=0.2
X15 drain_left.t0 plus.t5 source.t9 a_n1140_n3888# sky130_fd_pr__nfet_01v8 ad=2.475 pd=15.33 as=5.85 ps=30.78 w=15 l=0.2
R0 plus.n0 plus.t4 2005.05
R1 plus.n2 plus.t5 2005.05
R2 plus.n4 plus.t1 2005.05
R3 plus.n6 plus.t0 2005.05
R4 plus.n1 plus.t3 1964.15
R5 plus.n5 plus.t2 1964.15
R6 plus.n3 plus.n0 161.489
R7 plus.n7 plus.n4 161.489
R8 plus.n3 plus.n2 161.3
R9 plus.n7 plus.n6 161.3
R10 plus.n1 plus.n0 36.5157
R11 plus.n2 plus.n1 36.5157
R12 plus.n6 plus.n5 36.5157
R13 plus.n5 plus.n4 36.5157
R14 plus plus.n7 28.3949
R15 plus plus.n3 13.2183
R16 source.n3 source.t3 45.521
R17 source.n11 source.t2 45.5208
R18 source.n8 source.t8 45.5208
R19 source.n0 source.t9 45.5208
R20 source.n2 source.n1 44.201
R21 source.n5 source.n4 44.201
R22 source.n10 source.n9 44.2008
R23 source.n7 source.n6 44.2008
R24 source.n7 source.n5 24.4742
R25 source.n12 source.n0 18.526
R26 source.n12 source.n11 5.49188
R27 source.n9 source.t5 1.3205
R28 source.n9 source.t4 1.3205
R29 source.n6 source.t7 1.3205
R30 source.n6 source.t6 1.3205
R31 source.n1 source.t11 1.3205
R32 source.n1 source.t10 1.3205
R33 source.n4 source.t1 1.3205
R34 source.n4 source.t0 1.3205
R35 source.n3 source.n2 0.698776
R36 source.n10 source.n8 0.698776
R37 source.n5 source.n3 0.457397
R38 source.n2 source.n0 0.457397
R39 source.n8 source.n7 0.457397
R40 source.n11 source.n10 0.457397
R41 source source.n12 0.188
R42 drain_left.n3 drain_left.t1 62.6567
R43 drain_left.n1 drain_left.t5 62.4869
R44 drain_left.n1 drain_left.n0 60.9384
R45 drain_left.n3 drain_left.n2 60.8796
R46 drain_left drain_left.n1 30.8963
R47 drain_left drain_left.n3 6.11011
R48 drain_left.n0 drain_left.t3 1.3205
R49 drain_left.n0 drain_left.t4 1.3205
R50 drain_left.n2 drain_left.t2 1.3205
R51 drain_left.n2 drain_left.t0 1.3205
R52 minus.n2 minus.t0 2005.05
R53 minus.n0 minus.t5 2005.05
R54 minus.n6 minus.t1 2005.05
R55 minus.n4 minus.t3 2005.05
R56 minus.n1 minus.t2 1964.15
R57 minus.n5 minus.t4 1964.15
R58 minus.n3 minus.n0 161.489
R59 minus.n7 minus.n4 161.489
R60 minus.n3 minus.n2 161.3
R61 minus.n7 minus.n6 161.3
R62 minus.n2 minus.n1 36.5157
R63 minus.n1 minus.n0 36.5157
R64 minus.n5 minus.n4 36.5157
R65 minus.n6 minus.n5 36.5157
R66 minus.n8 minus.n3 35.6501
R67 minus.n8 minus.n7 6.438
R68 minus minus.n8 0.188
R69 drain_right.n1 drain_right.t2 62.4869
R70 drain_right.n3 drain_right.t5 62.1998
R71 drain_right.n3 drain_right.n2 61.3365
R72 drain_right.n1 drain_right.n0 60.9384
R73 drain_right drain_right.n1 30.343
R74 drain_right drain_right.n3 5.88166
R75 drain_right.n0 drain_right.t1 1.3205
R76 drain_right.n0 drain_right.t4 1.3205
R77 drain_right.n2 drain_right.t3 1.3205
R78 drain_right.n2 drain_right.t0 1.3205
C0 drain_left source 20.1038f
C1 drain_right plus 0.261837f
C2 minus drain_left 0.170484f
C3 source plus 1.99136f
C4 minus plus 5.13169f
C5 source drain_right 20.0882f
C6 minus drain_right 2.64234f
C7 minus source 1.97644f
C8 drain_left plus 2.74448f
C9 drain_left drain_right 0.536326f
C10 drain_right a_n1140_n3888# 7.438991f
C11 drain_left a_n1140_n3888# 7.61974f
C12 source a_n1140_n3888# 7.058882f
C13 minus a_n1140_n3888# 4.566799f
C14 plus a_n1140_n3888# 6.44839f
C15 drain_right.t2 a_n1140_n3888# 4.21043f
C16 drain_right.t1 a_n1140_n3888# 0.364779f
C17 drain_right.t4 a_n1140_n3888# 0.364779f
C18 drain_right.n0 a_n1140_n3888# 3.2975f
C19 drain_right.n1 a_n1140_n3888# 2.12547f
C20 drain_right.t3 a_n1140_n3888# 0.364779f
C21 drain_right.t0 a_n1140_n3888# 0.364779f
C22 drain_right.n2 a_n1140_n3888# 3.29982f
C23 drain_right.t5 a_n1140_n3888# 4.20869f
C24 drain_right.n3 a_n1140_n3888# 0.995657f
C25 minus.t5 a_n1140_n3888# 0.415602f
C26 minus.n0 a_n1140_n3888# 0.176572f
C27 minus.t0 a_n1140_n3888# 0.415602f
C28 minus.t2 a_n1140_n3888# 0.412283f
C29 minus.n1 a_n1140_n3888# 0.163366f
C30 minus.n2 a_n1140_n3888# 0.176506f
C31 minus.n3 a_n1140_n3888# 1.73528f
C32 minus.t3 a_n1140_n3888# 0.415602f
C33 minus.n4 a_n1140_n3888# 0.176572f
C34 minus.t4 a_n1140_n3888# 0.412283f
C35 minus.n5 a_n1140_n3888# 0.163366f
C36 minus.t1 a_n1140_n3888# 0.415602f
C37 minus.n6 a_n1140_n3888# 0.176506f
C38 minus.n7 a_n1140_n3888# 0.367794f
C39 minus.n8 a_n1140_n3888# 2.04507f
C40 drain_left.t5 a_n1140_n3888# 4.20667f
C41 drain_left.t3 a_n1140_n3888# 0.364454f
C42 drain_left.t4 a_n1140_n3888# 0.364454f
C43 drain_left.n0 a_n1140_n3888# 3.29455f
C44 drain_left.n1 a_n1140_n3888# 2.18839f
C45 drain_left.t1 a_n1140_n3888# 4.207799f
C46 drain_left.t2 a_n1140_n3888# 0.364454f
C47 drain_left.t0 a_n1140_n3888# 0.364454f
C48 drain_left.n2 a_n1140_n3888# 3.29423f
C49 drain_left.n3 a_n1140_n3888# 0.983893f
C50 source.t9 a_n1140_n3888# 3.78007f
C51 source.n0 a_n1140_n3888# 1.7381f
C52 source.t11 a_n1140_n3888# 0.337307f
C53 source.t10 a_n1140_n3888# 0.337307f
C54 source.n1 a_n1140_n3888# 2.96296f
C55 source.n2 a_n1140_n3888# 0.38622f
C56 source.t3 a_n1140_n3888# 3.78007f
C57 source.n3 a_n1140_n3888# 0.489035f
C58 source.t1 a_n1140_n3888# 0.337307f
C59 source.t0 a_n1140_n3888# 0.337307f
C60 source.n4 a_n1140_n3888# 2.96296f
C61 source.n5 a_n1140_n3888# 2.14723f
C62 source.t7 a_n1140_n3888# 0.337307f
C63 source.t6 a_n1140_n3888# 0.337307f
C64 source.n6 a_n1140_n3888# 2.96295f
C65 source.n7 a_n1140_n3888# 2.14724f
C66 source.t8 a_n1140_n3888# 3.78007f
C67 source.n8 a_n1140_n3888# 0.489039f
C68 source.t5 a_n1140_n3888# 0.337307f
C69 source.t4 a_n1140_n3888# 0.337307f
C70 source.n9 a_n1140_n3888# 2.96295f
C71 source.n10 a_n1140_n3888# 0.386224f
C72 source.t2 a_n1140_n3888# 3.78007f
C73 source.n11 a_n1140_n3888# 0.622392f
C74 source.n12 a_n1140_n3888# 2.07607f
C75 plus.t4 a_n1140_n3888# 0.426456f
C76 plus.n0 a_n1140_n3888# 0.181183f
C77 plus.t3 a_n1140_n3888# 0.423049f
C78 plus.n1 a_n1140_n3888# 0.167632f
C79 plus.t5 a_n1140_n3888# 0.426456f
C80 plus.n2 a_n1140_n3888# 0.181115f
C81 plus.n3 a_n1140_n3888# 0.682276f
C82 plus.t1 a_n1140_n3888# 0.426456f
C83 plus.n4 a_n1140_n3888# 0.181183f
C84 plus.t0 a_n1140_n3888# 0.426456f
C85 plus.t2 a_n1140_n3888# 0.423049f
C86 plus.n5 a_n1140_n3888# 0.167632f
C87 plus.n6 a_n1140_n3888# 0.181115f
C88 plus.n7 a_n1140_n3888# 1.46426f
.ends

