* NGSPICE file created from diffpair223.ext - technology: sky130A

.subckt diffpair223 minus drain_right drain_left source plus
X0 drain_right.t7 minus.t0 source.t15 a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X1 source.t14 minus.t1 drain_right.t6 a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X2 a_n1746_n1488# a_n1746_n1488# a_n1746_n1488# a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.7
X3 source.t7 plus.t0 drain_left.t7 a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X4 source.t12 minus.t2 drain_right.t5 a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X5 a_n1746_n1488# a_n1746_n1488# a_n1746_n1488# a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X6 source.t6 plus.t1 drain_left.t6 a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X7 drain_right.t4 minus.t3 source.t10 a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X8 source.t13 minus.t4 drain_right.t3 a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X9 drain_left.t5 plus.t2 source.t3 a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X10 source.t5 plus.t3 drain_left.t4 a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X11 drain_left.t3 plus.t4 source.t4 a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X12 drain_right.t2 minus.t5 source.t9 a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X13 drain_left.t2 plus.t5 source.t0 a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X14 drain_right.t1 minus.t6 source.t11 a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.7
X15 drain_left.t1 plus.t6 source.t2 a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.7
X16 a_n1746_n1488# a_n1746_n1488# a_n1746_n1488# a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X17 a_n1746_n1488# a_n1746_n1488# a_n1746_n1488# a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.7
X18 source.t1 plus.t7 drain_left.t0 a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
X19 source.t8 minus.t7 drain_right.t0 a_n1746_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.7
R0 minus.n3 minus.t6 181.583
R1 minus.n13 minus.t1 181.583
R2 minus.n9 minus.n8 161.3
R3 minus.n7 minus.n0 161.3
R4 minus.n6 minus.n5 161.3
R5 minus.n4 minus.n1 161.3
R6 minus.n19 minus.n18 161.3
R7 minus.n17 minus.n10 161.3
R8 minus.n16 minus.n15 161.3
R9 minus.n14 minus.n11 161.3
R10 minus.n2 minus.t2 159.405
R11 minus.n6 minus.t5 159.405
R12 minus.n8 minus.t7 159.405
R13 minus.n12 minus.t0 159.405
R14 minus.n16 minus.t4 159.405
R15 minus.n18 minus.t3 159.405
R16 minus.n4 minus.n3 44.862
R17 minus.n14 minus.n13 44.862
R18 minus.n20 minus.n9 29.0497
R19 minus.n8 minus.n7 28.4823
R20 minus.n18 minus.n17 28.4823
R21 minus.n6 minus.n1 24.1005
R22 minus.n2 minus.n1 24.1005
R23 minus.n12 minus.n11 24.1005
R24 minus.n16 minus.n11 24.1005
R25 minus.n7 minus.n6 19.7187
R26 minus.n17 minus.n16 19.7187
R27 minus.n3 minus.n2 19.7081
R28 minus.n13 minus.n12 19.7081
R29 minus.n20 minus.n19 6.63308
R30 minus.n9 minus.n0 0.189894
R31 minus.n5 minus.n0 0.189894
R32 minus.n5 minus.n4 0.189894
R33 minus.n15 minus.n14 0.189894
R34 minus.n15 minus.n10 0.189894
R35 minus.n19 minus.n10 0.189894
R36 minus minus.n20 0.188
R37 source.n0 source.t0 69.6943
R38 source.n3 source.t6 69.6943
R39 source.n4 source.t11 69.6943
R40 source.n7 source.t8 69.6943
R41 source.n15 source.t10 69.6942
R42 source.n12 source.t14 69.6942
R43 source.n11 source.t3 69.6942
R44 source.n8 source.t1 69.6942
R45 source.n2 source.n1 63.0943
R46 source.n6 source.n5 63.0943
R47 source.n14 source.n13 63.0942
R48 source.n10 source.n9 63.0942
R49 source.n8 source.n7 15.3575
R50 source.n16 source.n0 9.65058
R51 source.n13 source.t15 6.6005
R52 source.n13 source.t13 6.6005
R53 source.n9 source.t4 6.6005
R54 source.n9 source.t5 6.6005
R55 source.n1 source.t2 6.6005
R56 source.n1 source.t7 6.6005
R57 source.n5 source.t9 6.6005
R58 source.n5 source.t12 6.6005
R59 source.n16 source.n15 5.7074
R60 source.n7 source.n6 0.888431
R61 source.n6 source.n4 0.888431
R62 source.n3 source.n2 0.888431
R63 source.n2 source.n0 0.888431
R64 source.n10 source.n8 0.888431
R65 source.n11 source.n10 0.888431
R66 source.n14 source.n12 0.888431
R67 source.n15 source.n14 0.888431
R68 source.n4 source.n3 0.470328
R69 source.n12 source.n11 0.470328
R70 source source.n16 0.188
R71 drain_right.n5 drain_right.n3 80.661
R72 drain_right.n2 drain_right.n1 80.1616
R73 drain_right.n2 drain_right.n0 80.1616
R74 drain_right.n5 drain_right.n4 79.7731
R75 drain_right drain_right.n2 23.1034
R76 drain_right.n1 drain_right.t3 6.6005
R77 drain_right.n1 drain_right.t4 6.6005
R78 drain_right.n0 drain_right.t6 6.6005
R79 drain_right.n0 drain_right.t7 6.6005
R80 drain_right.n3 drain_right.t5 6.6005
R81 drain_right.n3 drain_right.t1 6.6005
R82 drain_right.n4 drain_right.t0 6.6005
R83 drain_right.n4 drain_right.t2 6.6005
R84 drain_right drain_right.n5 6.54115
R85 plus.n3 plus.t1 181.583
R86 plus.n13 plus.t2 181.583
R87 plus.n5 plus.n4 161.3
R88 plus.n6 plus.n1 161.3
R89 plus.n7 plus.n0 161.3
R90 plus.n9 plus.n8 161.3
R91 plus.n15 plus.n14 161.3
R92 plus.n16 plus.n11 161.3
R93 plus.n17 plus.n10 161.3
R94 plus.n19 plus.n18 161.3
R95 plus.n8 plus.t5 159.405
R96 plus.n6 plus.t0 159.405
R97 plus.n2 plus.t6 159.405
R98 plus.n18 plus.t7 159.405
R99 plus.n16 plus.t4 159.405
R100 plus.n12 plus.t3 159.405
R101 plus.n4 plus.n3 44.862
R102 plus.n14 plus.n13 44.862
R103 plus.n8 plus.n7 28.4823
R104 plus.n18 plus.n17 28.4823
R105 plus plus.n19 26.3399
R106 plus.n5 plus.n2 24.1005
R107 plus.n6 plus.n5 24.1005
R108 plus.n16 plus.n15 24.1005
R109 plus.n15 plus.n12 24.1005
R110 plus.n7 plus.n6 19.7187
R111 plus.n17 plus.n16 19.7187
R112 plus.n3 plus.n2 19.7081
R113 plus.n13 plus.n12 19.7081
R114 plus plus.n9 8.86792
R115 plus.n4 plus.n1 0.189894
R116 plus.n1 plus.n0 0.189894
R117 plus.n9 plus.n0 0.189894
R118 plus.n19 plus.n10 0.189894
R119 plus.n11 plus.n10 0.189894
R120 plus.n14 plus.n11 0.189894
R121 drain_left.n5 drain_left.n3 80.661
R122 drain_left.n2 drain_left.n1 80.1616
R123 drain_left.n2 drain_left.n0 80.1616
R124 drain_left.n5 drain_left.n4 79.7731
R125 drain_left drain_left.n2 23.6567
R126 drain_left.n1 drain_left.t4 6.6005
R127 drain_left.n1 drain_left.t5 6.6005
R128 drain_left.n0 drain_left.t0 6.6005
R129 drain_left.n0 drain_left.t3 6.6005
R130 drain_left.n4 drain_left.t7 6.6005
R131 drain_left.n4 drain_left.t2 6.6005
R132 drain_left.n3 drain_left.t6 6.6005
R133 drain_left.n3 drain_left.t1 6.6005
R134 drain_left drain_left.n5 6.54115
C0 source minus 1.88344f
C1 drain_left source 4.43614f
C2 drain_right source 4.43791f
C3 drain_left minus 0.17601f
C4 source plus 1.89743f
C5 drain_right minus 1.68047f
C6 drain_left drain_right 0.821811f
C7 plus minus 3.65923f
C8 drain_left plus 1.84929f
C9 drain_right plus 0.328414f
C10 drain_right a_n1746_n1488# 3.43584f
C11 drain_left a_n1746_n1488# 3.65213f
C12 source a_n1746_n1488# 3.655123f
C13 minus a_n1746_n1488# 6.027393f
C14 plus a_n1746_n1488# 6.560029f
C15 drain_left.t0 a_n1746_n1488# 0.043638f
C16 drain_left.t3 a_n1746_n1488# 0.043638f
C17 drain_left.n0 a_n1746_n1488# 0.315837f
C18 drain_left.t4 a_n1746_n1488# 0.043638f
C19 drain_left.t5 a_n1746_n1488# 0.043638f
C20 drain_left.n1 a_n1746_n1488# 0.315837f
C21 drain_left.n2 a_n1746_n1488# 1.01694f
C22 drain_left.t6 a_n1746_n1488# 0.043638f
C23 drain_left.t1 a_n1746_n1488# 0.043638f
C24 drain_left.n3 a_n1746_n1488# 0.317579f
C25 drain_left.t7 a_n1746_n1488# 0.043638f
C26 drain_left.t2 a_n1746_n1488# 0.043638f
C27 drain_left.n4 a_n1746_n1488# 0.314716f
C28 drain_left.n5 a_n1746_n1488# 0.672721f
C29 plus.n0 a_n1746_n1488# 0.024058f
C30 plus.t5 a_n1746_n1488# 0.151494f
C31 plus.t0 a_n1746_n1488# 0.151494f
C32 plus.n1 a_n1746_n1488# 0.024058f
C33 plus.t6 a_n1746_n1488# 0.151494f
C34 plus.n2 a_n1746_n1488# 0.090411f
C35 plus.t1 a_n1746_n1488# 0.162256f
C36 plus.n3 a_n1746_n1488# 0.079686f
C37 plus.n4 a_n1746_n1488# 0.100043f
C38 plus.n5 a_n1746_n1488# 0.005459f
C39 plus.n6 a_n1746_n1488# 0.088234f
C40 plus.n7 a_n1746_n1488# 0.005459f
C41 plus.n8 a_n1746_n1488# 0.086676f
C42 plus.n9 a_n1746_n1488# 0.187604f
C43 plus.n10 a_n1746_n1488# 0.024058f
C44 plus.t7 a_n1746_n1488# 0.151494f
C45 plus.n11 a_n1746_n1488# 0.024058f
C46 plus.t4 a_n1746_n1488# 0.151494f
C47 plus.t3 a_n1746_n1488# 0.151494f
C48 plus.n12 a_n1746_n1488# 0.090411f
C49 plus.t2 a_n1746_n1488# 0.162256f
C50 plus.n13 a_n1746_n1488# 0.079686f
C51 plus.n14 a_n1746_n1488# 0.100043f
C52 plus.n15 a_n1746_n1488# 0.005459f
C53 plus.n16 a_n1746_n1488# 0.088234f
C54 plus.n17 a_n1746_n1488# 0.005459f
C55 plus.n18 a_n1746_n1488# 0.086676f
C56 plus.n19 a_n1746_n1488# 0.560574f
C57 drain_right.t6 a_n1746_n1488# 0.044364f
C58 drain_right.t7 a_n1746_n1488# 0.044364f
C59 drain_right.n0 a_n1746_n1488# 0.321092f
C60 drain_right.t3 a_n1746_n1488# 0.044364f
C61 drain_right.t4 a_n1746_n1488# 0.044364f
C62 drain_right.n1 a_n1746_n1488# 0.321092f
C63 drain_right.n2 a_n1746_n1488# 0.996727f
C64 drain_right.t5 a_n1746_n1488# 0.044364f
C65 drain_right.t1 a_n1746_n1488# 0.044364f
C66 drain_right.n3 a_n1746_n1488# 0.322863f
C67 drain_right.t0 a_n1746_n1488# 0.044364f
C68 drain_right.t2 a_n1746_n1488# 0.044364f
C69 drain_right.n4 a_n1746_n1488# 0.319952f
C70 drain_right.n5 a_n1746_n1488# 0.683913f
C71 source.t0 a_n1746_n1488# 0.336828f
C72 source.n0 a_n1746_n1488# 0.492941f
C73 source.t2 a_n1746_n1488# 0.040563f
C74 source.t7 a_n1746_n1488# 0.040563f
C75 source.n1 a_n1746_n1488# 0.257193f
C76 source.n2 a_n1746_n1488# 0.246961f
C77 source.t6 a_n1746_n1488# 0.336828f
C78 source.n3 a_n1746_n1488# 0.2549f
C79 source.t11 a_n1746_n1488# 0.336828f
C80 source.n4 a_n1746_n1488# 0.2549f
C81 source.t9 a_n1746_n1488# 0.040563f
C82 source.t12 a_n1746_n1488# 0.040563f
C83 source.n5 a_n1746_n1488# 0.257193f
C84 source.n6 a_n1746_n1488# 0.246961f
C85 source.t8 a_n1746_n1488# 0.336828f
C86 source.n7 a_n1746_n1488# 0.67592f
C87 source.t1 a_n1746_n1488# 0.336827f
C88 source.n8 a_n1746_n1488# 0.675922f
C89 source.t4 a_n1746_n1488# 0.040563f
C90 source.t5 a_n1746_n1488# 0.040563f
C91 source.n9 a_n1746_n1488# 0.257191f
C92 source.n10 a_n1746_n1488# 0.246962f
C93 source.t3 a_n1746_n1488# 0.336827f
C94 source.n11 a_n1746_n1488# 0.254902f
C95 source.t14 a_n1746_n1488# 0.336827f
C96 source.n12 a_n1746_n1488# 0.254902f
C97 source.t15 a_n1746_n1488# 0.040563f
C98 source.t13 a_n1746_n1488# 0.040563f
C99 source.n13 a_n1746_n1488# 0.257191f
C100 source.n14 a_n1746_n1488# 0.246962f
C101 source.t10 a_n1746_n1488# 0.336827f
C102 source.n15 a_n1746_n1488# 0.366513f
C103 source.n16 a_n1746_n1488# 0.504559f
C104 minus.n0 a_n1746_n1488# 0.023745f
C105 minus.n1 a_n1746_n1488# 0.005388f
C106 minus.t5 a_n1746_n1488# 0.149528f
C107 minus.t6 a_n1746_n1488# 0.16015f
C108 minus.t2 a_n1746_n1488# 0.149528f
C109 minus.n2 a_n1746_n1488# 0.089237f
C110 minus.n3 a_n1746_n1488# 0.078652f
C111 minus.n4 a_n1746_n1488# 0.098745f
C112 minus.n5 a_n1746_n1488# 0.023745f
C113 minus.n6 a_n1746_n1488# 0.087089f
C114 minus.n7 a_n1746_n1488# 0.005388f
C115 minus.t7 a_n1746_n1488# 0.149528f
C116 minus.n8 a_n1746_n1488# 0.085551f
C117 minus.n9 a_n1746_n1488# 0.587452f
C118 minus.n10 a_n1746_n1488# 0.023745f
C119 minus.n11 a_n1746_n1488# 0.005388f
C120 minus.t1 a_n1746_n1488# 0.16015f
C121 minus.t0 a_n1746_n1488# 0.149528f
C122 minus.n12 a_n1746_n1488# 0.089237f
C123 minus.n13 a_n1746_n1488# 0.078652f
C124 minus.n14 a_n1746_n1488# 0.098745f
C125 minus.n15 a_n1746_n1488# 0.023745f
C126 minus.t4 a_n1746_n1488# 0.149528f
C127 minus.n16 a_n1746_n1488# 0.087089f
C128 minus.n17 a_n1746_n1488# 0.005388f
C129 minus.t3 a_n1746_n1488# 0.149528f
C130 minus.n18 a_n1746_n1488# 0.085551f
C131 minus.n19 a_n1746_n1488# 0.162639f
C132 minus.n20 a_n1746_n1488# 0.721766f
.ends

