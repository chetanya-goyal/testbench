* NGSPICE file created from diffpair378.ext - technology: sky130A

.subckt diffpair378 minus drain_right drain_left source plus
X0 drain_left.t19 plus.t0 source.t25 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X1 drain_left.t18 plus.t1 source.t38 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X2 source.t29 plus.t2 drain_left.t17 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X3 drain_left.t16 plus.t3 source.t31 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X4 source.t12 minus.t0 drain_right.t19 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X5 source.t21 plus.t4 drain_left.t15 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X6 drain_right.t18 minus.t1 source.t0 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X7 source.t15 minus.t2 drain_right.t17 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X8 drain_left.t14 plus.t5 source.t35 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X9 source.t2 minus.t3 drain_right.t16 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X10 source.t9 minus.t4 drain_right.t15 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X11 drain_right.t14 minus.t5 source.t3 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X12 drain_right.t13 minus.t6 source.t5 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X13 source.t24 plus.t6 drain_left.t13 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X14 source.t16 minus.t7 drain_right.t12 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X15 a_n2762_n2688# a_n2762_n2688# a_n2762_n2688# a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.6
X16 a_n2762_n2688# a_n2762_n2688# a_n2762_n2688# a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X17 source.t6 minus.t8 drain_right.t11 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X18 drain_right.t10 minus.t9 source.t10 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X19 source.t13 minus.t10 drain_right.t9 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X20 source.t37 plus.t7 drain_left.t12 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X21 drain_left.t11 plus.t8 source.t26 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X22 drain_left.t10 plus.t9 source.t23 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X23 source.t4 minus.t11 drain_right.t8 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X24 source.t20 plus.t10 drain_left.t9 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X25 drain_right.t7 minus.t12 source.t1 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X26 a_n2762_n2688# a_n2762_n2688# a_n2762_n2688# a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X27 drain_left.t8 plus.t11 source.t27 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X28 source.t17 minus.t13 drain_right.t6 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X29 source.t39 plus.t12 drain_left.t7 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X30 drain_right.t5 minus.t14 source.t11 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X31 drain_right.t4 minus.t15 source.t8 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X32 drain_left.t6 plus.t13 source.t36 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X33 source.t30 plus.t14 drain_left.t5 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.6
X34 drain_right.t3 minus.t16 source.t18 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X35 drain_left.t4 plus.t15 source.t22 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.6
X36 a_n2762_n2688# a_n2762_n2688# a_n2762_n2688# a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.6
X37 source.t28 plus.t16 drain_left.t3 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X38 source.t32 plus.t17 drain_left.t2 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X39 drain_right.t2 minus.t17 source.t19 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X40 drain_left.t1 plus.t18 source.t33 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X41 source.t7 minus.t18 drain_right.t1 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X42 drain_right.t0 minus.t19 source.t14 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
X43 source.t34 plus.t19 drain_left.t0 a_n2762_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.6
R0 plus.n8 plus.t14 453.793
R1 plus.n36 plus.t15 453.793
R2 plus.n26 plus.t0 426.973
R3 plus.n25 plus.t2 426.973
R4 plus.n24 plus.t3 426.973
R5 plus.n2 plus.t4 426.973
R6 plus.n18 plus.t5 426.973
R7 plus.n4 plus.t7 426.973
R8 plus.n12 plus.t11 426.973
R9 plus.n6 plus.t12 426.973
R10 plus.n7 plus.t13 426.973
R11 plus.n54 plus.t10 426.973
R12 plus.n53 plus.t1 426.973
R13 plus.n52 plus.t17 426.973
R14 plus.n30 plus.t9 426.973
R15 plus.n46 plus.t19 426.973
R16 plus.n32 plus.t18 426.973
R17 plus.n40 plus.t16 426.973
R18 plus.n34 plus.t8 426.973
R19 plus.n35 plus.t6 426.973
R20 plus.n9 plus.n6 161.3
R21 plus.n11 plus.n10 161.3
R22 plus.n12 plus.n5 161.3
R23 plus.n14 plus.n13 161.3
R24 plus.n15 plus.n4 161.3
R25 plus.n17 plus.n16 161.3
R26 plus.n18 plus.n3 161.3
R27 plus.n20 plus.n19 161.3
R28 plus.n21 plus.n2 161.3
R29 plus.n23 plus.n22 161.3
R30 plus.n24 plus.n1 161.3
R31 plus.n27 plus.n26 161.3
R32 plus.n37 plus.n34 161.3
R33 plus.n39 plus.n38 161.3
R34 plus.n40 plus.n33 161.3
R35 plus.n42 plus.n41 161.3
R36 plus.n43 plus.n32 161.3
R37 plus.n45 plus.n44 161.3
R38 plus.n46 plus.n31 161.3
R39 plus.n48 plus.n47 161.3
R40 plus.n49 plus.n30 161.3
R41 plus.n51 plus.n50 161.3
R42 plus.n52 plus.n29 161.3
R43 plus.n55 plus.n54 161.3
R44 plus.n25 plus.n0 80.6037
R45 plus.n53 plus.n28 80.6037
R46 plus.n26 plus.n25 48.2005
R47 plus.n25 plus.n24 48.2005
R48 plus.n7 plus.n6 48.2005
R49 plus.n54 plus.n53 48.2005
R50 plus.n53 plus.n52 48.2005
R51 plus.n35 plus.n34 48.2005
R52 plus.n9 plus.n8 45.1367
R53 plus.n37 plus.n36 45.1367
R54 plus.n23 plus.n2 44.549
R55 plus.n12 plus.n11 44.549
R56 plus.n51 plus.n30 44.549
R57 plus.n40 plus.n39 44.549
R58 plus.n19 plus.n18 34.3247
R59 plus.n13 plus.n4 34.3247
R60 plus.n47 plus.n46 34.3247
R61 plus.n41 plus.n32 34.3247
R62 plus plus.n55 32.4574
R63 plus.n17 plus.n4 24.1005
R64 plus.n18 plus.n17 24.1005
R65 plus.n46 plus.n45 24.1005
R66 plus.n45 plus.n32 24.1005
R67 plus.n19 plus.n2 13.8763
R68 plus.n13 plus.n12 13.8763
R69 plus.n47 plus.n30 13.8763
R70 plus.n41 plus.n40 13.8763
R71 plus.n8 plus.n7 13.3799
R72 plus.n36 plus.n35 13.3799
R73 plus plus.n27 11.1369
R74 plus.n24 plus.n23 3.65202
R75 plus.n11 plus.n6 3.65202
R76 plus.n52 plus.n51 3.65202
R77 plus.n39 plus.n34 3.65202
R78 plus.n1 plus.n0 0.285035
R79 plus.n27 plus.n0 0.285035
R80 plus.n55 plus.n28 0.285035
R81 plus.n29 plus.n28 0.285035
R82 plus.n10 plus.n9 0.189894
R83 plus.n10 plus.n5 0.189894
R84 plus.n14 plus.n5 0.189894
R85 plus.n15 plus.n14 0.189894
R86 plus.n16 plus.n15 0.189894
R87 plus.n16 plus.n3 0.189894
R88 plus.n20 plus.n3 0.189894
R89 plus.n21 plus.n20 0.189894
R90 plus.n22 plus.n21 0.189894
R91 plus.n22 plus.n1 0.189894
R92 plus.n50 plus.n29 0.189894
R93 plus.n50 plus.n49 0.189894
R94 plus.n49 plus.n48 0.189894
R95 plus.n48 plus.n31 0.189894
R96 plus.n44 plus.n31 0.189894
R97 plus.n44 plus.n43 0.189894
R98 plus.n43 plus.n42 0.189894
R99 plus.n42 plus.n33 0.189894
R100 plus.n38 plus.n33 0.189894
R101 plus.n38 plus.n37 0.189894
R102 source.n9 source.t30 51.0588
R103 source.n10 source.t11 51.0588
R104 source.n19 source.t12 51.0588
R105 source.n39 source.t10 51.0586
R106 source.n30 source.t13 51.0586
R107 source.n29 source.t22 51.0586
R108 source.n20 source.t20 51.0586
R109 source.n0 source.t25 51.0586
R110 source.n2 source.n1 48.8588
R111 source.n4 source.n3 48.8588
R112 source.n6 source.n5 48.8588
R113 source.n8 source.n7 48.8588
R114 source.n12 source.n11 48.8588
R115 source.n14 source.n13 48.8588
R116 source.n16 source.n15 48.8588
R117 source.n18 source.n17 48.8588
R118 source.n38 source.n37 48.8586
R119 source.n36 source.n35 48.8586
R120 source.n34 source.n33 48.8586
R121 source.n32 source.n31 48.8586
R122 source.n28 source.n27 48.8586
R123 source.n26 source.n25 48.8586
R124 source.n24 source.n23 48.8586
R125 source.n22 source.n21 48.8586
R126 source.n20 source.n19 19.8167
R127 source.n40 source.n0 14.1529
R128 source.n40 source.n39 5.66429
R129 source.n37 source.t8 2.2005
R130 source.n37 source.t15 2.2005
R131 source.n35 source.t19 2.2005
R132 source.n35 source.t6 2.2005
R133 source.n33 source.t18 2.2005
R134 source.n33 source.t7 2.2005
R135 source.n31 source.t14 2.2005
R136 source.n31 source.t9 2.2005
R137 source.n27 source.t26 2.2005
R138 source.n27 source.t24 2.2005
R139 source.n25 source.t33 2.2005
R140 source.n25 source.t28 2.2005
R141 source.n23 source.t23 2.2005
R142 source.n23 source.t34 2.2005
R143 source.n21 source.t38 2.2005
R144 source.n21 source.t32 2.2005
R145 source.n1 source.t31 2.2005
R146 source.n1 source.t29 2.2005
R147 source.n3 source.t35 2.2005
R148 source.n3 source.t21 2.2005
R149 source.n5 source.t27 2.2005
R150 source.n5 source.t37 2.2005
R151 source.n7 source.t36 2.2005
R152 source.n7 source.t39 2.2005
R153 source.n11 source.t1 2.2005
R154 source.n11 source.t17 2.2005
R155 source.n13 source.t3 2.2005
R156 source.n13 source.t4 2.2005
R157 source.n15 source.t5 2.2005
R158 source.n15 source.t16 2.2005
R159 source.n17 source.t0 2.2005
R160 source.n17 source.t2 2.2005
R161 source.n19 source.n18 0.802224
R162 source.n18 source.n16 0.802224
R163 source.n16 source.n14 0.802224
R164 source.n14 source.n12 0.802224
R165 source.n12 source.n10 0.802224
R166 source.n9 source.n8 0.802224
R167 source.n8 source.n6 0.802224
R168 source.n6 source.n4 0.802224
R169 source.n4 source.n2 0.802224
R170 source.n2 source.n0 0.802224
R171 source.n22 source.n20 0.802224
R172 source.n24 source.n22 0.802224
R173 source.n26 source.n24 0.802224
R174 source.n28 source.n26 0.802224
R175 source.n29 source.n28 0.802224
R176 source.n32 source.n30 0.802224
R177 source.n34 source.n32 0.802224
R178 source.n36 source.n34 0.802224
R179 source.n38 source.n36 0.802224
R180 source.n39 source.n38 0.802224
R181 source.n10 source.n9 0.470328
R182 source.n30 source.n29 0.470328
R183 source source.n40 0.188
R184 drain_left.n10 drain_left.n8 66.3393
R185 drain_left.n6 drain_left.n4 66.3391
R186 drain_left.n2 drain_left.n0 66.3391
R187 drain_left.n14 drain_left.n13 65.5376
R188 drain_left.n12 drain_left.n11 65.5376
R189 drain_left.n10 drain_left.n9 65.5376
R190 drain_left.n16 drain_left.n15 65.5374
R191 drain_left.n7 drain_left.n3 65.5373
R192 drain_left.n6 drain_left.n5 65.5373
R193 drain_left.n2 drain_left.n1 65.5373
R194 drain_left drain_left.n7 31.5081
R195 drain_left drain_left.n16 6.45494
R196 drain_left.n3 drain_left.t0 2.2005
R197 drain_left.n3 drain_left.t1 2.2005
R198 drain_left.n4 drain_left.t13 2.2005
R199 drain_left.n4 drain_left.t4 2.2005
R200 drain_left.n5 drain_left.t3 2.2005
R201 drain_left.n5 drain_left.t11 2.2005
R202 drain_left.n1 drain_left.t2 2.2005
R203 drain_left.n1 drain_left.t10 2.2005
R204 drain_left.n0 drain_left.t9 2.2005
R205 drain_left.n0 drain_left.t18 2.2005
R206 drain_left.n15 drain_left.t17 2.2005
R207 drain_left.n15 drain_left.t19 2.2005
R208 drain_left.n13 drain_left.t15 2.2005
R209 drain_left.n13 drain_left.t16 2.2005
R210 drain_left.n11 drain_left.t12 2.2005
R211 drain_left.n11 drain_left.t14 2.2005
R212 drain_left.n9 drain_left.t7 2.2005
R213 drain_left.n9 drain_left.t8 2.2005
R214 drain_left.n8 drain_left.t5 2.2005
R215 drain_left.n8 drain_left.t6 2.2005
R216 drain_left.n12 drain_left.n10 0.802224
R217 drain_left.n14 drain_left.n12 0.802224
R218 drain_left.n16 drain_left.n14 0.802224
R219 drain_left.n7 drain_left.n6 0.746878
R220 drain_left.n7 drain_left.n2 0.746878
R221 minus.n6 minus.t14 453.793
R222 minus.n34 minus.t10 453.793
R223 minus.n7 minus.t13 426.973
R224 minus.n8 minus.t12 426.973
R225 minus.n12 minus.t11 426.973
R226 minus.n14 minus.t5 426.973
R227 minus.n18 minus.t7 426.973
R228 minus.n20 minus.t6 426.973
R229 minus.n24 minus.t3 426.973
R230 minus.n25 minus.t1 426.973
R231 minus.n26 minus.t0 426.973
R232 minus.n35 minus.t19 426.973
R233 minus.n36 minus.t4 426.973
R234 minus.n40 minus.t16 426.973
R235 minus.n42 minus.t18 426.973
R236 minus.n46 minus.t17 426.973
R237 minus.n48 minus.t8 426.973
R238 minus.n52 minus.t15 426.973
R239 minus.n53 minus.t2 426.973
R240 minus.n54 minus.t9 426.973
R241 minus.n27 minus.n26 161.3
R242 minus.n24 minus.n23 161.3
R243 minus.n22 minus.n1 161.3
R244 minus.n21 minus.n20 161.3
R245 minus.n19 minus.n2 161.3
R246 minus.n18 minus.n17 161.3
R247 minus.n16 minus.n3 161.3
R248 minus.n15 minus.n14 161.3
R249 minus.n13 minus.n4 161.3
R250 minus.n12 minus.n11 161.3
R251 minus.n10 minus.n5 161.3
R252 minus.n9 minus.n8 161.3
R253 minus.n55 minus.n54 161.3
R254 minus.n52 minus.n51 161.3
R255 minus.n50 minus.n29 161.3
R256 minus.n49 minus.n48 161.3
R257 minus.n47 minus.n30 161.3
R258 minus.n46 minus.n45 161.3
R259 minus.n44 minus.n31 161.3
R260 minus.n43 minus.n42 161.3
R261 minus.n41 minus.n32 161.3
R262 minus.n40 minus.n39 161.3
R263 minus.n38 minus.n33 161.3
R264 minus.n37 minus.n36 161.3
R265 minus.n25 minus.n0 80.6037
R266 minus.n53 minus.n28 80.6037
R267 minus.n8 minus.n7 48.2005
R268 minus.n25 minus.n24 48.2005
R269 minus.n26 minus.n25 48.2005
R270 minus.n36 minus.n35 48.2005
R271 minus.n53 minus.n52 48.2005
R272 minus.n54 minus.n53 48.2005
R273 minus.n9 minus.n6 45.1367
R274 minus.n37 minus.n34 45.1367
R275 minus.n12 minus.n5 44.549
R276 minus.n20 minus.n1 44.549
R277 minus.n40 minus.n33 44.549
R278 minus.n48 minus.n29 44.549
R279 minus.n56 minus.n27 37.4399
R280 minus.n14 minus.n13 34.3247
R281 minus.n19 minus.n18 34.3247
R282 minus.n42 minus.n41 34.3247
R283 minus.n47 minus.n46 34.3247
R284 minus.n18 minus.n3 24.1005
R285 minus.n14 minus.n3 24.1005
R286 minus.n42 minus.n31 24.1005
R287 minus.n46 minus.n31 24.1005
R288 minus.n13 minus.n12 13.8763
R289 minus.n20 minus.n19 13.8763
R290 minus.n41 minus.n40 13.8763
R291 minus.n48 minus.n47 13.8763
R292 minus.n7 minus.n6 13.3799
R293 minus.n35 minus.n34 13.3799
R294 minus.n56 minus.n55 6.62929
R295 minus.n8 minus.n5 3.65202
R296 minus.n24 minus.n1 3.65202
R297 minus.n36 minus.n33 3.65202
R298 minus.n52 minus.n29 3.65202
R299 minus.n27 minus.n0 0.285035
R300 minus.n23 minus.n0 0.285035
R301 minus.n51 minus.n28 0.285035
R302 minus.n55 minus.n28 0.285035
R303 minus.n23 minus.n22 0.189894
R304 minus.n22 minus.n21 0.189894
R305 minus.n21 minus.n2 0.189894
R306 minus.n17 minus.n2 0.189894
R307 minus.n17 minus.n16 0.189894
R308 minus.n16 minus.n15 0.189894
R309 minus.n15 minus.n4 0.189894
R310 minus.n11 minus.n4 0.189894
R311 minus.n11 minus.n10 0.189894
R312 minus.n10 minus.n9 0.189894
R313 minus.n38 minus.n37 0.189894
R314 minus.n39 minus.n38 0.189894
R315 minus.n39 minus.n32 0.189894
R316 minus.n43 minus.n32 0.189894
R317 minus.n44 minus.n43 0.189894
R318 minus.n45 minus.n44 0.189894
R319 minus.n45 minus.n30 0.189894
R320 minus.n49 minus.n30 0.189894
R321 minus.n50 minus.n49 0.189894
R322 minus.n51 minus.n50 0.189894
R323 minus minus.n56 0.188
R324 drain_right.n10 drain_right.n8 66.3391
R325 drain_right.n6 drain_right.n4 66.3391
R326 drain_right.n2 drain_right.n0 66.3391
R327 drain_right.n10 drain_right.n9 65.5376
R328 drain_right.n12 drain_right.n11 65.5376
R329 drain_right.n14 drain_right.n13 65.5376
R330 drain_right.n16 drain_right.n15 65.5376
R331 drain_right.n7 drain_right.n3 65.5373
R332 drain_right.n6 drain_right.n5 65.5373
R333 drain_right.n2 drain_right.n1 65.5373
R334 drain_right drain_right.n7 30.9549
R335 drain_right drain_right.n16 6.45494
R336 drain_right.n3 drain_right.t1 2.2005
R337 drain_right.n3 drain_right.t2 2.2005
R338 drain_right.n4 drain_right.t17 2.2005
R339 drain_right.n4 drain_right.t10 2.2005
R340 drain_right.n5 drain_right.t11 2.2005
R341 drain_right.n5 drain_right.t4 2.2005
R342 drain_right.n1 drain_right.t15 2.2005
R343 drain_right.n1 drain_right.t3 2.2005
R344 drain_right.n0 drain_right.t9 2.2005
R345 drain_right.n0 drain_right.t0 2.2005
R346 drain_right.n8 drain_right.t6 2.2005
R347 drain_right.n8 drain_right.t5 2.2005
R348 drain_right.n9 drain_right.t8 2.2005
R349 drain_right.n9 drain_right.t7 2.2005
R350 drain_right.n11 drain_right.t12 2.2005
R351 drain_right.n11 drain_right.t14 2.2005
R352 drain_right.n13 drain_right.t16 2.2005
R353 drain_right.n13 drain_right.t13 2.2005
R354 drain_right.n15 drain_right.t19 2.2005
R355 drain_right.n15 drain_right.t18 2.2005
R356 drain_right.n16 drain_right.n14 0.802224
R357 drain_right.n14 drain_right.n12 0.802224
R358 drain_right.n12 drain_right.n10 0.802224
R359 drain_right.n7 drain_right.n6 0.746878
R360 drain_right.n7 drain_right.n2 0.746878
C0 drain_right plus 0.431663f
C1 drain_right drain_left 1.48676f
C2 drain_right source 20.5405f
C3 plus minus 6.0372f
C4 minus drain_left 0.173552f
C5 minus source 8.968571f
C6 plus drain_left 9.05917f
C7 plus source 8.982611f
C8 source drain_left 20.538599f
C9 drain_right minus 8.784531f
C10 drain_right a_n2762_n2688# 6.58157f
C11 drain_left a_n2762_n2688# 6.9782f
C12 source a_n2762_n2688# 7.638422f
C13 minus a_n2762_n2688# 10.853968f
C14 plus a_n2762_n2688# 12.56604f
C15 drain_right.t9 a_n2762_n2688# 0.198859f
C16 drain_right.t0 a_n2762_n2688# 0.198859f
C17 drain_right.n0 a_n2762_n2688# 1.74394f
C18 drain_right.t15 a_n2762_n2688# 0.198859f
C19 drain_right.t3 a_n2762_n2688# 0.198859f
C20 drain_right.n1 a_n2762_n2688# 1.73935f
C21 drain_right.n2 a_n2762_n2688# 0.739421f
C22 drain_right.t1 a_n2762_n2688# 0.198859f
C23 drain_right.t2 a_n2762_n2688# 0.198859f
C24 drain_right.n3 a_n2762_n2688# 1.73935f
C25 drain_right.t17 a_n2762_n2688# 0.198859f
C26 drain_right.t10 a_n2762_n2688# 0.198859f
C27 drain_right.n4 a_n2762_n2688# 1.74394f
C28 drain_right.t11 a_n2762_n2688# 0.198859f
C29 drain_right.t4 a_n2762_n2688# 0.198859f
C30 drain_right.n5 a_n2762_n2688# 1.73935f
C31 drain_right.n6 a_n2762_n2688# 0.739421f
C32 drain_right.n7 a_n2762_n2688# 1.70641f
C33 drain_right.t6 a_n2762_n2688# 0.198859f
C34 drain_right.t5 a_n2762_n2688# 0.198859f
C35 drain_right.n8 a_n2762_n2688# 1.74394f
C36 drain_right.t8 a_n2762_n2688# 0.198859f
C37 drain_right.t7 a_n2762_n2688# 0.198859f
C38 drain_right.n9 a_n2762_n2688# 1.73936f
C39 drain_right.n10 a_n2762_n2688# 0.743539f
C40 drain_right.t12 a_n2762_n2688# 0.198859f
C41 drain_right.t14 a_n2762_n2688# 0.198859f
C42 drain_right.n11 a_n2762_n2688# 1.73936f
C43 drain_right.n12 a_n2762_n2688# 0.368429f
C44 drain_right.t16 a_n2762_n2688# 0.198859f
C45 drain_right.t13 a_n2762_n2688# 0.198859f
C46 drain_right.n13 a_n2762_n2688# 1.73936f
C47 drain_right.n14 a_n2762_n2688# 0.368429f
C48 drain_right.t19 a_n2762_n2688# 0.198859f
C49 drain_right.t18 a_n2762_n2688# 0.198859f
C50 drain_right.n15 a_n2762_n2688# 1.73936f
C51 drain_right.n16 a_n2762_n2688# 0.612245f
C52 minus.n0 a_n2762_n2688# 0.055886f
C53 minus.n1 a_n2762_n2688# 0.009526f
C54 minus.t3 a_n2762_n2688# 0.650126f
C55 minus.n2 a_n2762_n2688# 0.04198f
C56 minus.n3 a_n2762_n2688# 0.009526f
C57 minus.t7 a_n2762_n2688# 0.650126f
C58 minus.n4 a_n2762_n2688# 0.04198f
C59 minus.n5 a_n2762_n2688# 0.009526f
C60 minus.t11 a_n2762_n2688# 0.650126f
C61 minus.t14 a_n2762_n2688# 0.666397f
C62 minus.n6 a_n2762_n2688# 0.259807f
C63 minus.t13 a_n2762_n2688# 0.650126f
C64 minus.n7 a_n2762_n2688# 0.284703f
C65 minus.t12 a_n2762_n2688# 0.650126f
C66 minus.n8 a_n2762_n2688# 0.275824f
C67 minus.n9 a_n2762_n2688# 0.179185f
C68 minus.n10 a_n2762_n2688# 0.04198f
C69 minus.n11 a_n2762_n2688# 0.04198f
C70 minus.n12 a_n2762_n2688# 0.276988f
C71 minus.n13 a_n2762_n2688# 0.009526f
C72 minus.t5 a_n2762_n2688# 0.650126f
C73 minus.n14 a_n2762_n2688# 0.276988f
C74 minus.n15 a_n2762_n2688# 0.04198f
C75 minus.n16 a_n2762_n2688# 0.04198f
C76 minus.n17 a_n2762_n2688# 0.04198f
C77 minus.n18 a_n2762_n2688# 0.276988f
C78 minus.n19 a_n2762_n2688# 0.009526f
C79 minus.t6 a_n2762_n2688# 0.650126f
C80 minus.n20 a_n2762_n2688# 0.276988f
C81 minus.n21 a_n2762_n2688# 0.04198f
C82 minus.n22 a_n2762_n2688# 0.04198f
C83 minus.n23 a_n2762_n2688# 0.056018f
C84 minus.n24 a_n2762_n2688# 0.275824f
C85 minus.t1 a_n2762_n2688# 0.650126f
C86 minus.n25 a_n2762_n2688# 0.284703f
C87 minus.t0 a_n2762_n2688# 0.650126f
C88 minus.n26 a_n2762_n2688# 0.275177f
C89 minus.n27 a_n2762_n2688# 1.58175f
C90 minus.n28 a_n2762_n2688# 0.055886f
C91 minus.n29 a_n2762_n2688# 0.009526f
C92 minus.n30 a_n2762_n2688# 0.04198f
C93 minus.n31 a_n2762_n2688# 0.009526f
C94 minus.n32 a_n2762_n2688# 0.04198f
C95 minus.n33 a_n2762_n2688# 0.009526f
C96 minus.t10 a_n2762_n2688# 0.666397f
C97 minus.n34 a_n2762_n2688# 0.259807f
C98 minus.t19 a_n2762_n2688# 0.650126f
C99 minus.n35 a_n2762_n2688# 0.284703f
C100 minus.t4 a_n2762_n2688# 0.650126f
C101 minus.n36 a_n2762_n2688# 0.275824f
C102 minus.n37 a_n2762_n2688# 0.179185f
C103 minus.n38 a_n2762_n2688# 0.04198f
C104 minus.n39 a_n2762_n2688# 0.04198f
C105 minus.t16 a_n2762_n2688# 0.650126f
C106 minus.n40 a_n2762_n2688# 0.276988f
C107 minus.n41 a_n2762_n2688# 0.009526f
C108 minus.t18 a_n2762_n2688# 0.650126f
C109 minus.n42 a_n2762_n2688# 0.276988f
C110 minus.n43 a_n2762_n2688# 0.04198f
C111 minus.n44 a_n2762_n2688# 0.04198f
C112 minus.n45 a_n2762_n2688# 0.04198f
C113 minus.t17 a_n2762_n2688# 0.650126f
C114 minus.n46 a_n2762_n2688# 0.276988f
C115 minus.n47 a_n2762_n2688# 0.009526f
C116 minus.t8 a_n2762_n2688# 0.650126f
C117 minus.n48 a_n2762_n2688# 0.276988f
C118 minus.n49 a_n2762_n2688# 0.04198f
C119 minus.n50 a_n2762_n2688# 0.04198f
C120 minus.n51 a_n2762_n2688# 0.056018f
C121 minus.t15 a_n2762_n2688# 0.650126f
C122 minus.n52 a_n2762_n2688# 0.275824f
C123 minus.t2 a_n2762_n2688# 0.650126f
C124 minus.n53 a_n2762_n2688# 0.284703f
C125 minus.t9 a_n2762_n2688# 0.650126f
C126 minus.n54 a_n2762_n2688# 0.275177f
C127 minus.n55 a_n2762_n2688# 0.301203f
C128 minus.n56 a_n2762_n2688# 1.89335f
C129 drain_left.t9 a_n2762_n2688# 0.200148f
C130 drain_left.t18 a_n2762_n2688# 0.200148f
C131 drain_left.n0 a_n2762_n2688# 1.75524f
C132 drain_left.t2 a_n2762_n2688# 0.200148f
C133 drain_left.t10 a_n2762_n2688# 0.200148f
C134 drain_left.n1 a_n2762_n2688# 1.75063f
C135 drain_left.n2 a_n2762_n2688# 0.744214f
C136 drain_left.t0 a_n2762_n2688# 0.200148f
C137 drain_left.t1 a_n2762_n2688# 0.200148f
C138 drain_left.n3 a_n2762_n2688# 1.75063f
C139 drain_left.t13 a_n2762_n2688# 0.200148f
C140 drain_left.t4 a_n2762_n2688# 0.200148f
C141 drain_left.n4 a_n2762_n2688# 1.75524f
C142 drain_left.t3 a_n2762_n2688# 0.200148f
C143 drain_left.t11 a_n2762_n2688# 0.200148f
C144 drain_left.n5 a_n2762_n2688# 1.75063f
C145 drain_left.n6 a_n2762_n2688# 0.744214f
C146 drain_left.n7 a_n2762_n2688# 1.77454f
C147 drain_left.t5 a_n2762_n2688# 0.200148f
C148 drain_left.t6 a_n2762_n2688# 0.200148f
C149 drain_left.n8 a_n2762_n2688# 1.75525f
C150 drain_left.t7 a_n2762_n2688# 0.200148f
C151 drain_left.t8 a_n2762_n2688# 0.200148f
C152 drain_left.n9 a_n2762_n2688# 1.75063f
C153 drain_left.n10 a_n2762_n2688# 0.748351f
C154 drain_left.t12 a_n2762_n2688# 0.200148f
C155 drain_left.t14 a_n2762_n2688# 0.200148f
C156 drain_left.n11 a_n2762_n2688# 1.75063f
C157 drain_left.n12 a_n2762_n2688# 0.370817f
C158 drain_left.t15 a_n2762_n2688# 0.200148f
C159 drain_left.t16 a_n2762_n2688# 0.200148f
C160 drain_left.n13 a_n2762_n2688# 1.75063f
C161 drain_left.n14 a_n2762_n2688# 0.370817f
C162 drain_left.t17 a_n2762_n2688# 0.200148f
C163 drain_left.t19 a_n2762_n2688# 0.200148f
C164 drain_left.n15 a_n2762_n2688# 1.75062f
C165 drain_left.n16 a_n2762_n2688# 0.616221f
C166 source.t25 a_n2762_n2688# 1.9234f
C167 source.n0 a_n2762_n2688# 1.14136f
C168 source.t31 a_n2762_n2688# 0.180373f
C169 source.t29 a_n2762_n2688# 0.180373f
C170 source.n1 a_n2762_n2688# 1.50996f
C171 source.n2 a_n2762_n2688# 0.367408f
C172 source.t35 a_n2762_n2688# 0.180373f
C173 source.t21 a_n2762_n2688# 0.180373f
C174 source.n3 a_n2762_n2688# 1.50996f
C175 source.n4 a_n2762_n2688# 0.367408f
C176 source.t27 a_n2762_n2688# 0.180373f
C177 source.t37 a_n2762_n2688# 0.180373f
C178 source.n5 a_n2762_n2688# 1.50996f
C179 source.n6 a_n2762_n2688# 0.367408f
C180 source.t36 a_n2762_n2688# 0.180373f
C181 source.t39 a_n2762_n2688# 0.180373f
C182 source.n7 a_n2762_n2688# 1.50996f
C183 source.n8 a_n2762_n2688# 0.367408f
C184 source.t30 a_n2762_n2688# 1.9234f
C185 source.n9 a_n2762_n2688# 0.418771f
C186 source.t11 a_n2762_n2688# 1.9234f
C187 source.n10 a_n2762_n2688# 0.418771f
C188 source.t1 a_n2762_n2688# 0.180373f
C189 source.t17 a_n2762_n2688# 0.180373f
C190 source.n11 a_n2762_n2688# 1.50996f
C191 source.n12 a_n2762_n2688# 0.367408f
C192 source.t3 a_n2762_n2688# 0.180373f
C193 source.t4 a_n2762_n2688# 0.180373f
C194 source.n13 a_n2762_n2688# 1.50996f
C195 source.n14 a_n2762_n2688# 0.367408f
C196 source.t5 a_n2762_n2688# 0.180373f
C197 source.t16 a_n2762_n2688# 0.180373f
C198 source.n15 a_n2762_n2688# 1.50996f
C199 source.n16 a_n2762_n2688# 0.367408f
C200 source.t0 a_n2762_n2688# 0.180373f
C201 source.t2 a_n2762_n2688# 0.180373f
C202 source.n17 a_n2762_n2688# 1.50996f
C203 source.n18 a_n2762_n2688# 0.367408f
C204 source.t12 a_n2762_n2688# 1.9234f
C205 source.n19 a_n2762_n2688# 1.51677f
C206 source.t20 a_n2762_n2688# 1.9234f
C207 source.n20 a_n2762_n2688# 1.51678f
C208 source.t38 a_n2762_n2688# 0.180373f
C209 source.t32 a_n2762_n2688# 0.180373f
C210 source.n21 a_n2762_n2688# 1.50996f
C211 source.n22 a_n2762_n2688# 0.367412f
C212 source.t23 a_n2762_n2688# 0.180373f
C213 source.t34 a_n2762_n2688# 0.180373f
C214 source.n23 a_n2762_n2688# 1.50996f
C215 source.n24 a_n2762_n2688# 0.367412f
C216 source.t33 a_n2762_n2688# 0.180373f
C217 source.t28 a_n2762_n2688# 0.180373f
C218 source.n25 a_n2762_n2688# 1.50996f
C219 source.n26 a_n2762_n2688# 0.367412f
C220 source.t26 a_n2762_n2688# 0.180373f
C221 source.t24 a_n2762_n2688# 0.180373f
C222 source.n27 a_n2762_n2688# 1.50996f
C223 source.n28 a_n2762_n2688# 0.367412f
C224 source.t22 a_n2762_n2688# 1.9234f
C225 source.n29 a_n2762_n2688# 0.418775f
C226 source.t13 a_n2762_n2688# 1.9234f
C227 source.n30 a_n2762_n2688# 0.418775f
C228 source.t14 a_n2762_n2688# 0.180373f
C229 source.t9 a_n2762_n2688# 0.180373f
C230 source.n31 a_n2762_n2688# 1.50996f
C231 source.n32 a_n2762_n2688# 0.367412f
C232 source.t18 a_n2762_n2688# 0.180373f
C233 source.t7 a_n2762_n2688# 0.180373f
C234 source.n33 a_n2762_n2688# 1.50996f
C235 source.n34 a_n2762_n2688# 0.367412f
C236 source.t19 a_n2762_n2688# 0.180373f
C237 source.t6 a_n2762_n2688# 0.180373f
C238 source.n35 a_n2762_n2688# 1.50996f
C239 source.n36 a_n2762_n2688# 0.367412f
C240 source.t8 a_n2762_n2688# 0.180373f
C241 source.t15 a_n2762_n2688# 0.180373f
C242 source.n37 a_n2762_n2688# 1.50996f
C243 source.n38 a_n2762_n2688# 0.367412f
C244 source.t10 a_n2762_n2688# 1.9234f
C245 source.n39 a_n2762_n2688# 0.578689f
C246 source.n40 a_n2762_n2688# 1.33155f
C247 plus.n0 a_n2762_n2688# 0.056793f
C248 plus.t0 a_n2762_n2688# 0.660677f
C249 plus.t2 a_n2762_n2688# 0.660677f
C250 plus.t3 a_n2762_n2688# 0.660677f
C251 plus.n1 a_n2762_n2688# 0.056927f
C252 plus.t4 a_n2762_n2688# 0.660677f
C253 plus.n2 a_n2762_n2688# 0.281484f
C254 plus.n3 a_n2762_n2688# 0.042662f
C255 plus.t5 a_n2762_n2688# 0.660677f
C256 plus.t7 a_n2762_n2688# 0.660677f
C257 plus.n4 a_n2762_n2688# 0.281484f
C258 plus.n5 a_n2762_n2688# 0.042662f
C259 plus.t11 a_n2762_n2688# 0.660677f
C260 plus.t12 a_n2762_n2688# 0.660677f
C261 plus.n6 a_n2762_n2688# 0.2803f
C262 plus.t13 a_n2762_n2688# 0.660677f
C263 plus.n7 a_n2762_n2688# 0.289324f
C264 plus.t14 a_n2762_n2688# 0.677213f
C265 plus.n8 a_n2762_n2688# 0.264023f
C266 plus.n9 a_n2762_n2688# 0.182093f
C267 plus.n10 a_n2762_n2688# 0.042662f
C268 plus.n11 a_n2762_n2688# 0.009681f
C269 plus.n12 a_n2762_n2688# 0.281484f
C270 plus.n13 a_n2762_n2688# 0.009681f
C271 plus.n14 a_n2762_n2688# 0.042662f
C272 plus.n15 a_n2762_n2688# 0.042662f
C273 plus.n16 a_n2762_n2688# 0.042662f
C274 plus.n17 a_n2762_n2688# 0.009681f
C275 plus.n18 a_n2762_n2688# 0.281484f
C276 plus.n19 a_n2762_n2688# 0.009681f
C277 plus.n20 a_n2762_n2688# 0.042662f
C278 plus.n21 a_n2762_n2688# 0.042662f
C279 plus.n22 a_n2762_n2688# 0.042662f
C280 plus.n23 a_n2762_n2688# 0.009681f
C281 plus.n24 a_n2762_n2688# 0.2803f
C282 plus.n25 a_n2762_n2688# 0.289324f
C283 plus.n26 a_n2762_n2688# 0.279643f
C284 plus.n27 a_n2762_n2688# 0.446658f
C285 plus.n28 a_n2762_n2688# 0.056793f
C286 plus.t10 a_n2762_n2688# 0.660677f
C287 plus.t1 a_n2762_n2688# 0.660677f
C288 plus.n29 a_n2762_n2688# 0.056927f
C289 plus.t17 a_n2762_n2688# 0.660677f
C290 plus.t9 a_n2762_n2688# 0.660677f
C291 plus.n30 a_n2762_n2688# 0.281484f
C292 plus.n31 a_n2762_n2688# 0.042662f
C293 plus.t19 a_n2762_n2688# 0.660677f
C294 plus.t18 a_n2762_n2688# 0.660677f
C295 plus.n32 a_n2762_n2688# 0.281484f
C296 plus.n33 a_n2762_n2688# 0.042662f
C297 plus.t16 a_n2762_n2688# 0.660677f
C298 plus.t8 a_n2762_n2688# 0.660677f
C299 plus.n34 a_n2762_n2688# 0.2803f
C300 plus.t6 a_n2762_n2688# 0.660677f
C301 plus.n35 a_n2762_n2688# 0.289324f
C302 plus.t15 a_n2762_n2688# 0.677213f
C303 plus.n36 a_n2762_n2688# 0.264023f
C304 plus.n37 a_n2762_n2688# 0.182093f
C305 plus.n38 a_n2762_n2688# 0.042662f
C306 plus.n39 a_n2762_n2688# 0.009681f
C307 plus.n40 a_n2762_n2688# 0.281484f
C308 plus.n41 a_n2762_n2688# 0.009681f
C309 plus.n42 a_n2762_n2688# 0.042662f
C310 plus.n43 a_n2762_n2688# 0.042662f
C311 plus.n44 a_n2762_n2688# 0.042662f
C312 plus.n45 a_n2762_n2688# 0.009681f
C313 plus.n46 a_n2762_n2688# 0.281484f
C314 plus.n47 a_n2762_n2688# 0.009681f
C315 plus.n48 a_n2762_n2688# 0.042662f
C316 plus.n49 a_n2762_n2688# 0.042662f
C317 plus.n50 a_n2762_n2688# 0.042662f
C318 plus.n51 a_n2762_n2688# 0.009681f
C319 plus.n52 a_n2762_n2688# 0.2803f
C320 plus.n53 a_n2762_n2688# 0.289324f
C321 plus.n54 a_n2762_n2688# 0.279643f
C322 plus.n55 a_n2762_n2688# 1.41314f
.ends

