* NGSPICE file created from diffpair561.ext - technology: sky130A

.subckt diffpair561 minus drain_right drain_left source plus
X0 drain_right minus source a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X1 drain_left plus source a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X2 source plus drain_left a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X3 drain_right minus source a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X4 a_n1106_n4892# a_n1106_n4892# a_n1106_n4892# a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=76 ps=327.6 w=20 l=0.15
X5 source plus drain_left a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X6 drain_left plus source a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X7 source minus drain_right a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X8 a_n1106_n4892# a_n1106_n4892# a_n1106_n4892# a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X9 a_n1106_n4892# a_n1106_n4892# a_n1106_n4892# a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X10 a_n1106_n4892# a_n1106_n4892# a_n1106_n4892# a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X11 source minus drain_right a_n1106_n4892# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
.ends

