* NGSPICE file created from diffpair489.ext - technology: sky130A

.subckt diffpair489 minus drain_right drain_left source plus
X0 source.t47 minus.t0 drain_right.t13 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X1 source.t46 minus.t1 drain_right.t12 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X2 drain_right.t17 minus.t2 source.t45 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X3 source.t0 plus.t0 drain_left.t23 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X4 drain_right.t16 minus.t3 source.t44 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X5 source.t43 minus.t4 drain_right.t23 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X6 source.t15 plus.t1 drain_left.t22 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X7 drain_left.t21 plus.t2 source.t19 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X8 drain_left.t20 plus.t3 source.t23 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X9 a_n2406_n3888# a_n2406_n3888# a_n2406_n3888# a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=57 ps=247.6 w=15 l=0.15
X10 a_n2406_n3888# a_n2406_n3888# a_n2406_n3888# a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X11 drain_left.t19 plus.t4 source.t16 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X12 source.t1 plus.t5 drain_left.t18 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X13 source.t42 minus.t5 drain_right.t22 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X14 source.t5 plus.t6 drain_left.t17 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X15 drain_right.t19 minus.t6 source.t41 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X16 drain_right.t18 minus.t7 source.t40 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X17 drain_right.t1 minus.t8 source.t39 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X18 source.t6 plus.t7 drain_left.t16 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X19 source.t38 minus.t9 drain_right.t0 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X20 source.t37 minus.t10 drain_right.t15 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X21 drain_left.t15 plus.t8 source.t11 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X22 drain_right.t14 minus.t11 source.t36 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X23 a_n2406_n3888# a_n2406_n3888# a_n2406_n3888# a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X24 drain_left.t14 plus.t9 source.t8 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X25 source.t2 plus.t10 drain_left.t13 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X26 drain_right.t5 minus.t12 source.t35 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X27 drain_right.t4 minus.t13 source.t34 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X28 source.t33 minus.t14 drain_right.t7 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X29 drain_left.t12 plus.t11 source.t10 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X30 source.t13 plus.t12 drain_left.t11 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X31 source.t32 minus.t15 drain_right.t6 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X32 source.t31 minus.t16 drain_right.t9 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X33 drain_left.t10 plus.t13 source.t18 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X34 source.t30 minus.t17 drain_right.t8 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X35 drain_right.t3 minus.t18 source.t29 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X36 drain_left.t9 plus.t14 source.t20 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X37 drain_right.t2 minus.t19 source.t28 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X38 drain_left.t8 plus.t15 source.t12 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X39 source.t17 plus.t16 drain_left.t7 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X40 source.t21 plus.t17 drain_left.t6 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X41 drain_right.t11 minus.t20 source.t27 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X42 source.t26 minus.t21 drain_right.t10 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X43 drain_right.t21 minus.t22 source.t25 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X44 source.t22 plus.t18 drain_left.t5 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X45 drain_left.t4 plus.t19 source.t4 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X46 drain_left.t3 plus.t20 source.t9 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X47 source.t3 plus.t21 drain_left.t2 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X48 drain_left.t1 plus.t22 source.t7 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X49 source.t14 plus.t23 drain_left.t0 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X50 source.t24 minus.t23 drain_right.t20 a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X51 a_n2406_n3888# a_n2406_n3888# a_n2406_n3888# a_n2406_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
R0 minus.n35 minus.t16 2666.34
R1 minus.n8 minus.t6 2666.34
R2 minus.n72 minus.t8 2666.34
R3 minus.n43 minus.t4 2666.34
R4 minus.n34 minus.t19 2618.87
R5 minus.n32 minus.t21 2618.87
R6 minus.n3 minus.t11 2618.87
R7 minus.n26 minus.t15 2618.87
R8 minus.n24 minus.t13 2618.87
R9 minus.n6 minus.t17 2618.87
R10 minus.n18 minus.t7 2618.87
R11 minus.n16 minus.t9 2618.87
R12 minus.n9 minus.t12 2618.87
R13 minus.n10 minus.t5 2618.87
R14 minus.n71 minus.t1 2618.87
R15 minus.n69 minus.t22 2618.87
R16 minus.n63 minus.t14 2618.87
R17 minus.n62 minus.t3 2618.87
R18 minus.n60 minus.t0 2618.87
R19 minus.n54 minus.t20 2618.87
R20 minus.n53 minus.t10 2618.87
R21 minus.n51 minus.t2 2618.87
R22 minus.n45 minus.t23 2618.87
R23 minus.n44 minus.t18 2618.87
R24 minus.n12 minus.n8 161.489
R25 minus.n47 minus.n43 161.489
R26 minus.n36 minus.n35 161.3
R27 minus.n33 minus.n0 161.3
R28 minus.n31 minus.n30 161.3
R29 minus.n29 minus.n1 161.3
R30 minus.n28 minus.n27 161.3
R31 minus.n25 minus.n2 161.3
R32 minus.n23 minus.n22 161.3
R33 minus.n21 minus.n4 161.3
R34 minus.n20 minus.n19 161.3
R35 minus.n17 minus.n5 161.3
R36 minus.n15 minus.n14 161.3
R37 minus.n13 minus.n7 161.3
R38 minus.n12 minus.n11 161.3
R39 minus.n73 minus.n72 161.3
R40 minus.n70 minus.n37 161.3
R41 minus.n68 minus.n67 161.3
R42 minus.n66 minus.n38 161.3
R43 minus.n65 minus.n64 161.3
R44 minus.n61 minus.n39 161.3
R45 minus.n59 minus.n58 161.3
R46 minus.n57 minus.n40 161.3
R47 minus.n56 minus.n55 161.3
R48 minus.n52 minus.n41 161.3
R49 minus.n50 minus.n49 161.3
R50 minus.n48 minus.n42 161.3
R51 minus.n47 minus.n46 161.3
R52 minus.n31 minus.n1 73.0308
R53 minus.n23 minus.n4 73.0308
R54 minus.n15 minus.n7 73.0308
R55 minus.n50 minus.n42 73.0308
R56 minus.n59 minus.n40 73.0308
R57 minus.n68 minus.n38 73.0308
R58 minus.n33 minus.n32 69.3793
R59 minus.n11 minus.n9 69.3793
R60 minus.n46 minus.n45 69.3793
R61 minus.n70 minus.n69 69.3793
R62 minus.n25 minus.n24 62.0763
R63 minus.n19 minus.n6 62.0763
R64 minus.n55 minus.n54 62.0763
R65 minus.n61 minus.n60 62.0763
R66 minus.n27 minus.n3 54.7732
R67 minus.n17 minus.n16 54.7732
R68 minus.n52 minus.n51 54.7732
R69 minus.n64 minus.n63 54.7732
R70 minus.n35 minus.n34 47.4702
R71 minus.n10 minus.n8 47.4702
R72 minus.n44 minus.n43 47.4702
R73 minus.n72 minus.n71 47.4702
R74 minus.n74 minus.n36 40.5308
R75 minus.n27 minus.n26 40.1672
R76 minus.n18 minus.n17 40.1672
R77 minus.n53 minus.n52 40.1672
R78 minus.n64 minus.n62 40.1672
R79 minus.n26 minus.n25 32.8641
R80 minus.n19 minus.n18 32.8641
R81 minus.n55 minus.n53 32.8641
R82 minus.n62 minus.n61 32.8641
R83 minus.n34 minus.n33 25.5611
R84 minus.n11 minus.n10 25.5611
R85 minus.n46 minus.n44 25.5611
R86 minus.n71 minus.n70 25.5611
R87 minus.n3 minus.n1 18.2581
R88 minus.n16 minus.n15 18.2581
R89 minus.n51 minus.n50 18.2581
R90 minus.n63 minus.n38 18.2581
R91 minus.n24 minus.n23 10.955
R92 minus.n6 minus.n4 10.955
R93 minus.n54 minus.n40 10.955
R94 minus.n60 minus.n59 10.955
R95 minus.n74 minus.n73 6.52323
R96 minus.n32 minus.n31 3.65202
R97 minus.n9 minus.n7 3.65202
R98 minus.n45 minus.n42 3.65202
R99 minus.n69 minus.n68 3.65202
R100 minus.n36 minus.n0 0.189894
R101 minus.n30 minus.n0 0.189894
R102 minus.n30 minus.n29 0.189894
R103 minus.n29 minus.n28 0.189894
R104 minus.n28 minus.n2 0.189894
R105 minus.n22 minus.n2 0.189894
R106 minus.n22 minus.n21 0.189894
R107 minus.n21 minus.n20 0.189894
R108 minus.n20 minus.n5 0.189894
R109 minus.n14 minus.n5 0.189894
R110 minus.n14 minus.n13 0.189894
R111 minus.n13 minus.n12 0.189894
R112 minus.n48 minus.n47 0.189894
R113 minus.n49 minus.n48 0.189894
R114 minus.n49 minus.n41 0.189894
R115 minus.n56 minus.n41 0.189894
R116 minus.n57 minus.n56 0.189894
R117 minus.n58 minus.n57 0.189894
R118 minus.n58 minus.n39 0.189894
R119 minus.n65 minus.n39 0.189894
R120 minus.n66 minus.n65 0.189894
R121 minus.n67 minus.n66 0.189894
R122 minus.n67 minus.n37 0.189894
R123 minus.n73 minus.n37 0.189894
R124 minus minus.n74 0.188
R125 drain_right.n13 drain_right.n11 61.44
R126 drain_right.n7 drain_right.n5 61.4399
R127 drain_right.n2 drain_right.n0 61.4399
R128 drain_right.n13 drain_right.n12 60.8798
R129 drain_right.n15 drain_right.n14 60.8798
R130 drain_right.n17 drain_right.n16 60.8798
R131 drain_right.n19 drain_right.n18 60.8798
R132 drain_right.n21 drain_right.n20 60.8798
R133 drain_right.n7 drain_right.n6 60.8796
R134 drain_right.n9 drain_right.n8 60.8796
R135 drain_right.n4 drain_right.n3 60.8796
R136 drain_right.n2 drain_right.n1 60.8796
R137 drain_right drain_right.n10 34.4098
R138 drain_right drain_right.n21 6.21356
R139 drain_right.n5 drain_right.t12 2.0005
R140 drain_right.n5 drain_right.t1 2.0005
R141 drain_right.n6 drain_right.t7 2.0005
R142 drain_right.n6 drain_right.t21 2.0005
R143 drain_right.n8 drain_right.t13 2.0005
R144 drain_right.n8 drain_right.t16 2.0005
R145 drain_right.n3 drain_right.t15 2.0005
R146 drain_right.n3 drain_right.t11 2.0005
R147 drain_right.n1 drain_right.t20 2.0005
R148 drain_right.n1 drain_right.t17 2.0005
R149 drain_right.n0 drain_right.t23 2.0005
R150 drain_right.n0 drain_right.t3 2.0005
R151 drain_right.n11 drain_right.t22 2.0005
R152 drain_right.n11 drain_right.t19 2.0005
R153 drain_right.n12 drain_right.t0 2.0005
R154 drain_right.n12 drain_right.t5 2.0005
R155 drain_right.n14 drain_right.t8 2.0005
R156 drain_right.n14 drain_right.t18 2.0005
R157 drain_right.n16 drain_right.t6 2.0005
R158 drain_right.n16 drain_right.t4 2.0005
R159 drain_right.n18 drain_right.t10 2.0005
R160 drain_right.n18 drain_right.t14 2.0005
R161 drain_right.n20 drain_right.t9 2.0005
R162 drain_right.n20 drain_right.t2 2.0005
R163 drain_right.n9 drain_right.n7 0.560845
R164 drain_right.n4 drain_right.n2 0.560845
R165 drain_right.n21 drain_right.n19 0.560845
R166 drain_right.n19 drain_right.n17 0.560845
R167 drain_right.n17 drain_right.n15 0.560845
R168 drain_right.n15 drain_right.n13 0.560845
R169 drain_right.n10 drain_right.n9 0.225326
R170 drain_right.n10 drain_right.n4 0.225326
R171 source.n11 source.t2 46.201
R172 source.n12 source.t41 46.201
R173 source.n23 source.t31 46.201
R174 source.n47 source.t39 46.2008
R175 source.n36 source.t43 46.2008
R176 source.n35 source.t10 46.2008
R177 source.n24 source.t5 46.2008
R178 source.n0 source.t7 46.2008
R179 source.n2 source.n1 44.201
R180 source.n4 source.n3 44.201
R181 source.n6 source.n5 44.201
R182 source.n8 source.n7 44.201
R183 source.n10 source.n9 44.201
R184 source.n14 source.n13 44.201
R185 source.n16 source.n15 44.201
R186 source.n18 source.n17 44.201
R187 source.n20 source.n19 44.201
R188 source.n22 source.n21 44.201
R189 source.n46 source.n45 44.2008
R190 source.n44 source.n43 44.2008
R191 source.n42 source.n41 44.2008
R192 source.n40 source.n39 44.2008
R193 source.n38 source.n37 44.2008
R194 source.n34 source.n33 44.2008
R195 source.n32 source.n31 44.2008
R196 source.n30 source.n29 44.2008
R197 source.n28 source.n27 44.2008
R198 source.n26 source.n25 44.2008
R199 source.n24 source.n23 24.1208
R200 source.n48 source.n0 18.5777
R201 source.n48 source.n47 5.5436
R202 source.n45 source.t25 2.0005
R203 source.n45 source.t46 2.0005
R204 source.n43 source.t44 2.0005
R205 source.n43 source.t33 2.0005
R206 source.n41 source.t27 2.0005
R207 source.n41 source.t47 2.0005
R208 source.n39 source.t45 2.0005
R209 source.n39 source.t37 2.0005
R210 source.n37 source.t29 2.0005
R211 source.n37 source.t24 2.0005
R212 source.n33 source.t23 2.0005
R213 source.n33 source.t3 2.0005
R214 source.n31 source.t20 2.0005
R215 source.n31 source.t6 2.0005
R216 source.n29 source.t16 2.0005
R217 source.n29 source.t15 2.0005
R218 source.n27 source.t11 2.0005
R219 source.n27 source.t1 2.0005
R220 source.n25 source.t19 2.0005
R221 source.n25 source.t0 2.0005
R222 source.n1 source.t12 2.0005
R223 source.n1 source.t13 2.0005
R224 source.n3 source.t8 2.0005
R225 source.n3 source.t22 2.0005
R226 source.n5 source.t4 2.0005
R227 source.n5 source.t17 2.0005
R228 source.n7 source.t18 2.0005
R229 source.n7 source.t14 2.0005
R230 source.n9 source.t9 2.0005
R231 source.n9 source.t21 2.0005
R232 source.n13 source.t35 2.0005
R233 source.n13 source.t42 2.0005
R234 source.n15 source.t40 2.0005
R235 source.n15 source.t38 2.0005
R236 source.n17 source.t34 2.0005
R237 source.n17 source.t30 2.0005
R238 source.n19 source.t36 2.0005
R239 source.n19 source.t32 2.0005
R240 source.n21 source.t28 2.0005
R241 source.n21 source.t26 2.0005
R242 source.n23 source.n22 0.560845
R243 source.n22 source.n20 0.560845
R244 source.n20 source.n18 0.560845
R245 source.n18 source.n16 0.560845
R246 source.n16 source.n14 0.560845
R247 source.n14 source.n12 0.560845
R248 source.n11 source.n10 0.560845
R249 source.n10 source.n8 0.560845
R250 source.n8 source.n6 0.560845
R251 source.n6 source.n4 0.560845
R252 source.n4 source.n2 0.560845
R253 source.n2 source.n0 0.560845
R254 source.n26 source.n24 0.560845
R255 source.n28 source.n26 0.560845
R256 source.n30 source.n28 0.560845
R257 source.n32 source.n30 0.560845
R258 source.n34 source.n32 0.560845
R259 source.n35 source.n34 0.560845
R260 source.n38 source.n36 0.560845
R261 source.n40 source.n38 0.560845
R262 source.n42 source.n40 0.560845
R263 source.n44 source.n42 0.560845
R264 source.n46 source.n44 0.560845
R265 source.n47 source.n46 0.560845
R266 source.n12 source.n11 0.470328
R267 source.n36 source.n35 0.470328
R268 source source.n48 0.188
R269 plus.n6 plus.t10 2666.34
R270 plus.n35 plus.t22 2666.34
R271 plus.n45 plus.t11 2666.34
R272 plus.n72 plus.t6 2666.34
R273 plus.n7 plus.t20 2618.87
R274 plus.n8 plus.t17 2618.87
R275 plus.n14 plus.t13 2618.87
R276 plus.n16 plus.t23 2618.87
R277 plus.n17 plus.t19 2618.87
R278 plus.n23 plus.t16 2618.87
R279 plus.n25 plus.t9 2618.87
R280 plus.n26 plus.t18 2618.87
R281 plus.n32 plus.t15 2618.87
R282 plus.n34 plus.t12 2618.87
R283 plus.n47 plus.t21 2618.87
R284 plus.n46 plus.t3 2618.87
R285 plus.n53 plus.t7 2618.87
R286 plus.n55 plus.t14 2618.87
R287 plus.n43 plus.t1 2618.87
R288 plus.n61 plus.t4 2618.87
R289 plus.n63 plus.t5 2618.87
R290 plus.n40 plus.t8 2618.87
R291 plus.n69 plus.t0 2618.87
R292 plus.n71 plus.t2 2618.87
R293 plus.n10 plus.n6 161.489
R294 plus.n49 plus.n45 161.489
R295 plus.n10 plus.n9 161.3
R296 plus.n11 plus.n5 161.3
R297 plus.n13 plus.n12 161.3
R298 plus.n15 plus.n4 161.3
R299 plus.n19 plus.n18 161.3
R300 plus.n20 plus.n3 161.3
R301 plus.n22 plus.n21 161.3
R302 plus.n24 plus.n2 161.3
R303 plus.n28 plus.n27 161.3
R304 plus.n29 plus.n1 161.3
R305 plus.n31 plus.n30 161.3
R306 plus.n33 plus.n0 161.3
R307 plus.n36 plus.n35 161.3
R308 plus.n49 plus.n48 161.3
R309 plus.n50 plus.n44 161.3
R310 plus.n52 plus.n51 161.3
R311 plus.n54 plus.n42 161.3
R312 plus.n57 plus.n56 161.3
R313 plus.n58 plus.n41 161.3
R314 plus.n60 plus.n59 161.3
R315 plus.n62 plus.n39 161.3
R316 plus.n65 plus.n64 161.3
R317 plus.n66 plus.n38 161.3
R318 plus.n68 plus.n67 161.3
R319 plus.n70 plus.n37 161.3
R320 plus.n73 plus.n72 161.3
R321 plus.n13 plus.n5 73.0308
R322 plus.n22 plus.n3 73.0308
R323 plus.n31 plus.n1 73.0308
R324 plus.n68 plus.n38 73.0308
R325 plus.n60 plus.n41 73.0308
R326 plus.n52 plus.n44 73.0308
R327 plus.n9 plus.n8 69.3793
R328 plus.n33 plus.n32 69.3793
R329 plus.n70 plus.n69 69.3793
R330 plus.n48 plus.n46 69.3793
R331 plus.n18 plus.n17 62.0763
R332 plus.n24 plus.n23 62.0763
R333 plus.n62 plus.n61 62.0763
R334 plus.n56 plus.n43 62.0763
R335 plus.n15 plus.n14 54.7732
R336 plus.n27 plus.n26 54.7732
R337 plus.n64 plus.n40 54.7732
R338 plus.n54 plus.n53 54.7732
R339 plus.n7 plus.n6 47.4702
R340 plus.n35 plus.n34 47.4702
R341 plus.n72 plus.n71 47.4702
R342 plus.n47 plus.n45 47.4702
R343 plus.n16 plus.n15 40.1672
R344 plus.n27 plus.n25 40.1672
R345 plus.n64 plus.n63 40.1672
R346 plus.n55 plus.n54 40.1672
R347 plus plus.n73 33.2755
R348 plus.n18 plus.n16 32.8641
R349 plus.n25 plus.n24 32.8641
R350 plus.n63 plus.n62 32.8641
R351 plus.n56 plus.n55 32.8641
R352 plus.n9 plus.n7 25.5611
R353 plus.n34 plus.n33 25.5611
R354 plus.n71 plus.n70 25.5611
R355 plus.n48 plus.n47 25.5611
R356 plus.n14 plus.n13 18.2581
R357 plus.n26 plus.n1 18.2581
R358 plus.n40 plus.n38 18.2581
R359 plus.n53 plus.n52 18.2581
R360 plus plus.n36 13.3035
R361 plus.n17 plus.n3 10.955
R362 plus.n23 plus.n22 10.955
R363 plus.n61 plus.n60 10.955
R364 plus.n43 plus.n41 10.955
R365 plus.n8 plus.n5 3.65202
R366 plus.n32 plus.n31 3.65202
R367 plus.n69 plus.n68 3.65202
R368 plus.n46 plus.n44 3.65202
R369 plus.n11 plus.n10 0.189894
R370 plus.n12 plus.n11 0.189894
R371 plus.n12 plus.n4 0.189894
R372 plus.n19 plus.n4 0.189894
R373 plus.n20 plus.n19 0.189894
R374 plus.n21 plus.n20 0.189894
R375 plus.n21 plus.n2 0.189894
R376 plus.n28 plus.n2 0.189894
R377 plus.n29 plus.n28 0.189894
R378 plus.n30 plus.n29 0.189894
R379 plus.n30 plus.n0 0.189894
R380 plus.n36 plus.n0 0.189894
R381 plus.n73 plus.n37 0.189894
R382 plus.n67 plus.n37 0.189894
R383 plus.n67 plus.n66 0.189894
R384 plus.n66 plus.n65 0.189894
R385 plus.n65 plus.n39 0.189894
R386 plus.n59 plus.n39 0.189894
R387 plus.n59 plus.n58 0.189894
R388 plus.n58 plus.n57 0.189894
R389 plus.n57 plus.n42 0.189894
R390 plus.n51 plus.n42 0.189894
R391 plus.n51 plus.n50 0.189894
R392 plus.n50 plus.n49 0.189894
R393 drain_left.n13 drain_left.n11 61.4402
R394 drain_left.n7 drain_left.n5 61.4399
R395 drain_left.n2 drain_left.n0 61.4399
R396 drain_left.n19 drain_left.n18 60.8798
R397 drain_left.n17 drain_left.n16 60.8798
R398 drain_left.n15 drain_left.n14 60.8798
R399 drain_left.n13 drain_left.n12 60.8798
R400 drain_left.n21 drain_left.n20 60.8796
R401 drain_left.n7 drain_left.n6 60.8796
R402 drain_left.n9 drain_left.n8 60.8796
R403 drain_left.n4 drain_left.n3 60.8796
R404 drain_left.n2 drain_left.n1 60.8796
R405 drain_left drain_left.n10 34.9631
R406 drain_left drain_left.n21 6.21356
R407 drain_left.n5 drain_left.t2 2.0005
R408 drain_left.n5 drain_left.t12 2.0005
R409 drain_left.n6 drain_left.t16 2.0005
R410 drain_left.n6 drain_left.t20 2.0005
R411 drain_left.n8 drain_left.t22 2.0005
R412 drain_left.n8 drain_left.t9 2.0005
R413 drain_left.n3 drain_left.t18 2.0005
R414 drain_left.n3 drain_left.t19 2.0005
R415 drain_left.n1 drain_left.t23 2.0005
R416 drain_left.n1 drain_left.t15 2.0005
R417 drain_left.n0 drain_left.t17 2.0005
R418 drain_left.n0 drain_left.t21 2.0005
R419 drain_left.n20 drain_left.t11 2.0005
R420 drain_left.n20 drain_left.t1 2.0005
R421 drain_left.n18 drain_left.t5 2.0005
R422 drain_left.n18 drain_left.t8 2.0005
R423 drain_left.n16 drain_left.t7 2.0005
R424 drain_left.n16 drain_left.t14 2.0005
R425 drain_left.n14 drain_left.t0 2.0005
R426 drain_left.n14 drain_left.t4 2.0005
R427 drain_left.n12 drain_left.t6 2.0005
R428 drain_left.n12 drain_left.t10 2.0005
R429 drain_left.n11 drain_left.t13 2.0005
R430 drain_left.n11 drain_left.t3 2.0005
R431 drain_left.n9 drain_left.n7 0.560845
R432 drain_left.n4 drain_left.n2 0.560845
R433 drain_left.n15 drain_left.n13 0.560845
R434 drain_left.n17 drain_left.n15 0.560845
R435 drain_left.n19 drain_left.n17 0.560845
R436 drain_left.n21 drain_left.n19 0.560845
R437 drain_left.n10 drain_left.n9 0.225326
R438 drain_left.n10 drain_left.n4 0.225326
C0 drain_left minus 0.171476f
C1 plus minus 6.69707f
C2 source drain_right 55.747803f
C3 drain_left drain_right 1.29455f
C4 source drain_left 55.7471f
C5 plus drain_right 0.392113f
C6 source plus 5.39649f
C7 drain_left plus 6.19527f
C8 minus drain_right 5.95749f
C9 source minus 5.38245f
C10 drain_right a_n2406_n3888# 7.39722f
C11 drain_left a_n2406_n3888# 7.74279f
C12 source a_n2406_n3888# 10.64225f
C13 minus a_n2406_n3888# 9.116482f
C14 plus a_n2406_n3888# 11.536811f
C15 drain_left.t17 a_n2406_n3888# 0.507454f
C16 drain_left.t21 a_n2406_n3888# 0.507454f
C17 drain_left.n0 a_n2406_n3888# 3.3755f
C18 drain_left.t23 a_n2406_n3888# 0.507454f
C19 drain_left.t15 a_n2406_n3888# 0.507454f
C20 drain_left.n1 a_n2406_n3888# 3.37235f
C21 drain_left.n2 a_n2406_n3888# 0.675152f
C22 drain_left.t18 a_n2406_n3888# 0.507454f
C23 drain_left.t19 a_n2406_n3888# 0.507454f
C24 drain_left.n3 a_n2406_n3888# 3.37235f
C25 drain_left.n4 a_n2406_n3888# 0.305825f
C26 drain_left.t2 a_n2406_n3888# 0.507454f
C27 drain_left.t12 a_n2406_n3888# 0.507454f
C28 drain_left.n5 a_n2406_n3888# 3.3755f
C29 drain_left.t16 a_n2406_n3888# 0.507454f
C30 drain_left.t20 a_n2406_n3888# 0.507454f
C31 drain_left.n6 a_n2406_n3888# 3.37235f
C32 drain_left.n7 a_n2406_n3888# 0.675152f
C33 drain_left.t22 a_n2406_n3888# 0.507454f
C34 drain_left.t9 a_n2406_n3888# 0.507454f
C35 drain_left.n8 a_n2406_n3888# 3.37235f
C36 drain_left.n9 a_n2406_n3888# 0.305825f
C37 drain_left.n10 a_n2406_n3888# 1.7513f
C38 drain_left.t13 a_n2406_n3888# 0.507454f
C39 drain_left.t3 a_n2406_n3888# 0.507454f
C40 drain_left.n11 a_n2406_n3888# 3.3755f
C41 drain_left.t6 a_n2406_n3888# 0.507454f
C42 drain_left.t10 a_n2406_n3888# 0.507454f
C43 drain_left.n12 a_n2406_n3888# 3.37235f
C44 drain_left.n13 a_n2406_n3888# 0.675147f
C45 drain_left.t0 a_n2406_n3888# 0.507454f
C46 drain_left.t4 a_n2406_n3888# 0.507454f
C47 drain_left.n14 a_n2406_n3888# 3.37235f
C48 drain_left.n15 a_n2406_n3888# 0.333456f
C49 drain_left.t7 a_n2406_n3888# 0.507454f
C50 drain_left.t14 a_n2406_n3888# 0.507454f
C51 drain_left.n16 a_n2406_n3888# 3.37235f
C52 drain_left.n17 a_n2406_n3888# 0.333456f
C53 drain_left.t5 a_n2406_n3888# 0.507454f
C54 drain_left.t8 a_n2406_n3888# 0.507454f
C55 drain_left.n18 a_n2406_n3888# 3.37235f
C56 drain_left.n19 a_n2406_n3888# 0.333456f
C57 drain_left.t11 a_n2406_n3888# 0.507454f
C58 drain_left.t1 a_n2406_n3888# 0.507454f
C59 drain_left.n20 a_n2406_n3888# 3.37234f
C60 drain_left.n21 a_n2406_n3888# 0.569426f
C61 plus.n0 a_n2406_n3888# 0.052312f
C62 plus.t12 a_n2406_n3888# 0.332054f
C63 plus.t15 a_n2406_n3888# 0.332054f
C64 plus.n1 a_n2406_n3888# 0.021385f
C65 plus.n2 a_n2406_n3888# 0.052312f
C66 plus.t9 a_n2406_n3888# 0.332054f
C67 plus.t16 a_n2406_n3888# 0.332054f
C68 plus.n3 a_n2406_n3888# 0.019772f
C69 plus.n4 a_n2406_n3888# 0.052312f
C70 plus.t23 a_n2406_n3888# 0.332054f
C71 plus.t13 a_n2406_n3888# 0.332054f
C72 plus.n5 a_n2406_n3888# 0.01816f
C73 plus.t10 a_n2406_n3888# 0.334454f
C74 plus.n6 a_n2406_n3888# 0.154665f
C75 plus.t20 a_n2406_n3888# 0.332054f
C76 plus.n7 a_n2406_n3888# 0.135607f
C77 plus.t17 a_n2406_n3888# 0.332054f
C78 plus.n8 a_n2406_n3888# 0.135607f
C79 plus.n9 a_n2406_n3888# 0.022191f
C80 plus.n10 a_n2406_n3888# 0.114227f
C81 plus.n11 a_n2406_n3888# 0.052312f
C82 plus.n12 a_n2406_n3888# 0.052312f
C83 plus.n13 a_n2406_n3888# 0.021385f
C84 plus.n14 a_n2406_n3888# 0.135607f
C85 plus.n15 a_n2406_n3888# 0.022191f
C86 plus.n16 a_n2406_n3888# 0.135607f
C87 plus.t19 a_n2406_n3888# 0.332054f
C88 plus.n17 a_n2406_n3888# 0.135607f
C89 plus.n18 a_n2406_n3888# 0.022191f
C90 plus.n19 a_n2406_n3888# 0.052312f
C91 plus.n20 a_n2406_n3888# 0.052312f
C92 plus.n21 a_n2406_n3888# 0.052312f
C93 plus.n22 a_n2406_n3888# 0.019772f
C94 plus.n23 a_n2406_n3888# 0.135607f
C95 plus.n24 a_n2406_n3888# 0.022191f
C96 plus.n25 a_n2406_n3888# 0.135607f
C97 plus.t18 a_n2406_n3888# 0.332054f
C98 plus.n26 a_n2406_n3888# 0.135607f
C99 plus.n27 a_n2406_n3888# 0.022191f
C100 plus.n28 a_n2406_n3888# 0.052312f
C101 plus.n29 a_n2406_n3888# 0.052312f
C102 plus.n30 a_n2406_n3888# 0.052312f
C103 plus.n31 a_n2406_n3888# 0.01816f
C104 plus.n32 a_n2406_n3888# 0.135607f
C105 plus.n33 a_n2406_n3888# 0.022191f
C106 plus.n34 a_n2406_n3888# 0.135607f
C107 plus.t22 a_n2406_n3888# 0.334454f
C108 plus.n35 a_n2406_n3888# 0.154592f
C109 plus.n36 a_n2406_n3888# 0.663918f
C110 plus.n37 a_n2406_n3888# 0.052312f
C111 plus.t6 a_n2406_n3888# 0.334454f
C112 plus.t2 a_n2406_n3888# 0.332054f
C113 plus.t0 a_n2406_n3888# 0.332054f
C114 plus.n38 a_n2406_n3888# 0.021385f
C115 plus.n39 a_n2406_n3888# 0.052312f
C116 plus.t8 a_n2406_n3888# 0.332054f
C117 plus.n40 a_n2406_n3888# 0.135607f
C118 plus.t5 a_n2406_n3888# 0.332054f
C119 plus.t4 a_n2406_n3888# 0.332054f
C120 plus.n41 a_n2406_n3888# 0.019772f
C121 plus.n42 a_n2406_n3888# 0.052312f
C122 plus.t1 a_n2406_n3888# 0.332054f
C123 plus.n43 a_n2406_n3888# 0.135607f
C124 plus.t14 a_n2406_n3888# 0.332054f
C125 plus.t7 a_n2406_n3888# 0.332054f
C126 plus.n44 a_n2406_n3888# 0.01816f
C127 plus.t11 a_n2406_n3888# 0.334454f
C128 plus.n45 a_n2406_n3888# 0.154665f
C129 plus.t3 a_n2406_n3888# 0.332054f
C130 plus.n46 a_n2406_n3888# 0.135607f
C131 plus.t21 a_n2406_n3888# 0.332054f
C132 plus.n47 a_n2406_n3888# 0.135607f
C133 plus.n48 a_n2406_n3888# 0.022191f
C134 plus.n49 a_n2406_n3888# 0.114227f
C135 plus.n50 a_n2406_n3888# 0.052312f
C136 plus.n51 a_n2406_n3888# 0.052312f
C137 plus.n52 a_n2406_n3888# 0.021385f
C138 plus.n53 a_n2406_n3888# 0.135607f
C139 plus.n54 a_n2406_n3888# 0.022191f
C140 plus.n55 a_n2406_n3888# 0.135607f
C141 plus.n56 a_n2406_n3888# 0.022191f
C142 plus.n57 a_n2406_n3888# 0.052312f
C143 plus.n58 a_n2406_n3888# 0.052312f
C144 plus.n59 a_n2406_n3888# 0.052312f
C145 plus.n60 a_n2406_n3888# 0.019772f
C146 plus.n61 a_n2406_n3888# 0.135607f
C147 plus.n62 a_n2406_n3888# 0.022191f
C148 plus.n63 a_n2406_n3888# 0.135607f
C149 plus.n64 a_n2406_n3888# 0.022191f
C150 plus.n65 a_n2406_n3888# 0.052312f
C151 plus.n66 a_n2406_n3888# 0.052312f
C152 plus.n67 a_n2406_n3888# 0.052312f
C153 plus.n68 a_n2406_n3888# 0.01816f
C154 plus.n69 a_n2406_n3888# 0.135607f
C155 plus.n70 a_n2406_n3888# 0.022191f
C156 plus.n71 a_n2406_n3888# 0.135607f
C157 plus.n72 a_n2406_n3888# 0.154592f
C158 plus.n73 a_n2406_n3888# 1.82095f
C159 source.t7 a_n2406_n3888# 3.59771f
C160 source.n0 a_n2406_n3888# 1.60161f
C161 source.t12 a_n2406_n3888# 0.451832f
C162 source.t13 a_n2406_n3888# 0.451832f
C163 source.n1 a_n2406_n3888# 2.92676f
C164 source.n2 a_n2406_n3888# 0.338658f
C165 source.t8 a_n2406_n3888# 0.451832f
C166 source.t22 a_n2406_n3888# 0.451832f
C167 source.n3 a_n2406_n3888# 2.92676f
C168 source.n4 a_n2406_n3888# 0.338658f
C169 source.t4 a_n2406_n3888# 0.451832f
C170 source.t17 a_n2406_n3888# 0.451832f
C171 source.n5 a_n2406_n3888# 2.92676f
C172 source.n6 a_n2406_n3888# 0.338658f
C173 source.t18 a_n2406_n3888# 0.451832f
C174 source.t14 a_n2406_n3888# 0.451832f
C175 source.n7 a_n2406_n3888# 2.92676f
C176 source.n8 a_n2406_n3888# 0.338658f
C177 source.t9 a_n2406_n3888# 0.451832f
C178 source.t21 a_n2406_n3888# 0.451832f
C179 source.n9 a_n2406_n3888# 2.92676f
C180 source.n10 a_n2406_n3888# 0.338658f
C181 source.t2 a_n2406_n3888# 3.59771f
C182 source.n11 a_n2406_n3888# 0.473666f
C183 source.t41 a_n2406_n3888# 3.59771f
C184 source.n12 a_n2406_n3888# 0.473666f
C185 source.t35 a_n2406_n3888# 0.451832f
C186 source.t42 a_n2406_n3888# 0.451832f
C187 source.n13 a_n2406_n3888# 2.92676f
C188 source.n14 a_n2406_n3888# 0.338658f
C189 source.t40 a_n2406_n3888# 0.451832f
C190 source.t38 a_n2406_n3888# 0.451832f
C191 source.n15 a_n2406_n3888# 2.92676f
C192 source.n16 a_n2406_n3888# 0.338658f
C193 source.t34 a_n2406_n3888# 0.451832f
C194 source.t30 a_n2406_n3888# 0.451832f
C195 source.n17 a_n2406_n3888# 2.92676f
C196 source.n18 a_n2406_n3888# 0.338658f
C197 source.t36 a_n2406_n3888# 0.451832f
C198 source.t32 a_n2406_n3888# 0.451832f
C199 source.n19 a_n2406_n3888# 2.92676f
C200 source.n20 a_n2406_n3888# 0.338658f
C201 source.t28 a_n2406_n3888# 0.451832f
C202 source.t26 a_n2406_n3888# 0.451832f
C203 source.n21 a_n2406_n3888# 2.92676f
C204 source.n22 a_n2406_n3888# 0.338658f
C205 source.t31 a_n2406_n3888# 3.59771f
C206 source.n23 a_n2406_n3888# 2.02043f
C207 source.t5 a_n2406_n3888# 3.59771f
C208 source.n24 a_n2406_n3888# 2.02043f
C209 source.t19 a_n2406_n3888# 0.451832f
C210 source.t0 a_n2406_n3888# 0.451832f
C211 source.n25 a_n2406_n3888# 2.92676f
C212 source.n26 a_n2406_n3888# 0.338661f
C213 source.t11 a_n2406_n3888# 0.451832f
C214 source.t1 a_n2406_n3888# 0.451832f
C215 source.n27 a_n2406_n3888# 2.92676f
C216 source.n28 a_n2406_n3888# 0.338661f
C217 source.t16 a_n2406_n3888# 0.451832f
C218 source.t15 a_n2406_n3888# 0.451832f
C219 source.n29 a_n2406_n3888# 2.92676f
C220 source.n30 a_n2406_n3888# 0.338661f
C221 source.t20 a_n2406_n3888# 0.451832f
C222 source.t6 a_n2406_n3888# 0.451832f
C223 source.n31 a_n2406_n3888# 2.92676f
C224 source.n32 a_n2406_n3888# 0.338661f
C225 source.t23 a_n2406_n3888# 0.451832f
C226 source.t3 a_n2406_n3888# 0.451832f
C227 source.n33 a_n2406_n3888# 2.92676f
C228 source.n34 a_n2406_n3888# 0.338661f
C229 source.t10 a_n2406_n3888# 3.59771f
C230 source.n35 a_n2406_n3888# 0.47367f
C231 source.t43 a_n2406_n3888# 3.59771f
C232 source.n36 a_n2406_n3888# 0.47367f
C233 source.t29 a_n2406_n3888# 0.451832f
C234 source.t24 a_n2406_n3888# 0.451832f
C235 source.n37 a_n2406_n3888# 2.92676f
C236 source.n38 a_n2406_n3888# 0.338661f
C237 source.t45 a_n2406_n3888# 0.451832f
C238 source.t37 a_n2406_n3888# 0.451832f
C239 source.n39 a_n2406_n3888# 2.92676f
C240 source.n40 a_n2406_n3888# 0.338661f
C241 source.t27 a_n2406_n3888# 0.451832f
C242 source.t47 a_n2406_n3888# 0.451832f
C243 source.n41 a_n2406_n3888# 2.92676f
C244 source.n42 a_n2406_n3888# 0.338661f
C245 source.t44 a_n2406_n3888# 0.451832f
C246 source.t33 a_n2406_n3888# 0.451832f
C247 source.n43 a_n2406_n3888# 2.92676f
C248 source.n44 a_n2406_n3888# 0.338661f
C249 source.t25 a_n2406_n3888# 0.451832f
C250 source.t46 a_n2406_n3888# 0.451832f
C251 source.n45 a_n2406_n3888# 2.92676f
C252 source.n46 a_n2406_n3888# 0.338661f
C253 source.t39 a_n2406_n3888# 3.59771f
C254 source.n47 a_n2406_n3888# 0.616803f
C255 source.n48 a_n2406_n3888# 1.84034f
C256 drain_right.t23 a_n2406_n3888# 0.506719f
C257 drain_right.t3 a_n2406_n3888# 0.506719f
C258 drain_right.n0 a_n2406_n3888# 3.37061f
C259 drain_right.t20 a_n2406_n3888# 0.506719f
C260 drain_right.t17 a_n2406_n3888# 0.506719f
C261 drain_right.n1 a_n2406_n3888# 3.36747f
C262 drain_right.n2 a_n2406_n3888# 0.674174f
C263 drain_right.t15 a_n2406_n3888# 0.506719f
C264 drain_right.t11 a_n2406_n3888# 0.506719f
C265 drain_right.n3 a_n2406_n3888# 3.36747f
C266 drain_right.n4 a_n2406_n3888# 0.305382f
C267 drain_right.t12 a_n2406_n3888# 0.506719f
C268 drain_right.t1 a_n2406_n3888# 0.506719f
C269 drain_right.n5 a_n2406_n3888# 3.37061f
C270 drain_right.t7 a_n2406_n3888# 0.506719f
C271 drain_right.t21 a_n2406_n3888# 0.506719f
C272 drain_right.n6 a_n2406_n3888# 3.36747f
C273 drain_right.n7 a_n2406_n3888# 0.674174f
C274 drain_right.t13 a_n2406_n3888# 0.506719f
C275 drain_right.t16 a_n2406_n3888# 0.506719f
C276 drain_right.n8 a_n2406_n3888# 3.36747f
C277 drain_right.n9 a_n2406_n3888# 0.305382f
C278 drain_right.n10 a_n2406_n3888# 1.69058f
C279 drain_right.t22 a_n2406_n3888# 0.506719f
C280 drain_right.t19 a_n2406_n3888# 0.506719f
C281 drain_right.n11 a_n2406_n3888# 3.3706f
C282 drain_right.t0 a_n2406_n3888# 0.506719f
C283 drain_right.t5 a_n2406_n3888# 0.506719f
C284 drain_right.n12 a_n2406_n3888# 3.36747f
C285 drain_right.n13 a_n2406_n3888# 0.67418f
C286 drain_right.t8 a_n2406_n3888# 0.506719f
C287 drain_right.t18 a_n2406_n3888# 0.506719f
C288 drain_right.n14 a_n2406_n3888# 3.36747f
C289 drain_right.n15 a_n2406_n3888# 0.332973f
C290 drain_right.t6 a_n2406_n3888# 0.506719f
C291 drain_right.t4 a_n2406_n3888# 0.506719f
C292 drain_right.n16 a_n2406_n3888# 3.36747f
C293 drain_right.n17 a_n2406_n3888# 0.332973f
C294 drain_right.t10 a_n2406_n3888# 0.506719f
C295 drain_right.t14 a_n2406_n3888# 0.506719f
C296 drain_right.n18 a_n2406_n3888# 3.36747f
C297 drain_right.n19 a_n2406_n3888# 0.332973f
C298 drain_right.t9 a_n2406_n3888# 0.506719f
C299 drain_right.t2 a_n2406_n3888# 0.506719f
C300 drain_right.n20 a_n2406_n3888# 3.36747f
C301 drain_right.n21 a_n2406_n3888# 0.56859f
C302 minus.n0 a_n2406_n3888# 0.051443f
C303 minus.t16 a_n2406_n3888# 0.328898f
C304 minus.t19 a_n2406_n3888# 0.326538f
C305 minus.t21 a_n2406_n3888# 0.326538f
C306 minus.n1 a_n2406_n3888# 0.02103f
C307 minus.n2 a_n2406_n3888# 0.051443f
C308 minus.t11 a_n2406_n3888# 0.326538f
C309 minus.n3 a_n2406_n3888# 0.133354f
C310 minus.t15 a_n2406_n3888# 0.326538f
C311 minus.t13 a_n2406_n3888# 0.326538f
C312 minus.n4 a_n2406_n3888# 0.019444f
C313 minus.n5 a_n2406_n3888# 0.051443f
C314 minus.t17 a_n2406_n3888# 0.326538f
C315 minus.n6 a_n2406_n3888# 0.133354f
C316 minus.t7 a_n2406_n3888# 0.326538f
C317 minus.t9 a_n2406_n3888# 0.326538f
C318 minus.n7 a_n2406_n3888# 0.017858f
C319 minus.t6 a_n2406_n3888# 0.328898f
C320 minus.n8 a_n2406_n3888# 0.152096f
C321 minus.t12 a_n2406_n3888# 0.326538f
C322 minus.n9 a_n2406_n3888# 0.133354f
C323 minus.t5 a_n2406_n3888# 0.326538f
C324 minus.n10 a_n2406_n3888# 0.133354f
C325 minus.n11 a_n2406_n3888# 0.021823f
C326 minus.n12 a_n2406_n3888# 0.112329f
C327 minus.n13 a_n2406_n3888# 0.051443f
C328 minus.n14 a_n2406_n3888# 0.051443f
C329 minus.n15 a_n2406_n3888# 0.02103f
C330 minus.n16 a_n2406_n3888# 0.133354f
C331 minus.n17 a_n2406_n3888# 0.021823f
C332 minus.n18 a_n2406_n3888# 0.133354f
C333 minus.n19 a_n2406_n3888# 0.021823f
C334 minus.n20 a_n2406_n3888# 0.051443f
C335 minus.n21 a_n2406_n3888# 0.051443f
C336 minus.n22 a_n2406_n3888# 0.051443f
C337 minus.n23 a_n2406_n3888# 0.019444f
C338 minus.n24 a_n2406_n3888# 0.133354f
C339 minus.n25 a_n2406_n3888# 0.021823f
C340 minus.n26 a_n2406_n3888# 0.133354f
C341 minus.n27 a_n2406_n3888# 0.021823f
C342 minus.n28 a_n2406_n3888# 0.051443f
C343 minus.n29 a_n2406_n3888# 0.051443f
C344 minus.n30 a_n2406_n3888# 0.051443f
C345 minus.n31 a_n2406_n3888# 0.017858f
C346 minus.n32 a_n2406_n3888# 0.133354f
C347 minus.n33 a_n2406_n3888# 0.021823f
C348 minus.n34 a_n2406_n3888# 0.133354f
C349 minus.n35 a_n2406_n3888# 0.152024f
C350 minus.n36 a_n2406_n3888# 2.1619f
C351 minus.n37 a_n2406_n3888# 0.051443f
C352 minus.t1 a_n2406_n3888# 0.326538f
C353 minus.t22 a_n2406_n3888# 0.326538f
C354 minus.n38 a_n2406_n3888# 0.02103f
C355 minus.n39 a_n2406_n3888# 0.051443f
C356 minus.t3 a_n2406_n3888# 0.326538f
C357 minus.t0 a_n2406_n3888# 0.326538f
C358 minus.n40 a_n2406_n3888# 0.019444f
C359 minus.n41 a_n2406_n3888# 0.051443f
C360 minus.t10 a_n2406_n3888# 0.326538f
C361 minus.t2 a_n2406_n3888# 0.326538f
C362 minus.n42 a_n2406_n3888# 0.017858f
C363 minus.t4 a_n2406_n3888# 0.328898f
C364 minus.n43 a_n2406_n3888# 0.152096f
C365 minus.t18 a_n2406_n3888# 0.326538f
C366 minus.n44 a_n2406_n3888# 0.133354f
C367 minus.t23 a_n2406_n3888# 0.326538f
C368 minus.n45 a_n2406_n3888# 0.133354f
C369 minus.n46 a_n2406_n3888# 0.021823f
C370 minus.n47 a_n2406_n3888# 0.112329f
C371 minus.n48 a_n2406_n3888# 0.051443f
C372 minus.n49 a_n2406_n3888# 0.051443f
C373 minus.n50 a_n2406_n3888# 0.02103f
C374 minus.n51 a_n2406_n3888# 0.133354f
C375 minus.n52 a_n2406_n3888# 0.021823f
C376 minus.n53 a_n2406_n3888# 0.133354f
C377 minus.t20 a_n2406_n3888# 0.326538f
C378 minus.n54 a_n2406_n3888# 0.133354f
C379 minus.n55 a_n2406_n3888# 0.021823f
C380 minus.n56 a_n2406_n3888# 0.051443f
C381 minus.n57 a_n2406_n3888# 0.051443f
C382 minus.n58 a_n2406_n3888# 0.051443f
C383 minus.n59 a_n2406_n3888# 0.019444f
C384 minus.n60 a_n2406_n3888# 0.133354f
C385 minus.n61 a_n2406_n3888# 0.021823f
C386 minus.n62 a_n2406_n3888# 0.133354f
C387 minus.t14 a_n2406_n3888# 0.326538f
C388 minus.n63 a_n2406_n3888# 0.133354f
C389 minus.n64 a_n2406_n3888# 0.021823f
C390 minus.n65 a_n2406_n3888# 0.051443f
C391 minus.n66 a_n2406_n3888# 0.051443f
C392 minus.n67 a_n2406_n3888# 0.051443f
C393 minus.n68 a_n2406_n3888# 0.017858f
C394 minus.n69 a_n2406_n3888# 0.133354f
C395 minus.n70 a_n2406_n3888# 0.021823f
C396 minus.n71 a_n2406_n3888# 0.133354f
C397 minus.t8 a_n2406_n3888# 0.328898f
C398 minus.n72 a_n2406_n3888# 0.152024f
C399 minus.n73 a_n2406_n3888# 0.339132f
C400 minus.n74 a_n2406_n3888# 2.59192f
.ends

