* NGSPICE file created from diffpair586.ext - technology: sky130A

.subckt diffpair586 minus drain_right drain_left source plus
X0 source.t27 plus.t0 drain_left.t4 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X1 source.t26 plus.t1 drain_left.t13 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X2 drain_left.t12 plus.t2 source.t25 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X3 source.t6 minus.t0 drain_right.t13 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X4 source.t8 minus.t1 drain_right.t12 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X5 drain_right.t11 minus.t2 source.t2 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X6 source.t0 minus.t3 drain_right.t10 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X7 source.t24 plus.t3 drain_left.t6 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X8 a_n1644_n4888# a_n1644_n4888# a_n1644_n4888# a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.25
X9 drain_left.t5 plus.t4 source.t23 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X10 source.t1 minus.t4 drain_right.t9 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X11 source.t3 minus.t5 drain_right.t8 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X12 drain_left.t11 plus.t5 source.t22 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X13 drain_right.t7 minus.t6 source.t10 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X14 drain_left.t9 plus.t6 source.t21 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X15 drain_left.t8 plus.t7 source.t20 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X16 drain_left.t7 plus.t8 source.t19 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X17 drain_left.t1 plus.t9 source.t18 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X18 drain_right.t6 minus.t7 source.t5 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X19 drain_right.t5 minus.t8 source.t12 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X20 a_n1644_n4888# a_n1644_n4888# a_n1644_n4888# a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X21 a_n1644_n4888# a_n1644_n4888# a_n1644_n4888# a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X22 source.t13 minus.t9 drain_right.t4 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X23 drain_left.t3 plus.t10 source.t17 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X24 drain_right.t3 minus.t10 source.t4 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X25 drain_right.t2 minus.t11 source.t9 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.25
X26 source.t16 plus.t11 drain_left.t2 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X27 drain_right.t1 minus.t12 source.t11 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.25
X28 drain_right.t0 minus.t13 source.t7 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X29 source.t15 plus.t12 drain_left.t10 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
X30 a_n1644_n4888# a_n1644_n4888# a_n1644_n4888# a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.25
X31 source.t14 plus.t13 drain_left.t0 a_n1644_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.25
R0 plus.n3 plus.t4 2088.37
R1 plus.n15 plus.t6 2088.37
R2 plus.n20 plus.t2 2088.37
R3 plus.n32 plus.t10 2088.37
R4 plus.n1 plus.t0 2053.32
R5 plus.n4 plus.t1 2053.32
R6 plus.n6 plus.t8 2053.32
R7 plus.n12 plus.t7 2053.32
R8 plus.n14 plus.t12 2053.32
R9 plus.n18 plus.t3 2053.32
R10 plus.n21 plus.t11 2053.32
R11 plus.n23 plus.t9 2053.32
R12 plus.n29 plus.t5 2053.32
R13 plus.n31 plus.t13 2053.32
R14 plus.n3 plus.n2 161.489
R15 plus.n20 plus.n19 161.489
R16 plus.n5 plus.n2 161.3
R17 plus.n8 plus.n7 161.3
R18 plus.n9 plus.n1 161.3
R19 plus.n11 plus.n10 161.3
R20 plus.n13 plus.n0 161.3
R21 plus.n16 plus.n15 161.3
R22 plus.n22 plus.n19 161.3
R23 plus.n25 plus.n24 161.3
R24 plus.n26 plus.n18 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n17 161.3
R27 plus.n33 plus.n32 161.3
R28 plus.n7 plus.n1 73.0308
R29 plus.n11 plus.n1 73.0308
R30 plus.n28 plus.n18 73.0308
R31 plus.n24 plus.n18 73.0308
R32 plus.n6 plus.n5 61.346
R33 plus.n13 plus.n12 61.346
R34 plus.n30 plus.n29 61.346
R35 plus.n23 plus.n22 61.346
R36 plus.n4 plus.n3 49.6611
R37 plus.n15 plus.n14 49.6611
R38 plus.n32 plus.n31 49.6611
R39 plus.n21 plus.n20 49.6611
R40 plus plus.n33 32.2111
R41 plus.n5 plus.n4 23.3702
R42 plus.n14 plus.n13 23.3702
R43 plus.n31 plus.n30 23.3702
R44 plus.n22 plus.n21 23.3702
R45 plus plus.n16 15.1255
R46 plus.n7 plus.n6 11.6853
R47 plus.n12 plus.n11 11.6853
R48 plus.n29 plus.n28 11.6853
R49 plus.n24 plus.n23 11.6853
R50 plus.n8 plus.n2 0.189894
R51 plus.n9 plus.n8 0.189894
R52 plus.n10 plus.n9 0.189894
R53 plus.n10 plus.n0 0.189894
R54 plus.n16 plus.n0 0.189894
R55 plus.n33 plus.n17 0.189894
R56 plus.n27 plus.n17 0.189894
R57 plus.n27 plus.n26 0.189894
R58 plus.n26 plus.n25 0.189894
R59 plus.n25 plus.n19 0.189894
R60 drain_left.n7 drain_left.t5 61.3084
R61 drain_left.n1 drain_left.t3 61.3083
R62 drain_left.n4 drain_left.n2 60.3184
R63 drain_left.n11 drain_left.n10 59.8185
R64 drain_left.n9 drain_left.n8 59.8185
R65 drain_left.n7 drain_left.n6 59.8185
R66 drain_left.n4 drain_left.n3 59.8184
R67 drain_left.n1 drain_left.n0 59.8184
R68 drain_left drain_left.n5 36.3027
R69 drain_left drain_left.n11 6.15322
R70 drain_left.n2 drain_left.t2 0.9905
R71 drain_left.n2 drain_left.t12 0.9905
R72 drain_left.n3 drain_left.t6 0.9905
R73 drain_left.n3 drain_left.t1 0.9905
R74 drain_left.n0 drain_left.t0 0.9905
R75 drain_left.n0 drain_left.t11 0.9905
R76 drain_left.n10 drain_left.t10 0.9905
R77 drain_left.n10 drain_left.t9 0.9905
R78 drain_left.n8 drain_left.t4 0.9905
R79 drain_left.n8 drain_left.t8 0.9905
R80 drain_left.n6 drain_left.t13 0.9905
R81 drain_left.n6 drain_left.t7 0.9905
R82 drain_left.n9 drain_left.n7 0.5005
R83 drain_left.n11 drain_left.n9 0.5005
R84 drain_left.n5 drain_left.n1 0.320154
R85 drain_left.n5 drain_left.n4 0.070154
R86 source.n0 source.t21 44.1297
R87 source.n7 source.t12 44.1296
R88 source.n27 source.t11 44.1295
R89 source.n20 source.t25 44.1295
R90 source.n2 source.n1 43.1397
R91 source.n4 source.n3 43.1397
R92 source.n6 source.n5 43.1397
R93 source.n9 source.n8 43.1397
R94 source.n11 source.n10 43.1397
R95 source.n13 source.n12 43.1397
R96 source.n26 source.n25 43.1396
R97 source.n24 source.n23 43.1396
R98 source.n22 source.n21 43.1396
R99 source.n19 source.n18 43.1396
R100 source.n17 source.n16 43.1396
R101 source.n15 source.n14 43.1396
R102 source.n15 source.n13 28.3483
R103 source.n28 source.n0 22.3354
R104 source.n28 source.n27 5.51343
R105 source.n25 source.t10 0.9905
R106 source.n25 source.t6 0.9905
R107 source.n23 source.t7 0.9905
R108 source.n23 source.t13 0.9905
R109 source.n21 source.t2 0.9905
R110 source.n21 source.t1 0.9905
R111 source.n18 source.t18 0.9905
R112 source.n18 source.t16 0.9905
R113 source.n16 source.t22 0.9905
R114 source.n16 source.t24 0.9905
R115 source.n14 source.t17 0.9905
R116 source.n14 source.t14 0.9905
R117 source.n1 source.t20 0.9905
R118 source.n1 source.t15 0.9905
R119 source.n3 source.t19 0.9905
R120 source.n3 source.t27 0.9905
R121 source.n5 source.t23 0.9905
R122 source.n5 source.t26 0.9905
R123 source.n8 source.t5 0.9905
R124 source.n8 source.t0 0.9905
R125 source.n10 source.t4 0.9905
R126 source.n10 source.t8 0.9905
R127 source.n12 source.t9 0.9905
R128 source.n12 source.t3 0.9905
R129 source.n7 source.n6 0.720328
R130 source.n22 source.n20 0.720328
R131 source.n13 source.n11 0.5005
R132 source.n11 source.n9 0.5005
R133 source.n9 source.n7 0.5005
R134 source.n6 source.n4 0.5005
R135 source.n4 source.n2 0.5005
R136 source.n2 source.n0 0.5005
R137 source.n17 source.n15 0.5005
R138 source.n19 source.n17 0.5005
R139 source.n20 source.n19 0.5005
R140 source.n24 source.n22 0.5005
R141 source.n26 source.n24 0.5005
R142 source.n27 source.n26 0.5005
R143 source source.n28 0.188
R144 minus.n15 minus.t11 2088.37
R145 minus.n3 minus.t8 2088.37
R146 minus.n32 minus.t12 2088.37
R147 minus.n20 minus.t2 2088.37
R148 minus.n1 minus.t1 2053.32
R149 minus.n14 minus.t5 2053.32
R150 minus.n12 minus.t10 2053.32
R151 minus.n6 minus.t7 2053.32
R152 minus.n4 minus.t3 2053.32
R153 minus.n18 minus.t9 2053.32
R154 minus.n31 minus.t0 2053.32
R155 minus.n29 minus.t6 2053.32
R156 minus.n23 minus.t13 2053.32
R157 minus.n21 minus.t4 2053.32
R158 minus.n3 minus.n2 161.489
R159 minus.n20 minus.n19 161.489
R160 minus.n16 minus.n15 161.3
R161 minus.n13 minus.n0 161.3
R162 minus.n11 minus.n10 161.3
R163 minus.n9 minus.n1 161.3
R164 minus.n8 minus.n7 161.3
R165 minus.n5 minus.n2 161.3
R166 minus.n33 minus.n32 161.3
R167 minus.n30 minus.n17 161.3
R168 minus.n28 minus.n27 161.3
R169 minus.n26 minus.n18 161.3
R170 minus.n25 minus.n24 161.3
R171 minus.n22 minus.n19 161.3
R172 minus.n11 minus.n1 73.0308
R173 minus.n7 minus.n1 73.0308
R174 minus.n24 minus.n18 73.0308
R175 minus.n28 minus.n18 73.0308
R176 minus.n13 minus.n12 61.346
R177 minus.n6 minus.n5 61.346
R178 minus.n23 minus.n22 61.346
R179 minus.n30 minus.n29 61.346
R180 minus.n15 minus.n14 49.6611
R181 minus.n4 minus.n3 49.6611
R182 minus.n21 minus.n20 49.6611
R183 minus.n32 minus.n31 49.6611
R184 minus.n34 minus.n16 41.3603
R185 minus.n14 minus.n13 23.3702
R186 minus.n5 minus.n4 23.3702
R187 minus.n22 minus.n21 23.3702
R188 minus.n31 minus.n30 23.3702
R189 minus.n12 minus.n11 11.6853
R190 minus.n7 minus.n6 11.6853
R191 minus.n24 minus.n23 11.6853
R192 minus.n29 minus.n28 11.6853
R193 minus.n34 minus.n33 6.45126
R194 minus.n16 minus.n0 0.189894
R195 minus.n10 minus.n0 0.189894
R196 minus.n10 minus.n9 0.189894
R197 minus.n9 minus.n8 0.189894
R198 minus.n8 minus.n2 0.189894
R199 minus.n25 minus.n19 0.189894
R200 minus.n26 minus.n25 0.189894
R201 minus.n27 minus.n26 0.189894
R202 minus.n27 minus.n17 0.189894
R203 minus.n33 minus.n17 0.189894
R204 minus minus.n34 0.188
R205 drain_right.n1 drain_right.t11 61.3083
R206 drain_right.n11 drain_right.t2 60.8084
R207 drain_right.n8 drain_right.n6 60.3185
R208 drain_right.n4 drain_right.n2 60.3184
R209 drain_right.n8 drain_right.n7 59.8185
R210 drain_right.n10 drain_right.n9 59.8185
R211 drain_right.n4 drain_right.n3 59.8184
R212 drain_right.n1 drain_right.n0 59.8184
R213 drain_right drain_right.n5 35.7495
R214 drain_right drain_right.n11 5.90322
R215 drain_right.n2 drain_right.t13 0.9905
R216 drain_right.n2 drain_right.t1 0.9905
R217 drain_right.n3 drain_right.t4 0.9905
R218 drain_right.n3 drain_right.t7 0.9905
R219 drain_right.n0 drain_right.t9 0.9905
R220 drain_right.n0 drain_right.t0 0.9905
R221 drain_right.n6 drain_right.t10 0.9905
R222 drain_right.n6 drain_right.t5 0.9905
R223 drain_right.n7 drain_right.t12 0.9905
R224 drain_right.n7 drain_right.t6 0.9905
R225 drain_right.n9 drain_right.t8 0.9905
R226 drain_right.n9 drain_right.t3 0.9905
R227 drain_right.n11 drain_right.n10 0.5005
R228 drain_right.n10 drain_right.n8 0.5005
R229 drain_right.n5 drain_right.n1 0.320154
R230 drain_right.n5 drain_right.n4 0.070154
C0 source drain_left 48.9652f
C1 drain_right minus 7.41951f
C2 drain_right plus 0.316461f
C3 plus minus 6.68769f
C4 drain_right drain_left 0.84441f
C5 drain_right source 48.9474f
C6 minus drain_left 0.171605f
C7 plus drain_left 7.57303f
C8 minus source 6.6944f
C9 plus source 6.70957f
C10 drain_right a_n1644_n4888# 9.889811f
C11 drain_left a_n1644_n4888# 10.17085f
C12 source a_n1644_n4888# 8.859434f
C13 minus a_n1644_n4888# 6.925898f
C14 plus a_n1644_n4888# 9.498509f
C15 drain_right.t11 a_n1644_n4888# 6.05439f
C16 drain_right.t9 a_n1644_n4888# 0.517499f
C17 drain_right.t0 a_n1644_n4888# 0.517499f
C18 drain_right.n0 a_n1644_n4888# 4.73109f
C19 drain_right.n1 a_n1644_n4888# 0.795475f
C20 drain_right.t13 a_n1644_n4888# 0.517499f
C21 drain_right.t1 a_n1644_n4888# 0.517499f
C22 drain_right.n2 a_n1644_n4888# 4.73437f
C23 drain_right.t4 a_n1644_n4888# 0.517499f
C24 drain_right.t7 a_n1644_n4888# 0.517499f
C25 drain_right.n3 a_n1644_n4888# 4.73109f
C26 drain_right.n4 a_n1644_n4888# 0.73904f
C27 drain_right.n5 a_n1644_n4888# 2.10036f
C28 drain_right.t10 a_n1644_n4888# 0.517499f
C29 drain_right.t5 a_n1644_n4888# 0.517499f
C30 drain_right.n6 a_n1644_n4888# 4.73436f
C31 drain_right.t12 a_n1644_n4888# 0.517499f
C32 drain_right.t6 a_n1644_n4888# 0.517499f
C33 drain_right.n7 a_n1644_n4888# 4.73109f
C34 drain_right.n8 a_n1644_n4888# 0.773559f
C35 drain_right.t8 a_n1644_n4888# 0.517499f
C36 drain_right.t3 a_n1644_n4888# 0.517499f
C37 drain_right.n9 a_n1644_n4888# 4.73109f
C38 drain_right.n10 a_n1644_n4888# 0.381823f
C39 drain_right.t2 a_n1644_n4888# 6.05088f
C40 drain_right.n11 a_n1644_n4888# 0.703478f
C41 minus.n0 a_n1644_n4888# 0.053234f
C42 minus.t11 a_n1644_n4888# 0.754371f
C43 minus.t5 a_n1644_n4888# 0.749656f
C44 minus.t10 a_n1644_n4888# 0.749656f
C45 minus.t1 a_n1644_n4888# 0.749656f
C46 minus.n1 a_n1644_n4888# 0.298874f
C47 minus.n2 a_n1644_n4888# 0.113945f
C48 minus.t7 a_n1644_n4888# 0.749656f
C49 minus.t3 a_n1644_n4888# 0.749656f
C50 minus.t8 a_n1644_n4888# 0.754371f
C51 minus.n3 a_n1644_n4888# 0.296528f
C52 minus.n4 a_n1644_n4888# 0.281214f
C53 minus.n5 a_n1644_n4888# 0.020285f
C54 minus.n6 a_n1644_n4888# 0.281214f
C55 minus.n7 a_n1644_n4888# 0.020285f
C56 minus.n8 a_n1644_n4888# 0.053234f
C57 minus.n9 a_n1644_n4888# 0.053234f
C58 minus.n10 a_n1644_n4888# 0.053234f
C59 minus.n11 a_n1644_n4888# 0.020285f
C60 minus.n12 a_n1644_n4888# 0.281214f
C61 minus.n13 a_n1644_n4888# 0.020285f
C62 minus.n14 a_n1644_n4888# 0.281214f
C63 minus.n15 a_n1644_n4888# 0.296456f
C64 minus.n16 a_n1644_n4888# 2.30294f
C65 minus.n17 a_n1644_n4888# 0.053234f
C66 minus.t0 a_n1644_n4888# 0.749656f
C67 minus.t6 a_n1644_n4888# 0.749656f
C68 minus.t9 a_n1644_n4888# 0.749656f
C69 minus.n18 a_n1644_n4888# 0.298874f
C70 minus.n19 a_n1644_n4888# 0.113945f
C71 minus.t13 a_n1644_n4888# 0.749656f
C72 minus.t4 a_n1644_n4888# 0.749656f
C73 minus.t2 a_n1644_n4888# 0.754371f
C74 minus.n20 a_n1644_n4888# 0.296528f
C75 minus.n21 a_n1644_n4888# 0.281214f
C76 minus.n22 a_n1644_n4888# 0.020285f
C77 minus.n23 a_n1644_n4888# 0.281214f
C78 minus.n24 a_n1644_n4888# 0.020285f
C79 minus.n25 a_n1644_n4888# 0.053234f
C80 minus.n26 a_n1644_n4888# 0.053234f
C81 minus.n27 a_n1644_n4888# 0.053234f
C82 minus.n28 a_n1644_n4888# 0.020285f
C83 minus.n29 a_n1644_n4888# 0.281214f
C84 minus.n30 a_n1644_n4888# 0.020285f
C85 minus.n31 a_n1644_n4888# 0.281214f
C86 minus.t12 a_n1644_n4888# 0.754371f
C87 minus.n32 a_n1644_n4888# 0.296456f
C88 minus.n33 a_n1644_n4888# 0.3419f
C89 minus.n34 a_n1644_n4888# 2.75668f
C90 source.t21 a_n1644_n4888# 6.01025f
C91 source.n0 a_n1644_n4888# 2.54908f
C92 source.t20 a_n1644_n4888# 0.525906f
C93 source.t15 a_n1644_n4888# 0.525906f
C94 source.n1 a_n1644_n4888# 4.70182f
C95 source.n2 a_n1644_n4888# 0.448914f
C96 source.t19 a_n1644_n4888# 0.525906f
C97 source.t27 a_n1644_n4888# 0.525906f
C98 source.n3 a_n1644_n4888# 4.70182f
C99 source.n4 a_n1644_n4888# 0.448914f
C100 source.t23 a_n1644_n4888# 0.525906f
C101 source.t26 a_n1644_n4888# 0.525906f
C102 source.n5 a_n1644_n4888# 4.70182f
C103 source.n6 a_n1644_n4888# 0.472484f
C104 source.t12 a_n1644_n4888# 6.01026f
C105 source.n7 a_n1644_n4888# 0.598331f
C106 source.t5 a_n1644_n4888# 0.525906f
C107 source.t0 a_n1644_n4888# 0.525906f
C108 source.n8 a_n1644_n4888# 4.70182f
C109 source.n9 a_n1644_n4888# 0.448914f
C110 source.t4 a_n1644_n4888# 0.525906f
C111 source.t8 a_n1644_n4888# 0.525906f
C112 source.n10 a_n1644_n4888# 4.70182f
C113 source.n11 a_n1644_n4888# 0.448914f
C114 source.t9 a_n1644_n4888# 0.525906f
C115 source.t3 a_n1644_n4888# 0.525906f
C116 source.n12 a_n1644_n4888# 4.70182f
C117 source.n13 a_n1644_n4888# 3.06456f
C118 source.t17 a_n1644_n4888# 0.525906f
C119 source.t14 a_n1644_n4888# 0.525906f
C120 source.n14 a_n1644_n4888# 4.70183f
C121 source.n15 a_n1644_n4888# 3.06455f
C122 source.t22 a_n1644_n4888# 0.525906f
C123 source.t24 a_n1644_n4888# 0.525906f
C124 source.n16 a_n1644_n4888# 4.70183f
C125 source.n17 a_n1644_n4888# 0.448905f
C126 source.t18 a_n1644_n4888# 0.525906f
C127 source.t16 a_n1644_n4888# 0.525906f
C128 source.n18 a_n1644_n4888# 4.70183f
C129 source.n19 a_n1644_n4888# 0.448905f
C130 source.t25 a_n1644_n4888# 6.01023f
C131 source.n20 a_n1644_n4888# 0.598365f
C132 source.t2 a_n1644_n4888# 0.525906f
C133 source.t1 a_n1644_n4888# 0.525906f
C134 source.n21 a_n1644_n4888# 4.70183f
C135 source.n22 a_n1644_n4888# 0.472475f
C136 source.t7 a_n1644_n4888# 0.525906f
C137 source.t13 a_n1644_n4888# 0.525906f
C138 source.n23 a_n1644_n4888# 4.70183f
C139 source.n24 a_n1644_n4888# 0.448905f
C140 source.t10 a_n1644_n4888# 0.525906f
C141 source.t6 a_n1644_n4888# 0.525906f
C142 source.n25 a_n1644_n4888# 4.70183f
C143 source.n26 a_n1644_n4888# 0.448905f
C144 source.t11 a_n1644_n4888# 6.01023f
C145 source.n27 a_n1644_n4888# 0.7557f
C146 source.n28 a_n1644_n4888# 2.99254f
C147 drain_left.t3 a_n1644_n4888# 6.07284f
C148 drain_left.t0 a_n1644_n4888# 0.519076f
C149 drain_left.t11 a_n1644_n4888# 0.519076f
C150 drain_left.n0 a_n1644_n4888# 4.74551f
C151 drain_left.n1 a_n1644_n4888# 0.797898f
C152 drain_left.t2 a_n1644_n4888# 0.519076f
C153 drain_left.t12 a_n1644_n4888# 0.519076f
C154 drain_left.n2 a_n1644_n4888# 4.74879f
C155 drain_left.t6 a_n1644_n4888# 0.519076f
C156 drain_left.t1 a_n1644_n4888# 0.519076f
C157 drain_left.n3 a_n1644_n4888# 4.74551f
C158 drain_left.n4 a_n1644_n4888# 0.741291f
C159 drain_left.n5 a_n1644_n4888# 2.17532f
C160 drain_left.t5 a_n1644_n4888# 6.07286f
C161 drain_left.t13 a_n1644_n4888# 0.519076f
C162 drain_left.t7 a_n1644_n4888# 0.519076f
C163 drain_left.n6 a_n1644_n4888# 4.7455f
C164 drain_left.n7 a_n1644_n4888# 0.814585f
C165 drain_left.t4 a_n1644_n4888# 0.519076f
C166 drain_left.t8 a_n1644_n4888# 0.519076f
C167 drain_left.n8 a_n1644_n4888# 4.7455f
C168 drain_left.n9 a_n1644_n4888# 0.382986f
C169 drain_left.t10 a_n1644_n4888# 0.519076f
C170 drain_left.t9 a_n1644_n4888# 0.519076f
C171 drain_left.n10 a_n1644_n4888# 4.7455f
C172 drain_left.n11 a_n1644_n4888# 0.654085f
C173 plus.n0 a_n1644_n4888# 0.054025f
C174 plus.t12 a_n1644_n4888# 0.760802f
C175 plus.t7 a_n1644_n4888# 0.760802f
C176 plus.t0 a_n1644_n4888# 0.760802f
C177 plus.n1 a_n1644_n4888# 0.303317f
C178 plus.n2 a_n1644_n4888# 0.115639f
C179 plus.t8 a_n1644_n4888# 0.760802f
C180 plus.t1 a_n1644_n4888# 0.760802f
C181 plus.t4 a_n1644_n4888# 0.765587f
C182 plus.n3 a_n1644_n4888# 0.300936f
C183 plus.n4 a_n1644_n4888# 0.285396f
C184 plus.n5 a_n1644_n4888# 0.020587f
C185 plus.n6 a_n1644_n4888# 0.285396f
C186 plus.n7 a_n1644_n4888# 0.020587f
C187 plus.n8 a_n1644_n4888# 0.054025f
C188 plus.n9 a_n1644_n4888# 0.054025f
C189 plus.n10 a_n1644_n4888# 0.054025f
C190 plus.n11 a_n1644_n4888# 0.020587f
C191 plus.n12 a_n1644_n4888# 0.285396f
C192 plus.n13 a_n1644_n4888# 0.020587f
C193 plus.n14 a_n1644_n4888# 0.285396f
C194 plus.t6 a_n1644_n4888# 0.765587f
C195 plus.n15 a_n1644_n4888# 0.300864f
C196 plus.n16 a_n1644_n4888# 0.814271f
C197 plus.n17 a_n1644_n4888# 0.054025f
C198 plus.t10 a_n1644_n4888# 0.765587f
C199 plus.t13 a_n1644_n4888# 0.760802f
C200 plus.t5 a_n1644_n4888# 0.760802f
C201 plus.t3 a_n1644_n4888# 0.760802f
C202 plus.n18 a_n1644_n4888# 0.303317f
C203 plus.n19 a_n1644_n4888# 0.115639f
C204 plus.t9 a_n1644_n4888# 0.760802f
C205 plus.t11 a_n1644_n4888# 0.760802f
C206 plus.t2 a_n1644_n4888# 0.765587f
C207 plus.n20 a_n1644_n4888# 0.300936f
C208 plus.n21 a_n1644_n4888# 0.285396f
C209 plus.n22 a_n1644_n4888# 0.020587f
C210 plus.n23 a_n1644_n4888# 0.285396f
C211 plus.n24 a_n1644_n4888# 0.020587f
C212 plus.n25 a_n1644_n4888# 0.054025f
C213 plus.n26 a_n1644_n4888# 0.054025f
C214 plus.n27 a_n1644_n4888# 0.054025f
C215 plus.n28 a_n1644_n4888# 0.020587f
C216 plus.n29 a_n1644_n4888# 0.285396f
C217 plus.n30 a_n1644_n4888# 0.020587f
C218 plus.n31 a_n1644_n4888# 0.285396f
C219 plus.n32 a_n1644_n4888# 0.300864f
C220 plus.n33 a_n1644_n4888# 1.84201f
.ends

