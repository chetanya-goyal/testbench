* NGSPICE file created from diffpair129.ext - technology: sky130A

.subckt diffpair129 minus drain_right drain_left source plus
X0 drain_right.t23 minus.t0 source.t34 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X1 a_n2874_n1288# a_n2874_n1288# a_n2874_n1288# a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.5
X2 drain_right.t22 minus.t1 source.t31 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X3 drain_right.t21 minus.t2 source.t33 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X4 drain_left.t23 plus.t0 source.t11 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X5 source.t15 plus.t1 drain_left.t22 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X6 source.t32 minus.t3 drain_right.t20 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X7 source.t19 plus.t2 drain_left.t21 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X8 source.t10 plus.t3 drain_left.t20 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X9 source.t23 minus.t4 drain_right.t19 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X10 source.t14 plus.t4 drain_left.t19 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X11 source.t20 plus.t5 drain_left.t18 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X12 source.t39 minus.t5 drain_right.t18 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X13 source.t21 plus.t6 drain_left.t17 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X14 source.t30 minus.t6 drain_right.t17 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X15 drain_left.t16 plus.t7 source.t2 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X16 drain_right.t16 minus.t7 source.t27 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X17 drain_right.t15 minus.t8 source.t36 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X18 source.t37 minus.t9 drain_right.t14 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X19 drain_left.t15 plus.t8 source.t7 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X20 drain_left.t14 plus.t9 source.t1 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X21 drain_left.t13 plus.t10 source.t5 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X22 source.t12 plus.t11 drain_left.t12 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X23 source.t16 plus.t12 drain_left.t11 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X24 source.t24 minus.t10 drain_right.t13 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X25 source.t38 minus.t11 drain_right.t12 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X26 drain_right.t11 minus.t12 source.t43 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X27 source.t17 plus.t13 drain_left.t10 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X28 a_n2874_n1288# a_n2874_n1288# a_n2874_n1288# a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X29 a_n2874_n1288# a_n2874_n1288# a_n2874_n1288# a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X30 drain_left.t9 plus.t14 source.t8 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X31 drain_right.t10 minus.t13 source.t44 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X32 drain_right.t9 minus.t14 source.t42 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X33 a_n2874_n1288# a_n2874_n1288# a_n2874_n1288# a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X34 drain_right.t8 minus.t15 source.t45 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X35 source.t46 plus.t15 drain_left.t8 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X36 drain_left.t7 plus.t16 source.t47 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X37 drain_right.t7 minus.t16 source.t35 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X38 source.t41 minus.t17 drain_right.t6 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X39 drain_right.t5 minus.t18 source.t28 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X40 source.t22 minus.t19 drain_right.t4 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X41 drain_left.t6 plus.t17 source.t4 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X42 source.t26 minus.t20 drain_right.t3 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X43 source.t0 plus.t18 drain_left.t5 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X44 source.t29 minus.t21 drain_right.t2 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X45 drain_right.t1 minus.t22 source.t25 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X46 drain_left.t4 plus.t19 source.t3 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X47 source.t18 plus.t20 drain_left.t3 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X48 drain_left.t2 plus.t21 source.t9 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X49 source.t40 minus.t23 drain_right.t0 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X50 drain_left.t1 plus.t22 source.t6 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X51 drain_left.t0 plus.t23 source.t13 a_n2874_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
R0 minus.n9 minus.t13 201.325
R1 minus.n43 minus.t20 201.325
R2 minus.n8 minus.t4 174.966
R3 minus.n7 minus.t8 174.966
R4 minus.n13 minus.t19 174.966
R5 minus.n5 minus.t7 174.966
R6 minus.n18 minus.t10 174.966
R7 minus.n20 minus.t1 174.966
R8 minus.n3 minus.t11 174.966
R9 minus.n25 minus.t16 174.966
R10 minus.n1 minus.t5 174.966
R11 minus.n30 minus.t14 174.966
R12 minus.n32 minus.t21 174.966
R13 minus.n42 minus.t0 174.966
R14 minus.n41 minus.t17 174.966
R15 minus.n47 minus.t22 174.966
R16 minus.n39 minus.t9 174.966
R17 minus.n52 minus.t2 174.966
R18 minus.n54 minus.t6 174.966
R19 minus.n37 minus.t15 174.966
R20 minus.n59 minus.t3 174.966
R21 minus.n35 minus.t12 174.966
R22 minus.n64 minus.t23 174.966
R23 minus.n66 minus.t18 174.966
R24 minus.n33 minus.n32 161.3
R25 minus.n31 minus.n0 161.3
R26 minus.n30 minus.n29 161.3
R27 minus.n28 minus.n1 161.3
R28 minus.n27 minus.n26 161.3
R29 minus.n25 minus.n2 161.3
R30 minus.n24 minus.n23 161.3
R31 minus.n22 minus.n3 161.3
R32 minus.n21 minus.n20 161.3
R33 minus.n19 minus.n4 161.3
R34 minus.n18 minus.n17 161.3
R35 minus.n16 minus.n5 161.3
R36 minus.n15 minus.n14 161.3
R37 minus.n13 minus.n6 161.3
R38 minus.n12 minus.n11 161.3
R39 minus.n10 minus.n7 161.3
R40 minus.n67 minus.n66 161.3
R41 minus.n65 minus.n34 161.3
R42 minus.n64 minus.n63 161.3
R43 minus.n62 minus.n35 161.3
R44 minus.n61 minus.n60 161.3
R45 minus.n59 minus.n36 161.3
R46 minus.n58 minus.n57 161.3
R47 minus.n56 minus.n37 161.3
R48 minus.n55 minus.n54 161.3
R49 minus.n53 minus.n38 161.3
R50 minus.n52 minus.n51 161.3
R51 minus.n50 minus.n39 161.3
R52 minus.n49 minus.n48 161.3
R53 minus.n47 minus.n40 161.3
R54 minus.n46 minus.n45 161.3
R55 minus.n44 minus.n41 161.3
R56 minus.n8 minus.n7 48.2005
R57 minus.n18 minus.n5 48.2005
R58 minus.n20 minus.n3 48.2005
R59 minus.n30 minus.n1 48.2005
R60 minus.n42 minus.n41 48.2005
R61 minus.n52 minus.n39 48.2005
R62 minus.n54 minus.n37 48.2005
R63 minus.n64 minus.n35 48.2005
R64 minus.n14 minus.n13 47.4702
R65 minus.n25 minus.n24 47.4702
R66 minus.n48 minus.n47 47.4702
R67 minus.n59 minus.n58 47.4702
R68 minus.n32 minus.n31 46.0096
R69 minus.n66 minus.n65 46.0096
R70 minus.n10 minus.n9 45.0871
R71 minus.n44 minus.n43 45.0871
R72 minus.n68 minus.n33 32.4588
R73 minus.n13 minus.n12 25.5611
R74 minus.n26 minus.n25 25.5611
R75 minus.n47 minus.n46 25.5611
R76 minus.n60 minus.n59 25.5611
R77 minus.n20 minus.n19 24.1005
R78 minus.n19 minus.n18 24.1005
R79 minus.n53 minus.n52 24.1005
R80 minus.n54 minus.n53 24.1005
R81 minus.n12 minus.n7 22.6399
R82 minus.n26 minus.n1 22.6399
R83 minus.n46 minus.n41 22.6399
R84 minus.n60 minus.n35 22.6399
R85 minus.n9 minus.n8 14.1472
R86 minus.n43 minus.n42 14.1472
R87 minus.n68 minus.n67 6.52702
R88 minus.n31 minus.n30 2.19141
R89 minus.n65 minus.n64 2.19141
R90 minus.n14 minus.n5 0.730803
R91 minus.n24 minus.n3 0.730803
R92 minus.n48 minus.n39 0.730803
R93 minus.n58 minus.n37 0.730803
R94 minus.n33 minus.n0 0.189894
R95 minus.n29 minus.n0 0.189894
R96 minus.n29 minus.n28 0.189894
R97 minus.n28 minus.n27 0.189894
R98 minus.n27 minus.n2 0.189894
R99 minus.n23 minus.n2 0.189894
R100 minus.n23 minus.n22 0.189894
R101 minus.n22 minus.n21 0.189894
R102 minus.n21 minus.n4 0.189894
R103 minus.n17 minus.n4 0.189894
R104 minus.n17 minus.n16 0.189894
R105 minus.n16 minus.n15 0.189894
R106 minus.n15 minus.n6 0.189894
R107 minus.n11 minus.n6 0.189894
R108 minus.n11 minus.n10 0.189894
R109 minus.n45 minus.n44 0.189894
R110 minus.n45 minus.n40 0.189894
R111 minus.n49 minus.n40 0.189894
R112 minus.n50 minus.n49 0.189894
R113 minus.n51 minus.n50 0.189894
R114 minus.n51 minus.n38 0.189894
R115 minus.n55 minus.n38 0.189894
R116 minus.n56 minus.n55 0.189894
R117 minus.n57 minus.n56 0.189894
R118 minus.n57 minus.n36 0.189894
R119 minus.n61 minus.n36 0.189894
R120 minus.n62 minus.n61 0.189894
R121 minus.n63 minus.n62 0.189894
R122 minus.n63 minus.n34 0.189894
R123 minus.n67 minus.n34 0.189894
R124 minus minus.n68 0.188
R125 source.n98 source.n96 289.615
R126 source.n80 source.n78 289.615
R127 source.n72 source.n70 289.615
R128 source.n54 source.n52 289.615
R129 source.n2 source.n0 289.615
R130 source.n20 source.n18 289.615
R131 source.n28 source.n26 289.615
R132 source.n46 source.n44 289.615
R133 source.n99 source.n98 185
R134 source.n81 source.n80 185
R135 source.n73 source.n72 185
R136 source.n55 source.n54 185
R137 source.n3 source.n2 185
R138 source.n21 source.n20 185
R139 source.n29 source.n28 185
R140 source.n47 source.n46 185
R141 source.t28 source.n97 167.117
R142 source.t26 source.n79 167.117
R143 source.t9 source.n71 167.117
R144 source.t12 source.n53 167.117
R145 source.t11 source.n1 167.117
R146 source.t20 source.n19 167.117
R147 source.t44 source.n27 167.117
R148 source.t29 source.n45 167.117
R149 source.n9 source.n8 84.1169
R150 source.n11 source.n10 84.1169
R151 source.n13 source.n12 84.1169
R152 source.n15 source.n14 84.1169
R153 source.n17 source.n16 84.1169
R154 source.n35 source.n34 84.1169
R155 source.n37 source.n36 84.1169
R156 source.n39 source.n38 84.1169
R157 source.n41 source.n40 84.1169
R158 source.n43 source.n42 84.1169
R159 source.n95 source.n94 84.1168
R160 source.n93 source.n92 84.1168
R161 source.n91 source.n90 84.1168
R162 source.n89 source.n88 84.1168
R163 source.n87 source.n86 84.1168
R164 source.n69 source.n68 84.1168
R165 source.n67 source.n66 84.1168
R166 source.n65 source.n64 84.1168
R167 source.n63 source.n62 84.1168
R168 source.n61 source.n60 84.1168
R169 source.n98 source.t28 52.3082
R170 source.n80 source.t26 52.3082
R171 source.n72 source.t9 52.3082
R172 source.n54 source.t12 52.3082
R173 source.n2 source.t11 52.3082
R174 source.n20 source.t20 52.3082
R175 source.n28 source.t44 52.3082
R176 source.n46 source.t29 52.3082
R177 source.n103 source.n102 31.4096
R178 source.n85 source.n84 31.4096
R179 source.n77 source.n76 31.4096
R180 source.n59 source.n58 31.4096
R181 source.n7 source.n6 31.4096
R182 source.n25 source.n24 31.4096
R183 source.n33 source.n32 31.4096
R184 source.n51 source.n50 31.4096
R185 source.n59 source.n51 14.4275
R186 source.n94 source.t43 9.9005
R187 source.n94 source.t40 9.9005
R188 source.n92 source.t45 9.9005
R189 source.n92 source.t32 9.9005
R190 source.n90 source.t33 9.9005
R191 source.n90 source.t30 9.9005
R192 source.n88 source.t25 9.9005
R193 source.n88 source.t37 9.9005
R194 source.n86 source.t34 9.9005
R195 source.n86 source.t41 9.9005
R196 source.n68 source.t4 9.9005
R197 source.n68 source.t10 9.9005
R198 source.n66 source.t5 9.9005
R199 source.n66 source.t21 9.9005
R200 source.n64 source.t2 9.9005
R201 source.n64 source.t19 9.9005
R202 source.n62 source.t7 9.9005
R203 source.n62 source.t46 9.9005
R204 source.n60 source.t6 9.9005
R205 source.n60 source.t17 9.9005
R206 source.n8 source.t8 9.9005
R207 source.n8 source.t15 9.9005
R208 source.n10 source.t3 9.9005
R209 source.n10 source.t14 9.9005
R210 source.n12 source.t13 9.9005
R211 source.n12 source.t16 9.9005
R212 source.n14 source.t1 9.9005
R213 source.n14 source.t0 9.9005
R214 source.n16 source.t47 9.9005
R215 source.n16 source.t18 9.9005
R216 source.n34 source.t36 9.9005
R217 source.n34 source.t23 9.9005
R218 source.n36 source.t27 9.9005
R219 source.n36 source.t22 9.9005
R220 source.n38 source.t31 9.9005
R221 source.n38 source.t24 9.9005
R222 source.n40 source.t35 9.9005
R223 source.n40 source.t38 9.9005
R224 source.n42 source.t42 9.9005
R225 source.n42 source.t39 9.9005
R226 source.n99 source.n97 9.71174
R227 source.n81 source.n79 9.71174
R228 source.n73 source.n71 9.71174
R229 source.n55 source.n53 9.71174
R230 source.n3 source.n1 9.71174
R231 source.n21 source.n19 9.71174
R232 source.n29 source.n27 9.71174
R233 source.n47 source.n45 9.71174
R234 source.n102 source.n101 9.45567
R235 source.n84 source.n83 9.45567
R236 source.n76 source.n75 9.45567
R237 source.n58 source.n57 9.45567
R238 source.n6 source.n5 9.45567
R239 source.n24 source.n23 9.45567
R240 source.n32 source.n31 9.45567
R241 source.n50 source.n49 9.45567
R242 source.n101 source.n100 9.3005
R243 source.n83 source.n82 9.3005
R244 source.n75 source.n74 9.3005
R245 source.n57 source.n56 9.3005
R246 source.n5 source.n4 9.3005
R247 source.n23 source.n22 9.3005
R248 source.n31 source.n30 9.3005
R249 source.n49 source.n48 9.3005
R250 source.n104 source.n7 8.8068
R251 source.n102 source.n96 8.14595
R252 source.n84 source.n78 8.14595
R253 source.n76 source.n70 8.14595
R254 source.n58 source.n52 8.14595
R255 source.n6 source.n0 8.14595
R256 source.n24 source.n18 8.14595
R257 source.n32 source.n26 8.14595
R258 source.n50 source.n44 8.14595
R259 source.n100 source.n99 7.3702
R260 source.n82 source.n81 7.3702
R261 source.n74 source.n73 7.3702
R262 source.n56 source.n55 7.3702
R263 source.n4 source.n3 7.3702
R264 source.n22 source.n21 7.3702
R265 source.n30 source.n29 7.3702
R266 source.n48 source.n47 7.3702
R267 source.n100 source.n96 5.81868
R268 source.n82 source.n78 5.81868
R269 source.n74 source.n70 5.81868
R270 source.n56 source.n52 5.81868
R271 source.n4 source.n0 5.81868
R272 source.n22 source.n18 5.81868
R273 source.n30 source.n26 5.81868
R274 source.n48 source.n44 5.81868
R275 source.n104 source.n103 5.62119
R276 source.n101 source.n97 3.44771
R277 source.n83 source.n79 3.44771
R278 source.n75 source.n71 3.44771
R279 source.n57 source.n53 3.44771
R280 source.n5 source.n1 3.44771
R281 source.n23 source.n19 3.44771
R282 source.n31 source.n27 3.44771
R283 source.n49 source.n45 3.44771
R284 source.n51 source.n43 0.716017
R285 source.n43 source.n41 0.716017
R286 source.n41 source.n39 0.716017
R287 source.n39 source.n37 0.716017
R288 source.n37 source.n35 0.716017
R289 source.n35 source.n33 0.716017
R290 source.n25 source.n17 0.716017
R291 source.n17 source.n15 0.716017
R292 source.n15 source.n13 0.716017
R293 source.n13 source.n11 0.716017
R294 source.n11 source.n9 0.716017
R295 source.n9 source.n7 0.716017
R296 source.n61 source.n59 0.716017
R297 source.n63 source.n61 0.716017
R298 source.n65 source.n63 0.716017
R299 source.n67 source.n65 0.716017
R300 source.n69 source.n67 0.716017
R301 source.n77 source.n69 0.716017
R302 source.n87 source.n85 0.716017
R303 source.n89 source.n87 0.716017
R304 source.n91 source.n89 0.716017
R305 source.n93 source.n91 0.716017
R306 source.n95 source.n93 0.716017
R307 source.n103 source.n95 0.716017
R308 source.n33 source.n25 0.470328
R309 source.n85 source.n77 0.470328
R310 source source.n104 0.188
R311 drain_right.n13 drain_right.n11 101.511
R312 drain_right.n7 drain_right.n5 101.511
R313 drain_right.n2 drain_right.n0 101.511
R314 drain_right.n13 drain_right.n12 100.796
R315 drain_right.n15 drain_right.n14 100.796
R316 drain_right.n17 drain_right.n16 100.796
R317 drain_right.n19 drain_right.n18 100.796
R318 drain_right.n21 drain_right.n20 100.796
R319 drain_right.n7 drain_right.n6 100.796
R320 drain_right.n9 drain_right.n8 100.796
R321 drain_right.n4 drain_right.n3 100.796
R322 drain_right.n2 drain_right.n1 100.796
R323 drain_right drain_right.n10 26.0355
R324 drain_right.n5 drain_right.t0 9.9005
R325 drain_right.n5 drain_right.t5 9.9005
R326 drain_right.n6 drain_right.t20 9.9005
R327 drain_right.n6 drain_right.t11 9.9005
R328 drain_right.n8 drain_right.t17 9.9005
R329 drain_right.n8 drain_right.t8 9.9005
R330 drain_right.n3 drain_right.t14 9.9005
R331 drain_right.n3 drain_right.t21 9.9005
R332 drain_right.n1 drain_right.t6 9.9005
R333 drain_right.n1 drain_right.t1 9.9005
R334 drain_right.n0 drain_right.t3 9.9005
R335 drain_right.n0 drain_right.t23 9.9005
R336 drain_right.n11 drain_right.t19 9.9005
R337 drain_right.n11 drain_right.t10 9.9005
R338 drain_right.n12 drain_right.t4 9.9005
R339 drain_right.n12 drain_right.t15 9.9005
R340 drain_right.n14 drain_right.t13 9.9005
R341 drain_right.n14 drain_right.t16 9.9005
R342 drain_right.n16 drain_right.t12 9.9005
R343 drain_right.n16 drain_right.t22 9.9005
R344 drain_right.n18 drain_right.t18 9.9005
R345 drain_right.n18 drain_right.t7 9.9005
R346 drain_right.n20 drain_right.t2 9.9005
R347 drain_right.n20 drain_right.t9 9.9005
R348 drain_right drain_right.n21 6.36873
R349 drain_right.n9 drain_right.n7 0.716017
R350 drain_right.n4 drain_right.n2 0.716017
R351 drain_right.n21 drain_right.n19 0.716017
R352 drain_right.n19 drain_right.n17 0.716017
R353 drain_right.n17 drain_right.n15 0.716017
R354 drain_right.n15 drain_right.n13 0.716017
R355 drain_right.n10 drain_right.n9 0.302913
R356 drain_right.n10 drain_right.n4 0.302913
R357 plus.n11 plus.t5 201.325
R358 plus.n45 plus.t21 201.325
R359 plus.n32 plus.t0 174.966
R360 plus.n30 plus.t1 174.966
R361 plus.n29 plus.t14 174.966
R362 plus.n3 plus.t4 174.966
R363 plus.n23 plus.t19 174.966
R364 plus.n22 plus.t12 174.966
R365 plus.n6 plus.t23 174.966
R366 plus.n17 plus.t18 174.966
R367 plus.n15 plus.t9 174.966
R368 plus.n9 plus.t20 174.966
R369 plus.n10 plus.t16 174.966
R370 plus.n66 plus.t11 174.966
R371 plus.n64 plus.t22 174.966
R372 plus.n63 plus.t13 174.966
R373 plus.n37 plus.t8 174.966
R374 plus.n57 plus.t15 174.966
R375 plus.n56 plus.t7 174.966
R376 plus.n40 plus.t2 174.966
R377 plus.n51 plus.t10 174.966
R378 plus.n49 plus.t6 174.966
R379 plus.n43 plus.t17 174.966
R380 plus.n44 plus.t3 174.966
R381 plus.n12 plus.n9 161.3
R382 plus.n14 plus.n13 161.3
R383 plus.n15 plus.n8 161.3
R384 plus.n16 plus.n7 161.3
R385 plus.n18 plus.n17 161.3
R386 plus.n19 plus.n6 161.3
R387 plus.n21 plus.n20 161.3
R388 plus.n22 plus.n5 161.3
R389 plus.n23 plus.n4 161.3
R390 plus.n25 plus.n24 161.3
R391 plus.n26 plus.n3 161.3
R392 plus.n28 plus.n27 161.3
R393 plus.n29 plus.n2 161.3
R394 plus.n30 plus.n1 161.3
R395 plus.n31 plus.n0 161.3
R396 plus.n33 plus.n32 161.3
R397 plus.n46 plus.n43 161.3
R398 plus.n48 plus.n47 161.3
R399 plus.n49 plus.n42 161.3
R400 plus.n50 plus.n41 161.3
R401 plus.n52 plus.n51 161.3
R402 plus.n53 plus.n40 161.3
R403 plus.n55 plus.n54 161.3
R404 plus.n56 plus.n39 161.3
R405 plus.n57 plus.n38 161.3
R406 plus.n59 plus.n58 161.3
R407 plus.n60 plus.n37 161.3
R408 plus.n62 plus.n61 161.3
R409 plus.n63 plus.n36 161.3
R410 plus.n64 plus.n35 161.3
R411 plus.n65 plus.n34 161.3
R412 plus.n67 plus.n66 161.3
R413 plus.n30 plus.n29 48.2005
R414 plus.n23 plus.n22 48.2005
R415 plus.n17 plus.n6 48.2005
R416 plus.n10 plus.n9 48.2005
R417 plus.n64 plus.n63 48.2005
R418 plus.n57 plus.n56 48.2005
R419 plus.n51 plus.n40 48.2005
R420 plus.n44 plus.n43 48.2005
R421 plus.n24 plus.n3 47.4702
R422 plus.n16 plus.n15 47.4702
R423 plus.n58 plus.n37 47.4702
R424 plus.n50 plus.n49 47.4702
R425 plus.n32 plus.n31 46.0096
R426 plus.n66 plus.n65 46.0096
R427 plus.n12 plus.n11 45.0871
R428 plus.n46 plus.n45 45.0871
R429 plus plus.n67 30.1278
R430 plus.n28 plus.n3 25.5611
R431 plus.n15 plus.n14 25.5611
R432 plus.n62 plus.n37 25.5611
R433 plus.n49 plus.n48 25.5611
R434 plus.n21 plus.n6 24.1005
R435 plus.n22 plus.n21 24.1005
R436 plus.n56 plus.n55 24.1005
R437 plus.n55 plus.n40 24.1005
R438 plus.n29 plus.n28 22.6399
R439 plus.n14 plus.n9 22.6399
R440 plus.n63 plus.n62 22.6399
R441 plus.n48 plus.n43 22.6399
R442 plus.n11 plus.n10 14.1472
R443 plus.n45 plus.n44 14.1472
R444 plus plus.n33 8.38308
R445 plus.n31 plus.n30 2.19141
R446 plus.n65 plus.n64 2.19141
R447 plus.n24 plus.n23 0.730803
R448 plus.n17 plus.n16 0.730803
R449 plus.n58 plus.n57 0.730803
R450 plus.n51 plus.n50 0.730803
R451 plus.n13 plus.n12 0.189894
R452 plus.n13 plus.n8 0.189894
R453 plus.n8 plus.n7 0.189894
R454 plus.n18 plus.n7 0.189894
R455 plus.n19 plus.n18 0.189894
R456 plus.n20 plus.n19 0.189894
R457 plus.n20 plus.n5 0.189894
R458 plus.n5 plus.n4 0.189894
R459 plus.n25 plus.n4 0.189894
R460 plus.n26 plus.n25 0.189894
R461 plus.n27 plus.n26 0.189894
R462 plus.n27 plus.n2 0.189894
R463 plus.n2 plus.n1 0.189894
R464 plus.n1 plus.n0 0.189894
R465 plus.n33 plus.n0 0.189894
R466 plus.n67 plus.n34 0.189894
R467 plus.n35 plus.n34 0.189894
R468 plus.n36 plus.n35 0.189894
R469 plus.n61 plus.n36 0.189894
R470 plus.n61 plus.n60 0.189894
R471 plus.n60 plus.n59 0.189894
R472 plus.n59 plus.n38 0.189894
R473 plus.n39 plus.n38 0.189894
R474 plus.n54 plus.n39 0.189894
R475 plus.n54 plus.n53 0.189894
R476 plus.n53 plus.n52 0.189894
R477 plus.n52 plus.n41 0.189894
R478 plus.n42 plus.n41 0.189894
R479 plus.n47 plus.n42 0.189894
R480 plus.n47 plus.n46 0.189894
R481 drain_left.n13 drain_left.n11 101.511
R482 drain_left.n7 drain_left.n5 101.511
R483 drain_left.n2 drain_left.n0 101.511
R484 drain_left.n21 drain_left.n20 100.796
R485 drain_left.n19 drain_left.n18 100.796
R486 drain_left.n17 drain_left.n16 100.796
R487 drain_left.n15 drain_left.n14 100.796
R488 drain_left.n13 drain_left.n12 100.796
R489 drain_left.n7 drain_left.n6 100.796
R490 drain_left.n9 drain_left.n8 100.796
R491 drain_left.n4 drain_left.n3 100.796
R492 drain_left.n2 drain_left.n1 100.796
R493 drain_left drain_left.n10 26.5887
R494 drain_left.n5 drain_left.t20 9.9005
R495 drain_left.n5 drain_left.t2 9.9005
R496 drain_left.n6 drain_left.t17 9.9005
R497 drain_left.n6 drain_left.t6 9.9005
R498 drain_left.n8 drain_left.t21 9.9005
R499 drain_left.n8 drain_left.t13 9.9005
R500 drain_left.n3 drain_left.t8 9.9005
R501 drain_left.n3 drain_left.t16 9.9005
R502 drain_left.n1 drain_left.t10 9.9005
R503 drain_left.n1 drain_left.t15 9.9005
R504 drain_left.n0 drain_left.t12 9.9005
R505 drain_left.n0 drain_left.t1 9.9005
R506 drain_left.n20 drain_left.t22 9.9005
R507 drain_left.n20 drain_left.t23 9.9005
R508 drain_left.n18 drain_left.t19 9.9005
R509 drain_left.n18 drain_left.t9 9.9005
R510 drain_left.n16 drain_left.t11 9.9005
R511 drain_left.n16 drain_left.t4 9.9005
R512 drain_left.n14 drain_left.t5 9.9005
R513 drain_left.n14 drain_left.t0 9.9005
R514 drain_left.n12 drain_left.t3 9.9005
R515 drain_left.n12 drain_left.t14 9.9005
R516 drain_left.n11 drain_left.t18 9.9005
R517 drain_left.n11 drain_left.t7 9.9005
R518 drain_left drain_left.n21 6.36873
R519 drain_left.n9 drain_left.n7 0.716017
R520 drain_left.n4 drain_left.n2 0.716017
R521 drain_left.n15 drain_left.n13 0.716017
R522 drain_left.n17 drain_left.n15 0.716017
R523 drain_left.n19 drain_left.n17 0.716017
R524 drain_left.n21 drain_left.n19 0.716017
R525 drain_left.n10 drain_left.n9 0.302913
R526 drain_left.n10 drain_left.n4 0.302913
C0 drain_right source 9.20647f
C1 plus minus 4.89787f
C2 plus drain_right 0.450398f
C3 plus source 3.26779f
C4 minus drain_left 0.179685f
C5 drain_left drain_right 1.55979f
C6 drain_left source 9.204929f
C7 minus drain_right 2.63813f
C8 plus drain_left 2.92432f
C9 minus source 3.25382f
C10 drain_right a_n2874_n1288# 5.45882f
C11 drain_left a_n2874_n1288# 5.88864f
C12 source a_n2874_n1288# 3.523933f
C13 minus a_n2874_n1288# 10.695829f
C14 plus a_n2874_n1288# 12.121819f
C15 drain_left.t12 a_n2874_n1288# 0.045758f
C16 drain_left.t1 a_n2874_n1288# 0.045758f
C17 drain_left.n0 a_n2874_n1288# 0.290049f
C18 drain_left.t10 a_n2874_n1288# 0.045758f
C19 drain_left.t15 a_n2874_n1288# 0.045758f
C20 drain_left.n1 a_n2874_n1288# 0.287464f
C21 drain_left.n2 a_n2874_n1288# 0.719274f
C22 drain_left.t8 a_n2874_n1288# 0.045758f
C23 drain_left.t16 a_n2874_n1288# 0.045758f
C24 drain_left.n3 a_n2874_n1288# 0.287464f
C25 drain_left.n4 a_n2874_n1288# 0.31878f
C26 drain_left.t20 a_n2874_n1288# 0.045758f
C27 drain_left.t2 a_n2874_n1288# 0.045758f
C28 drain_left.n5 a_n2874_n1288# 0.290049f
C29 drain_left.t17 a_n2874_n1288# 0.045758f
C30 drain_left.t6 a_n2874_n1288# 0.045758f
C31 drain_left.n6 a_n2874_n1288# 0.287464f
C32 drain_left.n7 a_n2874_n1288# 0.719274f
C33 drain_left.t21 a_n2874_n1288# 0.045758f
C34 drain_left.t13 a_n2874_n1288# 0.045758f
C35 drain_left.n8 a_n2874_n1288# 0.287464f
C36 drain_left.n9 a_n2874_n1288# 0.31878f
C37 drain_left.n10 a_n2874_n1288# 1.1348f
C38 drain_left.t18 a_n2874_n1288# 0.045758f
C39 drain_left.t7 a_n2874_n1288# 0.045758f
C40 drain_left.n11 a_n2874_n1288# 0.290051f
C41 drain_left.t3 a_n2874_n1288# 0.045758f
C42 drain_left.t14 a_n2874_n1288# 0.045758f
C43 drain_left.n12 a_n2874_n1288# 0.287465f
C44 drain_left.n13 a_n2874_n1288# 0.719271f
C45 drain_left.t5 a_n2874_n1288# 0.045758f
C46 drain_left.t0 a_n2874_n1288# 0.045758f
C47 drain_left.n14 a_n2874_n1288# 0.287465f
C48 drain_left.n15 a_n2874_n1288# 0.355098f
C49 drain_left.t11 a_n2874_n1288# 0.045758f
C50 drain_left.t4 a_n2874_n1288# 0.045758f
C51 drain_left.n16 a_n2874_n1288# 0.287465f
C52 drain_left.n17 a_n2874_n1288# 0.355098f
C53 drain_left.t19 a_n2874_n1288# 0.045758f
C54 drain_left.t9 a_n2874_n1288# 0.045758f
C55 drain_left.n18 a_n2874_n1288# 0.287465f
C56 drain_left.n19 a_n2874_n1288# 0.355098f
C57 drain_left.t22 a_n2874_n1288# 0.045758f
C58 drain_left.t23 a_n2874_n1288# 0.045758f
C59 drain_left.n20 a_n2874_n1288# 0.287465f
C60 drain_left.n21 a_n2874_n1288# 0.603837f
C61 plus.n0 a_n2874_n1288# 0.046291f
C62 plus.t0 a_n2874_n1288# 0.14335f
C63 plus.t1 a_n2874_n1288# 0.14335f
C64 plus.n1 a_n2874_n1288# 0.046291f
C65 plus.t14 a_n2874_n1288# 0.14335f
C66 plus.n2 a_n2874_n1288# 0.046291f
C67 plus.t4 a_n2874_n1288# 0.14335f
C68 plus.n3 a_n2874_n1288# 0.108112f
C69 plus.n4 a_n2874_n1288# 0.046291f
C70 plus.t19 a_n2874_n1288# 0.14335f
C71 plus.t12 a_n2874_n1288# 0.14335f
C72 plus.n5 a_n2874_n1288# 0.046291f
C73 plus.t23 a_n2874_n1288# 0.14335f
C74 plus.n6 a_n2874_n1288# 0.10797f
C75 plus.n7 a_n2874_n1288# 0.046291f
C76 plus.t18 a_n2874_n1288# 0.14335f
C77 plus.t9 a_n2874_n1288# 0.14335f
C78 plus.n8 a_n2874_n1288# 0.046291f
C79 plus.t20 a_n2874_n1288# 0.14335f
C80 plus.n9 a_n2874_n1288# 0.107684f
C81 plus.t16 a_n2874_n1288# 0.14335f
C82 plus.n10 a_n2874_n1288# 0.113162f
C83 plus.t5 a_n2874_n1288# 0.156861f
C84 plus.n11 a_n2874_n1288# 0.091267f
C85 plus.n12 a_n2874_n1288# 0.18796f
C86 plus.n13 a_n2874_n1288# 0.046291f
C87 plus.n14 a_n2874_n1288# 0.010504f
C88 plus.n15 a_n2874_n1288# 0.108112f
C89 plus.n16 a_n2874_n1288# 0.010504f
C90 plus.n17 a_n2874_n1288# 0.103403f
C91 plus.n18 a_n2874_n1288# 0.046291f
C92 plus.n19 a_n2874_n1288# 0.046291f
C93 plus.n20 a_n2874_n1288# 0.046291f
C94 plus.n21 a_n2874_n1288# 0.010504f
C95 plus.n22 a_n2874_n1288# 0.10797f
C96 plus.n23 a_n2874_n1288# 0.103403f
C97 plus.n24 a_n2874_n1288# 0.010504f
C98 plus.n25 a_n2874_n1288# 0.046291f
C99 plus.n26 a_n2874_n1288# 0.046291f
C100 plus.n27 a_n2874_n1288# 0.046291f
C101 plus.n28 a_n2874_n1288# 0.010504f
C102 plus.n29 a_n2874_n1288# 0.107684f
C103 plus.n30 a_n2874_n1288# 0.103689f
C104 plus.n31 a_n2874_n1288# 0.010504f
C105 plus.n32 a_n2874_n1288# 0.102832f
C106 plus.n33 a_n2874_n1288# 0.334031f
C107 plus.n34 a_n2874_n1288# 0.046291f
C108 plus.t11 a_n2874_n1288# 0.14335f
C109 plus.n35 a_n2874_n1288# 0.046291f
C110 plus.t22 a_n2874_n1288# 0.14335f
C111 plus.n36 a_n2874_n1288# 0.046291f
C112 plus.t13 a_n2874_n1288# 0.14335f
C113 plus.t8 a_n2874_n1288# 0.14335f
C114 plus.n37 a_n2874_n1288# 0.108112f
C115 plus.n38 a_n2874_n1288# 0.046291f
C116 plus.t15 a_n2874_n1288# 0.14335f
C117 plus.n39 a_n2874_n1288# 0.046291f
C118 plus.t7 a_n2874_n1288# 0.14335f
C119 plus.t2 a_n2874_n1288# 0.14335f
C120 plus.n40 a_n2874_n1288# 0.10797f
C121 plus.n41 a_n2874_n1288# 0.046291f
C122 plus.t10 a_n2874_n1288# 0.14335f
C123 plus.n42 a_n2874_n1288# 0.046291f
C124 plus.t6 a_n2874_n1288# 0.14335f
C125 plus.t17 a_n2874_n1288# 0.14335f
C126 plus.n43 a_n2874_n1288# 0.107684f
C127 plus.t21 a_n2874_n1288# 0.156861f
C128 plus.t3 a_n2874_n1288# 0.14335f
C129 plus.n44 a_n2874_n1288# 0.113162f
C130 plus.n45 a_n2874_n1288# 0.091267f
C131 plus.n46 a_n2874_n1288# 0.18796f
C132 plus.n47 a_n2874_n1288# 0.046291f
C133 plus.n48 a_n2874_n1288# 0.010504f
C134 plus.n49 a_n2874_n1288# 0.108112f
C135 plus.n50 a_n2874_n1288# 0.010504f
C136 plus.n51 a_n2874_n1288# 0.103403f
C137 plus.n52 a_n2874_n1288# 0.046291f
C138 plus.n53 a_n2874_n1288# 0.046291f
C139 plus.n54 a_n2874_n1288# 0.046291f
C140 plus.n55 a_n2874_n1288# 0.010504f
C141 plus.n56 a_n2874_n1288# 0.10797f
C142 plus.n57 a_n2874_n1288# 0.103403f
C143 plus.n58 a_n2874_n1288# 0.010504f
C144 plus.n59 a_n2874_n1288# 0.046291f
C145 plus.n60 a_n2874_n1288# 0.046291f
C146 plus.n61 a_n2874_n1288# 0.046291f
C147 plus.n62 a_n2874_n1288# 0.010504f
C148 plus.n63 a_n2874_n1288# 0.107684f
C149 plus.n64 a_n2874_n1288# 0.103689f
C150 plus.n65 a_n2874_n1288# 0.010504f
C151 plus.n66 a_n2874_n1288# 0.102832f
C152 plus.n67 a_n2874_n1288# 1.30682f
C153 drain_right.t3 a_n2874_n1288# 0.045045f
C154 drain_right.t23 a_n2874_n1288# 0.045045f
C155 drain_right.n0 a_n2874_n1288# 0.285531f
C156 drain_right.t6 a_n2874_n1288# 0.045045f
C157 drain_right.t1 a_n2874_n1288# 0.045045f
C158 drain_right.n1 a_n2874_n1288# 0.282986f
C159 drain_right.n2 a_n2874_n1288# 0.708068f
C160 drain_right.t14 a_n2874_n1288# 0.045045f
C161 drain_right.t21 a_n2874_n1288# 0.045045f
C162 drain_right.n3 a_n2874_n1288# 0.282986f
C163 drain_right.n4 a_n2874_n1288# 0.313813f
C164 drain_right.t0 a_n2874_n1288# 0.045045f
C165 drain_right.t5 a_n2874_n1288# 0.045045f
C166 drain_right.n5 a_n2874_n1288# 0.285531f
C167 drain_right.t20 a_n2874_n1288# 0.045045f
C168 drain_right.t11 a_n2874_n1288# 0.045045f
C169 drain_right.n6 a_n2874_n1288# 0.282986f
C170 drain_right.n7 a_n2874_n1288# 0.708068f
C171 drain_right.t17 a_n2874_n1288# 0.045045f
C172 drain_right.t8 a_n2874_n1288# 0.045045f
C173 drain_right.n8 a_n2874_n1288# 0.282986f
C174 drain_right.n9 a_n2874_n1288# 0.313813f
C175 drain_right.n10 a_n2874_n1288# 1.06184f
C176 drain_right.t19 a_n2874_n1288# 0.045045f
C177 drain_right.t10 a_n2874_n1288# 0.045045f
C178 drain_right.n11 a_n2874_n1288# 0.285532f
C179 drain_right.t4 a_n2874_n1288# 0.045045f
C180 drain_right.t15 a_n2874_n1288# 0.045045f
C181 drain_right.n12 a_n2874_n1288# 0.282987f
C182 drain_right.n13 a_n2874_n1288# 0.708066f
C183 drain_right.t13 a_n2874_n1288# 0.045045f
C184 drain_right.t16 a_n2874_n1288# 0.045045f
C185 drain_right.n14 a_n2874_n1288# 0.282987f
C186 drain_right.n15 a_n2874_n1288# 0.349565f
C187 drain_right.t12 a_n2874_n1288# 0.045045f
C188 drain_right.t22 a_n2874_n1288# 0.045045f
C189 drain_right.n16 a_n2874_n1288# 0.282987f
C190 drain_right.n17 a_n2874_n1288# 0.349565f
C191 drain_right.t18 a_n2874_n1288# 0.045045f
C192 drain_right.t7 a_n2874_n1288# 0.045045f
C193 drain_right.n18 a_n2874_n1288# 0.282987f
C194 drain_right.n19 a_n2874_n1288# 0.349565f
C195 drain_right.t2 a_n2874_n1288# 0.045045f
C196 drain_right.t9 a_n2874_n1288# 0.045045f
C197 drain_right.n20 a_n2874_n1288# 0.282987f
C198 drain_right.n21 a_n2874_n1288# 0.594429f
C199 source.n0 a_n2874_n1288# 0.047968f
C200 source.n1 a_n2874_n1288# 0.106135f
C201 source.t11 a_n2874_n1288# 0.079649f
C202 source.n2 a_n2874_n1288# 0.083066f
C203 source.n3 a_n2874_n1288# 0.026777f
C204 source.n4 a_n2874_n1288# 0.01766f
C205 source.n5 a_n2874_n1288# 0.233948f
C206 source.n6 a_n2874_n1288# 0.052584f
C207 source.n7 a_n2874_n1288# 0.528601f
C208 source.t8 a_n2874_n1288# 0.051941f
C209 source.t15 a_n2874_n1288# 0.051941f
C210 source.n8 a_n2874_n1288# 0.277677f
C211 source.n9 a_n2874_n1288# 0.407051f
C212 source.t3 a_n2874_n1288# 0.051941f
C213 source.t14 a_n2874_n1288# 0.051941f
C214 source.n10 a_n2874_n1288# 0.277677f
C215 source.n11 a_n2874_n1288# 0.407051f
C216 source.t13 a_n2874_n1288# 0.051941f
C217 source.t16 a_n2874_n1288# 0.051941f
C218 source.n12 a_n2874_n1288# 0.277677f
C219 source.n13 a_n2874_n1288# 0.407051f
C220 source.t1 a_n2874_n1288# 0.051941f
C221 source.t0 a_n2874_n1288# 0.051941f
C222 source.n14 a_n2874_n1288# 0.277677f
C223 source.n15 a_n2874_n1288# 0.407051f
C224 source.t47 a_n2874_n1288# 0.051941f
C225 source.t18 a_n2874_n1288# 0.051941f
C226 source.n16 a_n2874_n1288# 0.277677f
C227 source.n17 a_n2874_n1288# 0.407051f
C228 source.n18 a_n2874_n1288# 0.047968f
C229 source.n19 a_n2874_n1288# 0.106135f
C230 source.t20 a_n2874_n1288# 0.079649f
C231 source.n20 a_n2874_n1288# 0.083066f
C232 source.n21 a_n2874_n1288# 0.026777f
C233 source.n22 a_n2874_n1288# 0.01766f
C234 source.n23 a_n2874_n1288# 0.233948f
C235 source.n24 a_n2874_n1288# 0.052584f
C236 source.n25 a_n2874_n1288# 0.15258f
C237 source.n26 a_n2874_n1288# 0.047968f
C238 source.n27 a_n2874_n1288# 0.106135f
C239 source.t44 a_n2874_n1288# 0.079649f
C240 source.n28 a_n2874_n1288# 0.083066f
C241 source.n29 a_n2874_n1288# 0.026777f
C242 source.n30 a_n2874_n1288# 0.01766f
C243 source.n31 a_n2874_n1288# 0.233948f
C244 source.n32 a_n2874_n1288# 0.052584f
C245 source.n33 a_n2874_n1288# 0.15258f
C246 source.t36 a_n2874_n1288# 0.051941f
C247 source.t23 a_n2874_n1288# 0.051941f
C248 source.n34 a_n2874_n1288# 0.277677f
C249 source.n35 a_n2874_n1288# 0.407051f
C250 source.t27 a_n2874_n1288# 0.051941f
C251 source.t22 a_n2874_n1288# 0.051941f
C252 source.n36 a_n2874_n1288# 0.277677f
C253 source.n37 a_n2874_n1288# 0.407051f
C254 source.t31 a_n2874_n1288# 0.051941f
C255 source.t24 a_n2874_n1288# 0.051941f
C256 source.n38 a_n2874_n1288# 0.277677f
C257 source.n39 a_n2874_n1288# 0.407051f
C258 source.t35 a_n2874_n1288# 0.051941f
C259 source.t38 a_n2874_n1288# 0.051941f
C260 source.n40 a_n2874_n1288# 0.277677f
C261 source.n41 a_n2874_n1288# 0.407051f
C262 source.t42 a_n2874_n1288# 0.051941f
C263 source.t39 a_n2874_n1288# 0.051941f
C264 source.n42 a_n2874_n1288# 0.277677f
C265 source.n43 a_n2874_n1288# 0.407051f
C266 source.n44 a_n2874_n1288# 0.047968f
C267 source.n45 a_n2874_n1288# 0.106135f
C268 source.t29 a_n2874_n1288# 0.079649f
C269 source.n46 a_n2874_n1288# 0.083066f
C270 source.n47 a_n2874_n1288# 0.026777f
C271 source.n48 a_n2874_n1288# 0.01766f
C272 source.n49 a_n2874_n1288# 0.233948f
C273 source.n50 a_n2874_n1288# 0.052584f
C274 source.n51 a_n2874_n1288# 0.839118f
C275 source.n52 a_n2874_n1288# 0.047968f
C276 source.n53 a_n2874_n1288# 0.106135f
C277 source.t12 a_n2874_n1288# 0.079649f
C278 source.n54 a_n2874_n1288# 0.083066f
C279 source.n55 a_n2874_n1288# 0.026777f
C280 source.n56 a_n2874_n1288# 0.01766f
C281 source.n57 a_n2874_n1288# 0.233948f
C282 source.n58 a_n2874_n1288# 0.052584f
C283 source.n59 a_n2874_n1288# 0.839118f
C284 source.t6 a_n2874_n1288# 0.051941f
C285 source.t17 a_n2874_n1288# 0.051941f
C286 source.n60 a_n2874_n1288# 0.277675f
C287 source.n61 a_n2874_n1288# 0.407052f
C288 source.t7 a_n2874_n1288# 0.051941f
C289 source.t46 a_n2874_n1288# 0.051941f
C290 source.n62 a_n2874_n1288# 0.277675f
C291 source.n63 a_n2874_n1288# 0.407052f
C292 source.t2 a_n2874_n1288# 0.051941f
C293 source.t19 a_n2874_n1288# 0.051941f
C294 source.n64 a_n2874_n1288# 0.277675f
C295 source.n65 a_n2874_n1288# 0.407052f
C296 source.t5 a_n2874_n1288# 0.051941f
C297 source.t21 a_n2874_n1288# 0.051941f
C298 source.n66 a_n2874_n1288# 0.277675f
C299 source.n67 a_n2874_n1288# 0.407052f
C300 source.t4 a_n2874_n1288# 0.051941f
C301 source.t10 a_n2874_n1288# 0.051941f
C302 source.n68 a_n2874_n1288# 0.277675f
C303 source.n69 a_n2874_n1288# 0.407052f
C304 source.n70 a_n2874_n1288# 0.047968f
C305 source.n71 a_n2874_n1288# 0.106135f
C306 source.t9 a_n2874_n1288# 0.079649f
C307 source.n72 a_n2874_n1288# 0.083066f
C308 source.n73 a_n2874_n1288# 0.026777f
C309 source.n74 a_n2874_n1288# 0.01766f
C310 source.n75 a_n2874_n1288# 0.233948f
C311 source.n76 a_n2874_n1288# 0.052584f
C312 source.n77 a_n2874_n1288# 0.15258f
C313 source.n78 a_n2874_n1288# 0.047968f
C314 source.n79 a_n2874_n1288# 0.106135f
C315 source.t26 a_n2874_n1288# 0.079649f
C316 source.n80 a_n2874_n1288# 0.083066f
C317 source.n81 a_n2874_n1288# 0.026777f
C318 source.n82 a_n2874_n1288# 0.01766f
C319 source.n83 a_n2874_n1288# 0.233948f
C320 source.n84 a_n2874_n1288# 0.052584f
C321 source.n85 a_n2874_n1288# 0.15258f
C322 source.t34 a_n2874_n1288# 0.051941f
C323 source.t41 a_n2874_n1288# 0.051941f
C324 source.n86 a_n2874_n1288# 0.277675f
C325 source.n87 a_n2874_n1288# 0.407052f
C326 source.t25 a_n2874_n1288# 0.051941f
C327 source.t37 a_n2874_n1288# 0.051941f
C328 source.n88 a_n2874_n1288# 0.277675f
C329 source.n89 a_n2874_n1288# 0.407052f
C330 source.t33 a_n2874_n1288# 0.051941f
C331 source.t30 a_n2874_n1288# 0.051941f
C332 source.n90 a_n2874_n1288# 0.277675f
C333 source.n91 a_n2874_n1288# 0.407052f
C334 source.t45 a_n2874_n1288# 0.051941f
C335 source.t32 a_n2874_n1288# 0.051941f
C336 source.n92 a_n2874_n1288# 0.277675f
C337 source.n93 a_n2874_n1288# 0.407052f
C338 source.t43 a_n2874_n1288# 0.051941f
C339 source.t40 a_n2874_n1288# 0.051941f
C340 source.n94 a_n2874_n1288# 0.277675f
C341 source.n95 a_n2874_n1288# 0.407052f
C342 source.n96 a_n2874_n1288# 0.047968f
C343 source.n97 a_n2874_n1288# 0.106135f
C344 source.t28 a_n2874_n1288# 0.079649f
C345 source.n98 a_n2874_n1288# 0.083066f
C346 source.n99 a_n2874_n1288# 0.026777f
C347 source.n100 a_n2874_n1288# 0.01766f
C348 source.n101 a_n2874_n1288# 0.233948f
C349 source.n102 a_n2874_n1288# 0.052584f
C350 source.n103 a_n2874_n1288# 0.352611f
C351 source.n104 a_n2874_n1288# 0.820401f
C352 minus.n0 a_n2874_n1288# 0.044663f
C353 minus.t5 a_n2874_n1288# 0.13831f
C354 minus.n1 a_n2874_n1288# 0.103898f
C355 minus.t14 a_n2874_n1288# 0.13831f
C356 minus.n2 a_n2874_n1288# 0.044663f
C357 minus.t11 a_n2874_n1288# 0.13831f
C358 minus.n3 a_n2874_n1288# 0.099767f
C359 minus.n4 a_n2874_n1288# 0.044663f
C360 minus.t7 a_n2874_n1288# 0.13831f
C361 minus.n5 a_n2874_n1288# 0.099767f
C362 minus.t10 a_n2874_n1288# 0.13831f
C363 minus.n6 a_n2874_n1288# 0.044663f
C364 minus.t8 a_n2874_n1288# 0.13831f
C365 minus.n7 a_n2874_n1288# 0.103898f
C366 minus.t13 a_n2874_n1288# 0.151345f
C367 minus.t4 a_n2874_n1288# 0.13831f
C368 minus.n8 a_n2874_n1288# 0.109182f
C369 minus.n9 a_n2874_n1288# 0.088057f
C370 minus.n10 a_n2874_n1288# 0.181351f
C371 minus.n11 a_n2874_n1288# 0.044663f
C372 minus.n12 a_n2874_n1288# 0.010135f
C373 minus.t19 a_n2874_n1288# 0.13831f
C374 minus.n13 a_n2874_n1288# 0.104311f
C375 minus.n14 a_n2874_n1288# 0.010135f
C376 minus.n15 a_n2874_n1288# 0.044663f
C377 minus.n16 a_n2874_n1288# 0.044663f
C378 minus.n17 a_n2874_n1288# 0.044663f
C379 minus.n18 a_n2874_n1288# 0.104173f
C380 minus.n19 a_n2874_n1288# 0.010135f
C381 minus.t1 a_n2874_n1288# 0.13831f
C382 minus.n20 a_n2874_n1288# 0.104173f
C383 minus.n21 a_n2874_n1288# 0.044663f
C384 minus.n22 a_n2874_n1288# 0.044663f
C385 minus.n23 a_n2874_n1288# 0.044663f
C386 minus.n24 a_n2874_n1288# 0.010135f
C387 minus.t16 a_n2874_n1288# 0.13831f
C388 minus.n25 a_n2874_n1288# 0.104311f
C389 minus.n26 a_n2874_n1288# 0.010135f
C390 minus.n27 a_n2874_n1288# 0.044663f
C391 minus.n28 a_n2874_n1288# 0.044663f
C392 minus.n29 a_n2874_n1288# 0.044663f
C393 minus.n30 a_n2874_n1288# 0.100043f
C394 minus.n31 a_n2874_n1288# 0.010135f
C395 minus.t21 a_n2874_n1288# 0.13831f
C396 minus.n32 a_n2874_n1288# 0.099216f
C397 minus.n33 a_n2874_n1288# 1.32675f
C398 minus.n34 a_n2874_n1288# 0.044663f
C399 minus.t12 a_n2874_n1288# 0.13831f
C400 minus.n35 a_n2874_n1288# 0.103898f
C401 minus.n36 a_n2874_n1288# 0.044663f
C402 minus.t15 a_n2874_n1288# 0.13831f
C403 minus.n37 a_n2874_n1288# 0.099767f
C404 minus.n38 a_n2874_n1288# 0.044663f
C405 minus.t9 a_n2874_n1288# 0.13831f
C406 minus.n39 a_n2874_n1288# 0.099767f
C407 minus.n40 a_n2874_n1288# 0.044663f
C408 minus.t17 a_n2874_n1288# 0.13831f
C409 minus.n41 a_n2874_n1288# 0.103898f
C410 minus.t20 a_n2874_n1288# 0.151345f
C411 minus.t0 a_n2874_n1288# 0.13831f
C412 minus.n42 a_n2874_n1288# 0.109182f
C413 minus.n43 a_n2874_n1288# 0.088057f
C414 minus.n44 a_n2874_n1288# 0.181351f
C415 minus.n45 a_n2874_n1288# 0.044663f
C416 minus.n46 a_n2874_n1288# 0.010135f
C417 minus.t22 a_n2874_n1288# 0.13831f
C418 minus.n47 a_n2874_n1288# 0.104311f
C419 minus.n48 a_n2874_n1288# 0.010135f
C420 minus.n49 a_n2874_n1288# 0.044663f
C421 minus.n50 a_n2874_n1288# 0.044663f
C422 minus.n51 a_n2874_n1288# 0.044663f
C423 minus.t2 a_n2874_n1288# 0.13831f
C424 minus.n52 a_n2874_n1288# 0.104173f
C425 minus.n53 a_n2874_n1288# 0.010135f
C426 minus.t6 a_n2874_n1288# 0.13831f
C427 minus.n54 a_n2874_n1288# 0.104173f
C428 minus.n55 a_n2874_n1288# 0.044663f
C429 minus.n56 a_n2874_n1288# 0.044663f
C430 minus.n57 a_n2874_n1288# 0.044663f
C431 minus.n58 a_n2874_n1288# 0.010135f
C432 minus.t3 a_n2874_n1288# 0.13831f
C433 minus.n59 a_n2874_n1288# 0.104311f
C434 minus.n60 a_n2874_n1288# 0.010135f
C435 minus.n61 a_n2874_n1288# 0.044663f
C436 minus.n62 a_n2874_n1288# 0.044663f
C437 minus.n63 a_n2874_n1288# 0.044663f
C438 minus.t23 a_n2874_n1288# 0.13831f
C439 minus.n64 a_n2874_n1288# 0.100043f
C440 minus.n65 a_n2874_n1288# 0.010135f
C441 minus.t18 a_n2874_n1288# 0.13831f
C442 minus.n66 a_n2874_n1288# 0.099216f
C443 minus.n67 a_n2874_n1288# 0.294835f
C444 minus.n68 a_n2874_n1288# 1.62711f
.ends

