* NGSPICE file created from diffpair65.ext - technology: sky130A

.subckt diffpair65 minus drain_right drain_left source plus
X0 source.t23 plus.t0 drain_left.t2 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X1 source.t9 minus.t0 drain_right.t11 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X2 a_n2158_n1088# a_n2158_n1088# a_n2158_n1088# a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.7
X3 source.t22 plus.t1 drain_left.t9 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X4 source.t21 plus.t2 drain_left.t3 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X5 source.t20 plus.t3 drain_left.t4 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X6 drain_right.t10 minus.t1 source.t11 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X7 source.t2 minus.t2 drain_right.t9 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X8 drain_right.t8 minus.t3 source.t4 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X9 drain_right.t7 minus.t4 source.t1 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X10 source.t3 minus.t5 drain_right.t6 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X11 source.t7 minus.t6 drain_right.t5 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X12 source.t19 plus.t4 drain_left.t11 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X13 drain_right.t4 minus.t7 source.t8 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X14 drain_left.t10 plus.t5 source.t18 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X15 drain_left.t8 plus.t6 source.t17 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X16 a_n2158_n1088# a_n2158_n1088# a_n2158_n1088# a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X17 drain_left.t5 plus.t7 source.t16 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X18 a_n2158_n1088# a_n2158_n1088# a_n2158_n1088# a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X19 drain_right.t3 minus.t8 source.t10 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X20 drain_left.t1 plus.t8 source.t15 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X21 drain_right.t2 minus.t9 source.t0 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.7
X22 drain_left.t0 plus.t9 source.t14 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X23 source.t5 minus.t10 drain_right.t1 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X24 source.t6 minus.t11 drain_right.t0 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.7
X25 a_n2158_n1088# a_n2158_n1088# a_n2158_n1088# a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.7
X26 source.t13 plus.t10 drain_left.t7 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
X27 drain_left.t6 plus.t11 source.t12 a_n2158_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.7
R0 plus.n7 plus.n6 161.3
R1 plus.n8 plus.n3 161.3
R2 plus.n10 plus.n9 161.3
R3 plus.n11 plus.n2 161.3
R4 plus.n13 plus.n12 161.3
R5 plus.n14 plus.n1 161.3
R6 plus.n15 plus.n0 161.3
R7 plus.n17 plus.n16 161.3
R8 plus.n25 plus.n24 161.3
R9 plus.n26 plus.n21 161.3
R10 plus.n28 plus.n27 161.3
R11 plus.n29 plus.n20 161.3
R12 plus.n31 plus.n30 161.3
R13 plus.n32 plus.n19 161.3
R14 plus.n33 plus.n18 161.3
R15 plus.n35 plus.n34 161.3
R16 plus.n5 plus.t3 113.852
R17 plus.n23 plus.t5 113.852
R18 plus.n16 plus.t7 90.5476
R19 plus.n14 plus.t2 90.5476
R20 plus.n2 plus.t6 90.5476
R21 plus.n8 plus.t0 90.5476
R22 plus.n4 plus.t8 90.5476
R23 plus.n34 plus.t1 90.5476
R24 plus.n32 plus.t11 90.5476
R25 plus.n20 plus.t10 90.5476
R26 plus.n26 plus.t9 90.5476
R27 plus.n22 plus.t4 90.5476
R28 plus.n6 plus.n5 44.8907
R29 plus.n24 plus.n23 44.8907
R30 plus.n16 plus.n15 32.8641
R31 plus.n34 plus.n33 32.8641
R32 plus.n14 plus.n13 28.4823
R33 plus.n7 plus.n4 28.4823
R34 plus.n32 plus.n31 28.4823
R35 plus.n25 plus.n22 28.4823
R36 plus plus.n35 27.1543
R37 plus.n9 plus.n8 24.1005
R38 plus.n9 plus.n2 24.1005
R39 plus.n27 plus.n20 24.1005
R40 plus.n27 plus.n26 24.1005
R41 plus.n13 plus.n2 19.7187
R42 plus.n8 plus.n7 19.7187
R43 plus.n31 plus.n20 19.7187
R44 plus.n26 plus.n25 19.7187
R45 plus.n5 plus.n4 18.4104
R46 plus.n23 plus.n22 18.4104
R47 plus.n15 plus.n14 15.3369
R48 plus.n33 plus.n32 15.3369
R49 plus plus.n17 8.12171
R50 plus.n6 plus.n3 0.189894
R51 plus.n10 plus.n3 0.189894
R52 plus.n11 plus.n10 0.189894
R53 plus.n12 plus.n11 0.189894
R54 plus.n12 plus.n1 0.189894
R55 plus.n1 plus.n0 0.189894
R56 plus.n17 plus.n0 0.189894
R57 plus.n35 plus.n18 0.189894
R58 plus.n19 plus.n18 0.189894
R59 plus.n30 plus.n19 0.189894
R60 plus.n30 plus.n29 0.189894
R61 plus.n29 plus.n28 0.189894
R62 plus.n28 plus.n21 0.189894
R63 plus.n24 plus.n21 0.189894
R64 drain_left.n6 drain_left.n4 241.02
R65 drain_left.n3 drain_left.n2 240.964
R66 drain_left.n3 drain_left.n0 240.964
R67 drain_left.n8 drain_left.n7 240.132
R68 drain_left.n6 drain_left.n5 240.132
R69 drain_left.n3 drain_left.n1 240.131
R70 drain_left drain_left.n3 23.4734
R71 drain_left.n1 drain_left.t7 19.8005
R72 drain_left.n1 drain_left.t0 19.8005
R73 drain_left.n2 drain_left.t11 19.8005
R74 drain_left.n2 drain_left.t10 19.8005
R75 drain_left.n0 drain_left.t9 19.8005
R76 drain_left.n0 drain_left.t6 19.8005
R77 drain_left.n7 drain_left.t3 19.8005
R78 drain_left.n7 drain_left.t5 19.8005
R79 drain_left.n5 drain_left.t2 19.8005
R80 drain_left.n5 drain_left.t8 19.8005
R81 drain_left.n4 drain_left.t4 19.8005
R82 drain_left.n4 drain_left.t1 19.8005
R83 drain_left drain_left.n8 6.54115
R84 drain_left.n8 drain_left.n6 0.888431
R85 source.n0 source.t16 243.255
R86 source.n5 source.t20 243.255
R87 source.n6 source.t10 243.255
R88 source.n11 source.t6 243.255
R89 source.n23 source.t0 243.254
R90 source.n18 source.t2 243.254
R91 source.n17 source.t18 243.254
R92 source.n12 source.t22 243.254
R93 source.n2 source.n1 223.454
R94 source.n4 source.n3 223.454
R95 source.n8 source.n7 223.454
R96 source.n10 source.n9 223.454
R97 source.n22 source.n21 223.453
R98 source.n20 source.n19 223.453
R99 source.n16 source.n15 223.453
R100 source.n14 source.n13 223.453
R101 source.n21 source.t1 19.8005
R102 source.n21 source.t7 19.8005
R103 source.n19 source.t11 19.8005
R104 source.n19 source.t3 19.8005
R105 source.n15 source.t14 19.8005
R106 source.n15 source.t19 19.8005
R107 source.n13 source.t12 19.8005
R108 source.n13 source.t13 19.8005
R109 source.n1 source.t17 19.8005
R110 source.n1 source.t21 19.8005
R111 source.n3 source.t15 19.8005
R112 source.n3 source.t23 19.8005
R113 source.n7 source.t8 19.8005
R114 source.n7 source.t9 19.8005
R115 source.n9 source.t4 19.8005
R116 source.n9 source.t5 19.8005
R117 source.n12 source.n11 13.8423
R118 source.n24 source.n0 8.13543
R119 source.n24 source.n23 5.7074
R120 source.n11 source.n10 0.888431
R121 source.n10 source.n8 0.888431
R122 source.n8 source.n6 0.888431
R123 source.n5 source.n4 0.888431
R124 source.n4 source.n2 0.888431
R125 source.n2 source.n0 0.888431
R126 source.n14 source.n12 0.888431
R127 source.n16 source.n14 0.888431
R128 source.n17 source.n16 0.888431
R129 source.n20 source.n18 0.888431
R130 source.n22 source.n20 0.888431
R131 source.n23 source.n22 0.888431
R132 source.n6 source.n5 0.470328
R133 source.n18 source.n17 0.470328
R134 source source.n24 0.188
R135 minus.n17 minus.n16 161.3
R136 minus.n15 minus.n0 161.3
R137 minus.n14 minus.n13 161.3
R138 minus.n12 minus.n1 161.3
R139 minus.n11 minus.n10 161.3
R140 minus.n9 minus.n2 161.3
R141 minus.n8 minus.n7 161.3
R142 minus.n6 minus.n3 161.3
R143 minus.n35 minus.n34 161.3
R144 minus.n33 minus.n18 161.3
R145 minus.n32 minus.n31 161.3
R146 minus.n30 minus.n19 161.3
R147 minus.n29 minus.n28 161.3
R148 minus.n27 minus.n20 161.3
R149 minus.n26 minus.n25 161.3
R150 minus.n24 minus.n21 161.3
R151 minus.n5 minus.t8 113.852
R152 minus.n23 minus.t2 113.852
R153 minus.n4 minus.t0 90.5476
R154 minus.n8 minus.t7 90.5476
R155 minus.n10 minus.t10 90.5476
R156 minus.n14 minus.t3 90.5476
R157 minus.n16 minus.t11 90.5476
R158 minus.n22 minus.t1 90.5476
R159 minus.n26 minus.t5 90.5476
R160 minus.n28 minus.t4 90.5476
R161 minus.n32 minus.t6 90.5476
R162 minus.n34 minus.t9 90.5476
R163 minus.n6 minus.n5 44.8907
R164 minus.n24 minus.n23 44.8907
R165 minus.n16 minus.n15 32.8641
R166 minus.n34 minus.n33 32.8641
R167 minus.n36 minus.n17 29.1066
R168 minus.n4 minus.n3 28.4823
R169 minus.n14 minus.n1 28.4823
R170 minus.n22 minus.n21 28.4823
R171 minus.n32 minus.n19 28.4823
R172 minus.n10 minus.n9 24.1005
R173 minus.n9 minus.n8 24.1005
R174 minus.n27 minus.n26 24.1005
R175 minus.n28 minus.n27 24.1005
R176 minus.n8 minus.n3 19.7187
R177 minus.n10 minus.n1 19.7187
R178 minus.n26 minus.n21 19.7187
R179 minus.n28 minus.n19 19.7187
R180 minus.n5 minus.n4 18.4104
R181 minus.n23 minus.n22 18.4104
R182 minus.n15 minus.n14 15.3369
R183 minus.n33 minus.n32 15.3369
R184 minus.n36 minus.n35 6.64444
R185 minus.n17 minus.n0 0.189894
R186 minus.n13 minus.n0 0.189894
R187 minus.n13 minus.n12 0.189894
R188 minus.n12 minus.n11 0.189894
R189 minus.n11 minus.n2 0.189894
R190 minus.n7 minus.n2 0.189894
R191 minus.n7 minus.n6 0.189894
R192 minus.n25 minus.n24 0.189894
R193 minus.n25 minus.n20 0.189894
R194 minus.n29 minus.n20 0.189894
R195 minus.n30 minus.n29 0.189894
R196 minus.n31 minus.n30 0.189894
R197 minus.n31 minus.n18 0.189894
R198 minus.n35 minus.n18 0.189894
R199 minus minus.n36 0.188
R200 drain_right.n6 drain_right.n4 241.02
R201 drain_right.n3 drain_right.n2 240.964
R202 drain_right.n3 drain_right.n0 240.964
R203 drain_right.n6 drain_right.n5 240.132
R204 drain_right.n8 drain_right.n7 240.132
R205 drain_right.n3 drain_right.n1 240.131
R206 drain_right drain_right.n3 22.9202
R207 drain_right.n1 drain_right.t6 19.8005
R208 drain_right.n1 drain_right.t7 19.8005
R209 drain_right.n2 drain_right.t5 19.8005
R210 drain_right.n2 drain_right.t2 19.8005
R211 drain_right.n0 drain_right.t9 19.8005
R212 drain_right.n0 drain_right.t10 19.8005
R213 drain_right.n4 drain_right.t11 19.8005
R214 drain_right.n4 drain_right.t3 19.8005
R215 drain_right.n5 drain_right.t1 19.8005
R216 drain_right.n5 drain_right.t4 19.8005
R217 drain_right.n7 drain_right.t0 19.8005
R218 drain_right.n7 drain_right.t8 19.8005
R219 drain_right drain_right.n8 6.54115
R220 drain_right.n8 drain_right.n6 0.888431
C0 drain_right plus 0.375212f
C1 minus drain_right 1.11541f
C2 source drain_left 3.86767f
C3 source drain_right 3.8697f
C4 minus plus 3.80715f
C5 drain_left drain_right 1.0854f
C6 source plus 1.64744f
C7 drain_left plus 1.32703f
C8 minus source 1.63358f
C9 minus drain_left 0.178985f
C10 drain_right a_n2158_n1088# 3.69623f
C11 drain_left a_n2158_n1088# 3.96417f
C12 source a_n2158_n1088# 2.581302f
C13 minus a_n2158_n1088# 7.584761f
C14 plus a_n2158_n1088# 8.188752f
C15 drain_right.t9 a_n2158_n1088# 0.015968f
C16 drain_right.t10 a_n2158_n1088# 0.015968f
C17 drain_right.n0 a_n2158_n1088# 0.062954f
C18 drain_right.t6 a_n2158_n1088# 0.015968f
C19 drain_right.t7 a_n2158_n1088# 0.015968f
C20 drain_right.n1 a_n2158_n1088# 0.062049f
C21 drain_right.t5 a_n2158_n1088# 0.015968f
C22 drain_right.t2 a_n2158_n1088# 0.015968f
C23 drain_right.n2 a_n2158_n1088# 0.062954f
C24 drain_right.n3 a_n2158_n1088# 1.30773f
C25 drain_right.t11 a_n2158_n1088# 0.015968f
C26 drain_right.t3 a_n2158_n1088# 0.015968f
C27 drain_right.n4 a_n2158_n1088# 0.063026f
C28 drain_right.t1 a_n2158_n1088# 0.015968f
C29 drain_right.t4 a_n2158_n1088# 0.015968f
C30 drain_right.n5 a_n2158_n1088# 0.062049f
C31 drain_right.n6 a_n2158_n1088# 0.521051f
C32 drain_right.t0 a_n2158_n1088# 0.015968f
C33 drain_right.t8 a_n2158_n1088# 0.015968f
C34 drain_right.n7 a_n2158_n1088# 0.062049f
C35 drain_right.n8 a_n2158_n1088# 0.43568f
C36 minus.n0 a_n2158_n1088# 0.026726f
C37 minus.n1 a_n2158_n1088# 0.006065f
C38 minus.t3 a_n2158_n1088# 0.06344f
C39 minus.n2 a_n2158_n1088# 0.026726f
C40 minus.n3 a_n2158_n1088# 0.006065f
C41 minus.t7 a_n2158_n1088# 0.06344f
C42 minus.t8 a_n2158_n1088# 0.076342f
C43 minus.t0 a_n2158_n1088# 0.06344f
C44 minus.n4 a_n2158_n1088# 0.066058f
C45 minus.n5 a_n2158_n1088# 0.052559f
C46 minus.n6 a_n2158_n1088# 0.112121f
C47 minus.n7 a_n2158_n1088# 0.026726f
C48 minus.n8 a_n2158_n1088# 0.063069f
C49 minus.n9 a_n2158_n1088# 0.006065f
C50 minus.t10 a_n2158_n1088# 0.06344f
C51 minus.n10 a_n2158_n1088# 0.063069f
C52 minus.n11 a_n2158_n1088# 0.026726f
C53 minus.n12 a_n2158_n1088# 0.026726f
C54 minus.n13 a_n2158_n1088# 0.026726f
C55 minus.n14 a_n2158_n1088# 0.063069f
C56 minus.n15 a_n2158_n1088# 0.006065f
C57 minus.t11 a_n2158_n1088# 0.06344f
C58 minus.n16 a_n2158_n1088# 0.061833f
C59 minus.n17 a_n2158_n1088# 0.663722f
C60 minus.n18 a_n2158_n1088# 0.026726f
C61 minus.n19 a_n2158_n1088# 0.006065f
C62 minus.n20 a_n2158_n1088# 0.026726f
C63 minus.n21 a_n2158_n1088# 0.006065f
C64 minus.t2 a_n2158_n1088# 0.076342f
C65 minus.t1 a_n2158_n1088# 0.06344f
C66 minus.n22 a_n2158_n1088# 0.066058f
C67 minus.n23 a_n2158_n1088# 0.052559f
C68 minus.n24 a_n2158_n1088# 0.112121f
C69 minus.n25 a_n2158_n1088# 0.026726f
C70 minus.t5 a_n2158_n1088# 0.06344f
C71 minus.n26 a_n2158_n1088# 0.063069f
C72 minus.n27 a_n2158_n1088# 0.006065f
C73 minus.t4 a_n2158_n1088# 0.06344f
C74 minus.n28 a_n2158_n1088# 0.063069f
C75 minus.n29 a_n2158_n1088# 0.026726f
C76 minus.n30 a_n2158_n1088# 0.026726f
C77 minus.n31 a_n2158_n1088# 0.026726f
C78 minus.t6 a_n2158_n1088# 0.06344f
C79 minus.n32 a_n2158_n1088# 0.063069f
C80 minus.n33 a_n2158_n1088# 0.006065f
C81 minus.t9 a_n2158_n1088# 0.06344f
C82 minus.n34 a_n2158_n1088# 0.061833f
C83 minus.n35 a_n2158_n1088# 0.183764f
C84 minus.n36 a_n2158_n1088# 0.815086f
C85 source.t16 a_n2158_n1088# 0.105408f
C86 source.n0 a_n2158_n1088# 0.500157f
C87 source.t17 a_n2158_n1088# 0.018938f
C88 source.t21 a_n2158_n1088# 0.018938f
C89 source.n1 a_n2158_n1088# 0.06142f
C90 source.n2 a_n2158_n1088# 0.284324f
C91 source.t15 a_n2158_n1088# 0.018938f
C92 source.t23 a_n2158_n1088# 0.018938f
C93 source.n3 a_n2158_n1088# 0.06142f
C94 source.n4 a_n2158_n1088# 0.284324f
C95 source.t20 a_n2158_n1088# 0.105408f
C96 source.n5 a_n2158_n1088# 0.259699f
C97 source.t10 a_n2158_n1088# 0.105408f
C98 source.n6 a_n2158_n1088# 0.259699f
C99 source.t8 a_n2158_n1088# 0.018938f
C100 source.t9 a_n2158_n1088# 0.018938f
C101 source.n7 a_n2158_n1088# 0.06142f
C102 source.n8 a_n2158_n1088# 0.284324f
C103 source.t4 a_n2158_n1088# 0.018938f
C104 source.t5 a_n2158_n1088# 0.018938f
C105 source.n9 a_n2158_n1088# 0.06142f
C106 source.n10 a_n2158_n1088# 0.284324f
C107 source.t6 a_n2158_n1088# 0.105408f
C108 source.n11 a_n2158_n1088# 0.697897f
C109 source.t22 a_n2158_n1088# 0.105408f
C110 source.n12 a_n2158_n1088# 0.697897f
C111 source.t12 a_n2158_n1088# 0.018938f
C112 source.t13 a_n2158_n1088# 0.018938f
C113 source.n13 a_n2158_n1088# 0.06142f
C114 source.n14 a_n2158_n1088# 0.284324f
C115 source.t14 a_n2158_n1088# 0.018938f
C116 source.t19 a_n2158_n1088# 0.018938f
C117 source.n15 a_n2158_n1088# 0.06142f
C118 source.n16 a_n2158_n1088# 0.284324f
C119 source.t18 a_n2158_n1088# 0.105408f
C120 source.n17 a_n2158_n1088# 0.259699f
C121 source.t2 a_n2158_n1088# 0.105408f
C122 source.n18 a_n2158_n1088# 0.259699f
C123 source.t11 a_n2158_n1088# 0.018938f
C124 source.t3 a_n2158_n1088# 0.018938f
C125 source.n19 a_n2158_n1088# 0.06142f
C126 source.n20 a_n2158_n1088# 0.284324f
C127 source.t1 a_n2158_n1088# 0.018938f
C128 source.t7 a_n2158_n1088# 0.018938f
C129 source.n21 a_n2158_n1088# 0.06142f
C130 source.n22 a_n2158_n1088# 0.284324f
C131 source.t0 a_n2158_n1088# 0.105408f
C132 source.n23 a_n2158_n1088# 0.416027f
C133 source.n24 a_n2158_n1088# 0.496656f
C134 drain_left.t9 a_n2158_n1088# 0.015651f
C135 drain_left.t6 a_n2158_n1088# 0.015651f
C136 drain_left.n0 a_n2158_n1088# 0.061704f
C137 drain_left.t7 a_n2158_n1088# 0.015651f
C138 drain_left.t0 a_n2158_n1088# 0.015651f
C139 drain_left.n1 a_n2158_n1088# 0.060816f
C140 drain_left.t11 a_n2158_n1088# 0.015651f
C141 drain_left.t10 a_n2158_n1088# 0.015651f
C142 drain_left.n2 a_n2158_n1088# 0.061704f
C143 drain_left.n3 a_n2158_n1088# 1.31995f
C144 drain_left.t4 a_n2158_n1088# 0.015651f
C145 drain_left.t1 a_n2158_n1088# 0.015651f
C146 drain_left.n4 a_n2158_n1088# 0.061773f
C147 drain_left.t2 a_n2158_n1088# 0.015651f
C148 drain_left.t8 a_n2158_n1088# 0.015651f
C149 drain_left.n5 a_n2158_n1088# 0.060816f
C150 drain_left.n6 a_n2158_n1088# 0.5107f
C151 drain_left.t3 a_n2158_n1088# 0.015651f
C152 drain_left.t5 a_n2158_n1088# 0.015651f
C153 drain_left.n7 a_n2158_n1088# 0.060816f
C154 drain_left.n8 a_n2158_n1088# 0.427025f
C155 plus.n0 a_n2158_n1088# 0.027112f
C156 plus.t7 a_n2158_n1088# 0.064356f
C157 plus.t2 a_n2158_n1088# 0.064356f
C158 plus.n1 a_n2158_n1088# 0.027112f
C159 plus.t6 a_n2158_n1088# 0.064356f
C160 plus.n2 a_n2158_n1088# 0.063979f
C161 plus.n3 a_n2158_n1088# 0.027112f
C162 plus.t0 a_n2158_n1088# 0.064356f
C163 plus.t8 a_n2158_n1088# 0.064356f
C164 plus.n4 a_n2158_n1088# 0.067011f
C165 plus.t3 a_n2158_n1088# 0.077444f
C166 plus.n5 a_n2158_n1088# 0.053318f
C167 plus.n6 a_n2158_n1088# 0.113738f
C168 plus.n7 a_n2158_n1088# 0.006152f
C169 plus.n8 a_n2158_n1088# 0.063979f
C170 plus.n9 a_n2158_n1088# 0.006152f
C171 plus.n10 a_n2158_n1088# 0.027112f
C172 plus.n11 a_n2158_n1088# 0.027112f
C173 plus.n12 a_n2158_n1088# 0.027112f
C174 plus.n13 a_n2158_n1088# 0.006152f
C175 plus.n14 a_n2158_n1088# 0.063979f
C176 plus.n15 a_n2158_n1088# 0.006152f
C177 plus.n16 a_n2158_n1088# 0.062725f
C178 plus.n17 a_n2158_n1088# 0.195543f
C179 plus.n18 a_n2158_n1088# 0.027112f
C180 plus.t1 a_n2158_n1088# 0.064356f
C181 plus.n19 a_n2158_n1088# 0.027112f
C182 plus.t11 a_n2158_n1088# 0.064356f
C183 plus.t10 a_n2158_n1088# 0.064356f
C184 plus.n20 a_n2158_n1088# 0.063979f
C185 plus.n21 a_n2158_n1088# 0.027112f
C186 plus.t9 a_n2158_n1088# 0.064356f
C187 plus.t4 a_n2158_n1088# 0.064356f
C188 plus.n22 a_n2158_n1088# 0.067011f
C189 plus.t5 a_n2158_n1088# 0.077444f
C190 plus.n23 a_n2158_n1088# 0.053318f
C191 plus.n24 a_n2158_n1088# 0.113738f
C192 plus.n25 a_n2158_n1088# 0.006152f
C193 plus.n26 a_n2158_n1088# 0.063979f
C194 plus.n27 a_n2158_n1088# 0.006152f
C195 plus.n28 a_n2158_n1088# 0.027112f
C196 plus.n29 a_n2158_n1088# 0.027112f
C197 plus.n30 a_n2158_n1088# 0.027112f
C198 plus.n31 a_n2158_n1088# 0.006152f
C199 plus.n32 a_n2158_n1088# 0.063979f
C200 plus.n33 a_n2158_n1088# 0.006152f
C201 plus.n34 a_n2158_n1088# 0.062725f
C202 plus.n35 a_n2158_n1088# 0.651222f
.ends

