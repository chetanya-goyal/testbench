* NGSPICE file created from diffpair266.ext - technology: sky130A

.subckt diffpair266 minus drain_right drain_left source plus
X0 source.t27 plus.t0 drain_left.t12 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X1 source.t26 plus.t1 drain_left.t2 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X2 drain_left.t13 plus.t2 source.t25 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X3 source.t7 minus.t0 drain_right.t13 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X4 source.t10 minus.t1 drain_right.t12 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X5 drain_left.t7 plus.t3 source.t24 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X6 a_n1644_n2088# a_n1644_n2088# a_n1644_n2088# a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.25
X7 source.t5 minus.t2 drain_right.t11 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X8 drain_left.t8 plus.t4 source.t23 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X9 source.t6 minus.t3 drain_right.t10 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X10 drain_right.t9 minus.t4 source.t13 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X11 source.t22 plus.t5 drain_left.t9 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X12 drain_right.t8 minus.t5 source.t8 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X13 source.t21 plus.t6 drain_left.t10 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X14 drain_left.t0 plus.t7 source.t20 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X15 drain_left.t3 plus.t8 source.t19 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X16 drain_left.t1 plus.t9 source.t18 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X17 drain_left.t6 plus.t10 source.t17 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X18 source.t3 minus.t6 drain_right.t7 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X19 drain_right.t6 minus.t7 source.t4 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X20 drain_right.t5 minus.t8 source.t9 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X21 drain_right.t4 minus.t9 source.t11 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X22 source.t16 plus.t11 drain_left.t11 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X23 a_n1644_n2088# a_n1644_n2088# a_n1644_n2088# a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X24 a_n1644_n2088# a_n1644_n2088# a_n1644_n2088# a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X25 source.t0 minus.t10 drain_right.t3 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X26 drain_left.t4 plus.t12 source.t15 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X27 drain_right.t2 minus.t11 source.t12 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X28 drain_right.t1 minus.t12 source.t2 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X29 drain_right.t0 minus.t13 source.t1 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X30 source.t14 plus.t13 drain_left.t5 a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X31 a_n1644_n2088# a_n1644_n2088# a_n1644_n2088# a_n1644_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
R0 plus.n3 plus.t3 738.775
R1 plus.n15 plus.t7 738.775
R2 plus.n20 plus.t10 738.775
R3 plus.n32 plus.t4 738.775
R4 plus.n1 plus.t0 703.721
R5 plus.n4 plus.t1 703.721
R6 plus.n6 plus.t9 703.721
R7 plus.n12 plus.t8 703.721
R8 plus.n14 plus.t13 703.721
R9 plus.n18 plus.t11 703.721
R10 plus.n21 plus.t5 703.721
R11 plus.n23 plus.t2 703.721
R12 plus.n29 plus.t12 703.721
R13 plus.n31 plus.t6 703.721
R14 plus.n3 plus.n2 161.489
R15 plus.n20 plus.n19 161.489
R16 plus.n5 plus.n2 161.3
R17 plus.n8 plus.n7 161.3
R18 plus.n9 plus.n1 161.3
R19 plus.n11 plus.n10 161.3
R20 plus.n13 plus.n0 161.3
R21 plus.n16 plus.n15 161.3
R22 plus.n22 plus.n19 161.3
R23 plus.n25 plus.n24 161.3
R24 plus.n26 plus.n18 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n17 161.3
R27 plus.n33 plus.n32 161.3
R28 plus.n7 plus.n1 73.0308
R29 plus.n11 plus.n1 73.0308
R30 plus.n28 plus.n18 73.0308
R31 plus.n24 plus.n18 73.0308
R32 plus.n6 plus.n5 61.346
R33 plus.n13 plus.n12 61.346
R34 plus.n30 plus.n29 61.346
R35 plus.n23 plus.n22 61.346
R36 plus.n4 plus.n3 49.6611
R37 plus.n15 plus.n14 49.6611
R38 plus.n32 plus.n31 49.6611
R39 plus.n21 plus.n20 49.6611
R40 plus plus.n33 26.9081
R41 plus.n5 plus.n4 23.3702
R42 plus.n14 plus.n13 23.3702
R43 plus.n31 plus.n30 23.3702
R44 plus.n22 plus.n21 23.3702
R45 plus.n7 plus.n6 11.6853
R46 plus.n12 plus.n11 11.6853
R47 plus.n29 plus.n28 11.6853
R48 plus.n24 plus.n23 11.6853
R49 plus plus.n16 9.82247
R50 plus.n8 plus.n2 0.189894
R51 plus.n9 plus.n8 0.189894
R52 plus.n10 plus.n9 0.189894
R53 plus.n10 plus.n0 0.189894
R54 plus.n16 plus.n0 0.189894
R55 plus.n33 plus.n17 0.189894
R56 plus.n27 plus.n17 0.189894
R57 plus.n27 plus.n26 0.189894
R58 plus.n26 plus.n25 0.189894
R59 plus.n25 plus.n19 0.189894
R60 drain_left.n26 drain_left.n0 289.615
R61 drain_left.n63 drain_left.n37 289.615
R62 drain_left.n11 drain_left.n10 185
R63 drain_left.n8 drain_left.n7 185
R64 drain_left.n17 drain_left.n16 185
R65 drain_left.n19 drain_left.n18 185
R66 drain_left.n4 drain_left.n3 185
R67 drain_left.n25 drain_left.n24 185
R68 drain_left.n27 drain_left.n26 185
R69 drain_left.n64 drain_left.n63 185
R70 drain_left.n62 drain_left.n61 185
R71 drain_left.n41 drain_left.n40 185
R72 drain_left.n56 drain_left.n55 185
R73 drain_left.n54 drain_left.n53 185
R74 drain_left.n45 drain_left.n44 185
R75 drain_left.n48 drain_left.n47 185
R76 drain_left.t8 drain_left.n9 147.661
R77 drain_left.t7 drain_left.n46 147.661
R78 drain_left.n10 drain_left.n7 104.615
R79 drain_left.n17 drain_left.n7 104.615
R80 drain_left.n18 drain_left.n17 104.615
R81 drain_left.n18 drain_left.n3 104.615
R82 drain_left.n25 drain_left.n3 104.615
R83 drain_left.n26 drain_left.n25 104.615
R84 drain_left.n63 drain_left.n62 104.615
R85 drain_left.n62 drain_left.n40 104.615
R86 drain_left.n55 drain_left.n40 104.615
R87 drain_left.n55 drain_left.n54 104.615
R88 drain_left.n54 drain_left.n44 104.615
R89 drain_left.n47 drain_left.n44 104.615
R90 drain_left.n35 drain_left.n33 67.6907
R91 drain_left.n71 drain_left.n70 67.1908
R92 drain_left.n69 drain_left.n68 67.1908
R93 drain_left.n73 drain_left.n72 67.1907
R94 drain_left.n35 drain_left.n34 67.1907
R95 drain_left.n32 drain_left.n31 67.1907
R96 drain_left.n10 drain_left.t8 52.3082
R97 drain_left.n47 drain_left.t7 52.3082
R98 drain_left.n32 drain_left.n30 49.3641
R99 drain_left.n69 drain_left.n67 49.3641
R100 drain_left drain_left.n36 25.6966
R101 drain_left.n11 drain_left.n9 15.6674
R102 drain_left.n48 drain_left.n46 15.6674
R103 drain_left.n12 drain_left.n8 12.8005
R104 drain_left.n49 drain_left.n45 12.8005
R105 drain_left.n16 drain_left.n15 12.0247
R106 drain_left.n53 drain_left.n52 12.0247
R107 drain_left.n19 drain_left.n6 11.249
R108 drain_left.n56 drain_left.n43 11.249
R109 drain_left.n20 drain_left.n4 10.4732
R110 drain_left.n57 drain_left.n41 10.4732
R111 drain_left.n24 drain_left.n23 9.69747
R112 drain_left.n61 drain_left.n60 9.69747
R113 drain_left.n30 drain_left.n29 9.45567
R114 drain_left.n67 drain_left.n66 9.45567
R115 drain_left.n29 drain_left.n28 9.3005
R116 drain_left.n2 drain_left.n1 9.3005
R117 drain_left.n23 drain_left.n22 9.3005
R118 drain_left.n21 drain_left.n20 9.3005
R119 drain_left.n6 drain_left.n5 9.3005
R120 drain_left.n15 drain_left.n14 9.3005
R121 drain_left.n13 drain_left.n12 9.3005
R122 drain_left.n66 drain_left.n65 9.3005
R123 drain_left.n39 drain_left.n38 9.3005
R124 drain_left.n60 drain_left.n59 9.3005
R125 drain_left.n58 drain_left.n57 9.3005
R126 drain_left.n43 drain_left.n42 9.3005
R127 drain_left.n52 drain_left.n51 9.3005
R128 drain_left.n50 drain_left.n49 9.3005
R129 drain_left.n27 drain_left.n2 8.92171
R130 drain_left.n64 drain_left.n39 8.92171
R131 drain_left.n28 drain_left.n0 8.14595
R132 drain_left.n65 drain_left.n37 8.14595
R133 drain_left drain_left.n73 6.15322
R134 drain_left.n30 drain_left.n0 5.81868
R135 drain_left.n67 drain_left.n37 5.81868
R136 drain_left.n28 drain_left.n27 5.04292
R137 drain_left.n65 drain_left.n64 5.04292
R138 drain_left.n13 drain_left.n9 4.38594
R139 drain_left.n50 drain_left.n46 4.38594
R140 drain_left.n24 drain_left.n2 4.26717
R141 drain_left.n61 drain_left.n39 4.26717
R142 drain_left.n23 drain_left.n4 3.49141
R143 drain_left.n60 drain_left.n41 3.49141
R144 drain_left.n33 drain_left.t9 3.3005
R145 drain_left.n33 drain_left.t6 3.3005
R146 drain_left.n34 drain_left.t11 3.3005
R147 drain_left.n34 drain_left.t13 3.3005
R148 drain_left.n31 drain_left.t10 3.3005
R149 drain_left.n31 drain_left.t4 3.3005
R150 drain_left.n72 drain_left.t5 3.3005
R151 drain_left.n72 drain_left.t0 3.3005
R152 drain_left.n70 drain_left.t12 3.3005
R153 drain_left.n70 drain_left.t3 3.3005
R154 drain_left.n68 drain_left.t2 3.3005
R155 drain_left.n68 drain_left.t1 3.3005
R156 drain_left.n20 drain_left.n19 2.71565
R157 drain_left.n57 drain_left.n56 2.71565
R158 drain_left.n16 drain_left.n6 1.93989
R159 drain_left.n53 drain_left.n43 1.93989
R160 drain_left.n15 drain_left.n8 1.16414
R161 drain_left.n52 drain_left.n45 1.16414
R162 drain_left.n71 drain_left.n69 0.5005
R163 drain_left.n73 drain_left.n71 0.5005
R164 drain_left.n12 drain_left.n11 0.388379
R165 drain_left.n49 drain_left.n48 0.388379
R166 drain_left.n36 drain_left.n32 0.320154
R167 drain_left.n14 drain_left.n13 0.155672
R168 drain_left.n14 drain_left.n5 0.155672
R169 drain_left.n21 drain_left.n5 0.155672
R170 drain_left.n22 drain_left.n21 0.155672
R171 drain_left.n22 drain_left.n1 0.155672
R172 drain_left.n29 drain_left.n1 0.155672
R173 drain_left.n66 drain_left.n38 0.155672
R174 drain_left.n59 drain_left.n38 0.155672
R175 drain_left.n59 drain_left.n58 0.155672
R176 drain_left.n58 drain_left.n42 0.155672
R177 drain_left.n51 drain_left.n42 0.155672
R178 drain_left.n51 drain_left.n50 0.155672
R179 drain_left.n36 drain_left.n35 0.070154
R180 source.n146 source.n120 289.615
R181 source.n108 source.n82 289.615
R182 source.n26 source.n0 289.615
R183 source.n64 source.n38 289.615
R184 source.n131 source.n130 185
R185 source.n128 source.n127 185
R186 source.n137 source.n136 185
R187 source.n139 source.n138 185
R188 source.n124 source.n123 185
R189 source.n145 source.n144 185
R190 source.n147 source.n146 185
R191 source.n93 source.n92 185
R192 source.n90 source.n89 185
R193 source.n99 source.n98 185
R194 source.n101 source.n100 185
R195 source.n86 source.n85 185
R196 source.n107 source.n106 185
R197 source.n109 source.n108 185
R198 source.n27 source.n26 185
R199 source.n25 source.n24 185
R200 source.n4 source.n3 185
R201 source.n19 source.n18 185
R202 source.n17 source.n16 185
R203 source.n8 source.n7 185
R204 source.n11 source.n10 185
R205 source.n65 source.n64 185
R206 source.n63 source.n62 185
R207 source.n42 source.n41 185
R208 source.n57 source.n56 185
R209 source.n55 source.n54 185
R210 source.n46 source.n45 185
R211 source.n49 source.n48 185
R212 source.t13 source.n129 147.661
R213 source.t17 source.n91 147.661
R214 source.t20 source.n9 147.661
R215 source.t11 source.n47 147.661
R216 source.n130 source.n127 104.615
R217 source.n137 source.n127 104.615
R218 source.n138 source.n137 104.615
R219 source.n138 source.n123 104.615
R220 source.n145 source.n123 104.615
R221 source.n146 source.n145 104.615
R222 source.n92 source.n89 104.615
R223 source.n99 source.n89 104.615
R224 source.n100 source.n99 104.615
R225 source.n100 source.n85 104.615
R226 source.n107 source.n85 104.615
R227 source.n108 source.n107 104.615
R228 source.n26 source.n25 104.615
R229 source.n25 source.n3 104.615
R230 source.n18 source.n3 104.615
R231 source.n18 source.n17 104.615
R232 source.n17 source.n7 104.615
R233 source.n10 source.n7 104.615
R234 source.n64 source.n63 104.615
R235 source.n63 source.n41 104.615
R236 source.n56 source.n41 104.615
R237 source.n56 source.n55 104.615
R238 source.n55 source.n45 104.615
R239 source.n48 source.n45 104.615
R240 source.n130 source.t13 52.3082
R241 source.n92 source.t17 52.3082
R242 source.n10 source.t20 52.3082
R243 source.n48 source.t11 52.3082
R244 source.n33 source.n32 50.512
R245 source.n35 source.n34 50.512
R246 source.n37 source.n36 50.512
R247 source.n71 source.n70 50.512
R248 source.n73 source.n72 50.512
R249 source.n75 source.n74 50.512
R250 source.n119 source.n118 50.5119
R251 source.n117 source.n116 50.5119
R252 source.n115 source.n114 50.5119
R253 source.n81 source.n80 50.5119
R254 source.n79 source.n78 50.5119
R255 source.n77 source.n76 50.5119
R256 source.n151 source.n150 32.1853
R257 source.n113 source.n112 32.1853
R258 source.n31 source.n30 32.1853
R259 source.n69 source.n68 32.1853
R260 source.n77 source.n75 17.7423
R261 source.n131 source.n129 15.6674
R262 source.n93 source.n91 15.6674
R263 source.n11 source.n9 15.6674
R264 source.n49 source.n47 15.6674
R265 source.n132 source.n128 12.8005
R266 source.n94 source.n90 12.8005
R267 source.n12 source.n8 12.8005
R268 source.n50 source.n46 12.8005
R269 source.n136 source.n135 12.0247
R270 source.n98 source.n97 12.0247
R271 source.n16 source.n15 12.0247
R272 source.n54 source.n53 12.0247
R273 source.n152 source.n31 11.7293
R274 source.n139 source.n126 11.249
R275 source.n101 source.n88 11.249
R276 source.n19 source.n6 11.249
R277 source.n57 source.n44 11.249
R278 source.n140 source.n124 10.4732
R279 source.n102 source.n86 10.4732
R280 source.n20 source.n4 10.4732
R281 source.n58 source.n42 10.4732
R282 source.n144 source.n143 9.69747
R283 source.n106 source.n105 9.69747
R284 source.n24 source.n23 9.69747
R285 source.n62 source.n61 9.69747
R286 source.n150 source.n149 9.45567
R287 source.n112 source.n111 9.45567
R288 source.n30 source.n29 9.45567
R289 source.n68 source.n67 9.45567
R290 source.n149 source.n148 9.3005
R291 source.n122 source.n121 9.3005
R292 source.n143 source.n142 9.3005
R293 source.n141 source.n140 9.3005
R294 source.n126 source.n125 9.3005
R295 source.n135 source.n134 9.3005
R296 source.n133 source.n132 9.3005
R297 source.n111 source.n110 9.3005
R298 source.n84 source.n83 9.3005
R299 source.n105 source.n104 9.3005
R300 source.n103 source.n102 9.3005
R301 source.n88 source.n87 9.3005
R302 source.n97 source.n96 9.3005
R303 source.n95 source.n94 9.3005
R304 source.n29 source.n28 9.3005
R305 source.n2 source.n1 9.3005
R306 source.n23 source.n22 9.3005
R307 source.n21 source.n20 9.3005
R308 source.n6 source.n5 9.3005
R309 source.n15 source.n14 9.3005
R310 source.n13 source.n12 9.3005
R311 source.n67 source.n66 9.3005
R312 source.n40 source.n39 9.3005
R313 source.n61 source.n60 9.3005
R314 source.n59 source.n58 9.3005
R315 source.n44 source.n43 9.3005
R316 source.n53 source.n52 9.3005
R317 source.n51 source.n50 9.3005
R318 source.n147 source.n122 8.92171
R319 source.n109 source.n84 8.92171
R320 source.n27 source.n2 8.92171
R321 source.n65 source.n40 8.92171
R322 source.n148 source.n120 8.14595
R323 source.n110 source.n82 8.14595
R324 source.n28 source.n0 8.14595
R325 source.n66 source.n38 8.14595
R326 source.n150 source.n120 5.81868
R327 source.n112 source.n82 5.81868
R328 source.n30 source.n0 5.81868
R329 source.n68 source.n38 5.81868
R330 source.n152 source.n151 5.51343
R331 source.n148 source.n147 5.04292
R332 source.n110 source.n109 5.04292
R333 source.n28 source.n27 5.04292
R334 source.n66 source.n65 5.04292
R335 source.n133 source.n129 4.38594
R336 source.n95 source.n91 4.38594
R337 source.n13 source.n9 4.38594
R338 source.n51 source.n47 4.38594
R339 source.n144 source.n122 4.26717
R340 source.n106 source.n84 4.26717
R341 source.n24 source.n2 4.26717
R342 source.n62 source.n40 4.26717
R343 source.n143 source.n124 3.49141
R344 source.n105 source.n86 3.49141
R345 source.n23 source.n4 3.49141
R346 source.n61 source.n42 3.49141
R347 source.n118 source.t1 3.3005
R348 source.n118 source.t3 3.3005
R349 source.n116 source.t8 3.3005
R350 source.n116 source.t5 3.3005
R351 source.n114 source.t9 3.3005
R352 source.n114 source.t0 3.3005
R353 source.n80 source.t25 3.3005
R354 source.n80 source.t22 3.3005
R355 source.n78 source.t15 3.3005
R356 source.n78 source.t16 3.3005
R357 source.n76 source.t23 3.3005
R358 source.n76 source.t21 3.3005
R359 source.n32 source.t19 3.3005
R360 source.n32 source.t14 3.3005
R361 source.n34 source.t18 3.3005
R362 source.n34 source.t27 3.3005
R363 source.n36 source.t24 3.3005
R364 source.n36 source.t26 3.3005
R365 source.n70 source.t4 3.3005
R366 source.n70 source.t10 3.3005
R367 source.n72 source.t12 3.3005
R368 source.n72 source.t7 3.3005
R369 source.n74 source.t2 3.3005
R370 source.n74 source.t6 3.3005
R371 source.n140 source.n139 2.71565
R372 source.n102 source.n101 2.71565
R373 source.n20 source.n19 2.71565
R374 source.n58 source.n57 2.71565
R375 source.n136 source.n126 1.93989
R376 source.n98 source.n88 1.93989
R377 source.n16 source.n6 1.93989
R378 source.n54 source.n44 1.93989
R379 source.n135 source.n128 1.16414
R380 source.n97 source.n90 1.16414
R381 source.n15 source.n8 1.16414
R382 source.n53 source.n46 1.16414
R383 source.n69 source.n37 0.720328
R384 source.n115 source.n113 0.720328
R385 source.n75 source.n73 0.5005
R386 source.n73 source.n71 0.5005
R387 source.n71 source.n69 0.5005
R388 source.n37 source.n35 0.5005
R389 source.n35 source.n33 0.5005
R390 source.n33 source.n31 0.5005
R391 source.n79 source.n77 0.5005
R392 source.n81 source.n79 0.5005
R393 source.n113 source.n81 0.5005
R394 source.n117 source.n115 0.5005
R395 source.n119 source.n117 0.5005
R396 source.n151 source.n119 0.5005
R397 source.n132 source.n131 0.388379
R398 source.n94 source.n93 0.388379
R399 source.n12 source.n11 0.388379
R400 source.n50 source.n49 0.388379
R401 source source.n152 0.188
R402 source.n134 source.n133 0.155672
R403 source.n134 source.n125 0.155672
R404 source.n141 source.n125 0.155672
R405 source.n142 source.n141 0.155672
R406 source.n142 source.n121 0.155672
R407 source.n149 source.n121 0.155672
R408 source.n96 source.n95 0.155672
R409 source.n96 source.n87 0.155672
R410 source.n103 source.n87 0.155672
R411 source.n104 source.n103 0.155672
R412 source.n104 source.n83 0.155672
R413 source.n111 source.n83 0.155672
R414 source.n29 source.n1 0.155672
R415 source.n22 source.n1 0.155672
R416 source.n22 source.n21 0.155672
R417 source.n21 source.n5 0.155672
R418 source.n14 source.n5 0.155672
R419 source.n14 source.n13 0.155672
R420 source.n67 source.n39 0.155672
R421 source.n60 source.n39 0.155672
R422 source.n60 source.n59 0.155672
R423 source.n59 source.n43 0.155672
R424 source.n52 source.n43 0.155672
R425 source.n52 source.n51 0.155672
R426 minus.n15 minus.t12 738.775
R427 minus.n3 minus.t9 738.775
R428 minus.n32 minus.t4 738.775
R429 minus.n20 minus.t8 738.775
R430 minus.n1 minus.t0 703.721
R431 minus.n14 minus.t3 703.721
R432 minus.n12 minus.t11 703.721
R433 minus.n6 minus.t7 703.721
R434 minus.n4 minus.t1 703.721
R435 minus.n18 minus.t2 703.721
R436 minus.n31 minus.t6 703.721
R437 minus.n29 minus.t13 703.721
R438 minus.n23 minus.t5 703.721
R439 minus.n21 minus.t10 703.721
R440 minus.n3 minus.n2 161.489
R441 minus.n20 minus.n19 161.489
R442 minus.n16 minus.n15 161.3
R443 minus.n13 minus.n0 161.3
R444 minus.n11 minus.n10 161.3
R445 minus.n9 minus.n1 161.3
R446 minus.n8 minus.n7 161.3
R447 minus.n5 minus.n2 161.3
R448 minus.n33 minus.n32 161.3
R449 minus.n30 minus.n17 161.3
R450 minus.n28 minus.n27 161.3
R451 minus.n26 minus.n18 161.3
R452 minus.n25 minus.n24 161.3
R453 minus.n22 minus.n19 161.3
R454 minus.n11 minus.n1 73.0308
R455 minus.n7 minus.n1 73.0308
R456 minus.n24 minus.n18 73.0308
R457 minus.n28 minus.n18 73.0308
R458 minus.n13 minus.n12 61.346
R459 minus.n6 minus.n5 61.346
R460 minus.n23 minus.n22 61.346
R461 minus.n30 minus.n29 61.346
R462 minus.n15 minus.n14 49.6611
R463 minus.n4 minus.n3 49.6611
R464 minus.n21 minus.n20 49.6611
R465 minus.n32 minus.n31 49.6611
R466 minus.n34 minus.n16 30.7543
R467 minus.n14 minus.n13 23.3702
R468 minus.n5 minus.n4 23.3702
R469 minus.n22 minus.n21 23.3702
R470 minus.n31 minus.n30 23.3702
R471 minus.n12 minus.n11 11.6853
R472 minus.n7 minus.n6 11.6853
R473 minus.n24 minus.n23 11.6853
R474 minus.n29 minus.n28 11.6853
R475 minus.n34 minus.n33 6.45126
R476 minus.n16 minus.n0 0.189894
R477 minus.n10 minus.n0 0.189894
R478 minus.n10 minus.n9 0.189894
R479 minus.n9 minus.n8 0.189894
R480 minus.n8 minus.n2 0.189894
R481 minus.n25 minus.n19 0.189894
R482 minus.n26 minus.n25 0.189894
R483 minus.n27 minus.n26 0.189894
R484 minus.n27 minus.n17 0.189894
R485 minus.n33 minus.n17 0.189894
R486 minus minus.n34 0.188
R487 drain_right.n26 drain_right.n0 289.615
R488 drain_right.n68 drain_right.n42 289.615
R489 drain_right.n11 drain_right.n10 185
R490 drain_right.n8 drain_right.n7 185
R491 drain_right.n17 drain_right.n16 185
R492 drain_right.n19 drain_right.n18 185
R493 drain_right.n4 drain_right.n3 185
R494 drain_right.n25 drain_right.n24 185
R495 drain_right.n27 drain_right.n26 185
R496 drain_right.n69 drain_right.n68 185
R497 drain_right.n67 drain_right.n66 185
R498 drain_right.n46 drain_right.n45 185
R499 drain_right.n61 drain_right.n60 185
R500 drain_right.n59 drain_right.n58 185
R501 drain_right.n50 drain_right.n49 185
R502 drain_right.n53 drain_right.n52 185
R503 drain_right.t5 drain_right.n9 147.661
R504 drain_right.t1 drain_right.n51 147.661
R505 drain_right.n10 drain_right.n7 104.615
R506 drain_right.n17 drain_right.n7 104.615
R507 drain_right.n18 drain_right.n17 104.615
R508 drain_right.n18 drain_right.n3 104.615
R509 drain_right.n25 drain_right.n3 104.615
R510 drain_right.n26 drain_right.n25 104.615
R511 drain_right.n68 drain_right.n67 104.615
R512 drain_right.n67 drain_right.n45 104.615
R513 drain_right.n60 drain_right.n45 104.615
R514 drain_right.n60 drain_right.n59 104.615
R515 drain_right.n59 drain_right.n49 104.615
R516 drain_right.n52 drain_right.n49 104.615
R517 drain_right.n39 drain_right.n37 67.6907
R518 drain_right.n35 drain_right.n33 67.6907
R519 drain_right.n39 drain_right.n38 67.1908
R520 drain_right.n41 drain_right.n40 67.1908
R521 drain_right.n35 drain_right.n34 67.1907
R522 drain_right.n32 drain_right.n31 67.1907
R523 drain_right.n10 drain_right.t5 52.3082
R524 drain_right.n52 drain_right.t1 52.3082
R525 drain_right.n32 drain_right.n30 49.3641
R526 drain_right.n73 drain_right.n72 48.8641
R527 drain_right drain_right.n36 25.1434
R528 drain_right.n11 drain_right.n9 15.6674
R529 drain_right.n53 drain_right.n51 15.6674
R530 drain_right.n12 drain_right.n8 12.8005
R531 drain_right.n54 drain_right.n50 12.8005
R532 drain_right.n16 drain_right.n15 12.0247
R533 drain_right.n58 drain_right.n57 12.0247
R534 drain_right.n19 drain_right.n6 11.249
R535 drain_right.n61 drain_right.n48 11.249
R536 drain_right.n20 drain_right.n4 10.4732
R537 drain_right.n62 drain_right.n46 10.4732
R538 drain_right.n24 drain_right.n23 9.69747
R539 drain_right.n66 drain_right.n65 9.69747
R540 drain_right.n30 drain_right.n29 9.45567
R541 drain_right.n72 drain_right.n71 9.45567
R542 drain_right.n29 drain_right.n28 9.3005
R543 drain_right.n2 drain_right.n1 9.3005
R544 drain_right.n23 drain_right.n22 9.3005
R545 drain_right.n21 drain_right.n20 9.3005
R546 drain_right.n6 drain_right.n5 9.3005
R547 drain_right.n15 drain_right.n14 9.3005
R548 drain_right.n13 drain_right.n12 9.3005
R549 drain_right.n71 drain_right.n70 9.3005
R550 drain_right.n44 drain_right.n43 9.3005
R551 drain_right.n65 drain_right.n64 9.3005
R552 drain_right.n63 drain_right.n62 9.3005
R553 drain_right.n48 drain_right.n47 9.3005
R554 drain_right.n57 drain_right.n56 9.3005
R555 drain_right.n55 drain_right.n54 9.3005
R556 drain_right.n27 drain_right.n2 8.92171
R557 drain_right.n69 drain_right.n44 8.92171
R558 drain_right.n28 drain_right.n0 8.14595
R559 drain_right.n70 drain_right.n42 8.14595
R560 drain_right drain_right.n73 5.90322
R561 drain_right.n30 drain_right.n0 5.81868
R562 drain_right.n72 drain_right.n42 5.81868
R563 drain_right.n28 drain_right.n27 5.04292
R564 drain_right.n70 drain_right.n69 5.04292
R565 drain_right.n13 drain_right.n9 4.38594
R566 drain_right.n55 drain_right.n51 4.38594
R567 drain_right.n24 drain_right.n2 4.26717
R568 drain_right.n66 drain_right.n44 4.26717
R569 drain_right.n23 drain_right.n4 3.49141
R570 drain_right.n65 drain_right.n46 3.49141
R571 drain_right.n33 drain_right.t7 3.3005
R572 drain_right.n33 drain_right.t9 3.3005
R573 drain_right.n34 drain_right.t11 3.3005
R574 drain_right.n34 drain_right.t0 3.3005
R575 drain_right.n31 drain_right.t3 3.3005
R576 drain_right.n31 drain_right.t8 3.3005
R577 drain_right.n37 drain_right.t12 3.3005
R578 drain_right.n37 drain_right.t4 3.3005
R579 drain_right.n38 drain_right.t13 3.3005
R580 drain_right.n38 drain_right.t6 3.3005
R581 drain_right.n40 drain_right.t10 3.3005
R582 drain_right.n40 drain_right.t2 3.3005
R583 drain_right.n20 drain_right.n19 2.71565
R584 drain_right.n62 drain_right.n61 2.71565
R585 drain_right.n16 drain_right.n6 1.93989
R586 drain_right.n58 drain_right.n48 1.93989
R587 drain_right.n15 drain_right.n8 1.16414
R588 drain_right.n57 drain_right.n50 1.16414
R589 drain_right.n73 drain_right.n41 0.5005
R590 drain_right.n41 drain_right.n39 0.5005
R591 drain_right.n12 drain_right.n11 0.388379
R592 drain_right.n54 drain_right.n53 0.388379
R593 drain_right.n36 drain_right.n32 0.320154
R594 drain_right.n14 drain_right.n13 0.155672
R595 drain_right.n14 drain_right.n5 0.155672
R596 drain_right.n21 drain_right.n5 0.155672
R597 drain_right.n22 drain_right.n21 0.155672
R598 drain_right.n22 drain_right.n1 0.155672
R599 drain_right.n29 drain_right.n1 0.155672
R600 drain_right.n71 drain_right.n43 0.155672
R601 drain_right.n64 drain_right.n43 0.155672
R602 drain_right.n64 drain_right.n63 0.155672
R603 drain_right.n63 drain_right.n47 0.155672
R604 drain_right.n56 drain_right.n47 0.155672
R605 drain_right.n56 drain_right.n55 0.155672
R606 drain_right.n36 drain_right.n35 0.070154
C0 source plus 2.4938f
C1 drain_left drain_right 0.838543f
C2 source drain_right 16.5003f
C3 plus minus 4.09509f
C4 minus drain_right 2.54935f
C5 plus drain_right 0.31389f
C6 drain_left source 16.506401f
C7 drain_left minus 0.171605f
C8 source minus 2.47944f
C9 drain_left plus 2.70623f
C10 drain_right a_n1644_n2088# 5.50034f
C11 drain_left a_n1644_n2088# 5.77742f
C12 source a_n1644_n2088# 3.954995f
C13 minus a_n1644_n2088# 5.91924f
C14 plus a_n1644_n2088# 7.51596f
C15 drain_right.n0 a_n1644_n2088# 0.044834f
C16 drain_right.n1 a_n1644_n2088# 0.031897f
C17 drain_right.n2 a_n1644_n2088# 0.01714f
C18 drain_right.n3 a_n1644_n2088# 0.040513f
C19 drain_right.n4 a_n1644_n2088# 0.018148f
C20 drain_right.n5 a_n1644_n2088# 0.031897f
C21 drain_right.n6 a_n1644_n2088# 0.01714f
C22 drain_right.n7 a_n1644_n2088# 0.040513f
C23 drain_right.n8 a_n1644_n2088# 0.018148f
C24 drain_right.n9 a_n1644_n2088# 0.136497f
C25 drain_right.t5 a_n1644_n2088# 0.066031f
C26 drain_right.n10 a_n1644_n2088# 0.030385f
C27 drain_right.n11 a_n1644_n2088# 0.023931f
C28 drain_right.n12 a_n1644_n2088# 0.01714f
C29 drain_right.n13 a_n1644_n2088# 0.75896f
C30 drain_right.n14 a_n1644_n2088# 0.031897f
C31 drain_right.n15 a_n1644_n2088# 0.01714f
C32 drain_right.n16 a_n1644_n2088# 0.018148f
C33 drain_right.n17 a_n1644_n2088# 0.040513f
C34 drain_right.n18 a_n1644_n2088# 0.040513f
C35 drain_right.n19 a_n1644_n2088# 0.018148f
C36 drain_right.n20 a_n1644_n2088# 0.01714f
C37 drain_right.n21 a_n1644_n2088# 0.031897f
C38 drain_right.n22 a_n1644_n2088# 0.031897f
C39 drain_right.n23 a_n1644_n2088# 0.01714f
C40 drain_right.n24 a_n1644_n2088# 0.018148f
C41 drain_right.n25 a_n1644_n2088# 0.040513f
C42 drain_right.n26 a_n1644_n2088# 0.087704f
C43 drain_right.n27 a_n1644_n2088# 0.018148f
C44 drain_right.n28 a_n1644_n2088# 0.01714f
C45 drain_right.n29 a_n1644_n2088# 0.073729f
C46 drain_right.n30 a_n1644_n2088# 0.07224f
C47 drain_right.t3 a_n1644_n2088# 0.151236f
C48 drain_right.t8 a_n1644_n2088# 0.151236f
C49 drain_right.n31 a_n1644_n2088# 1.26131f
C50 drain_right.n32 a_n1644_n2088# 0.457112f
C51 drain_right.t7 a_n1644_n2088# 0.151236f
C52 drain_right.t9 a_n1644_n2088# 0.151236f
C53 drain_right.n33 a_n1644_n2088# 1.26408f
C54 drain_right.t11 a_n1644_n2088# 0.151236f
C55 drain_right.t0 a_n1644_n2088# 0.151236f
C56 drain_right.n34 a_n1644_n2088# 1.26131f
C57 drain_right.n35 a_n1644_n2088# 0.699802f
C58 drain_right.n36 a_n1644_n2088# 1.00632f
C59 drain_right.t12 a_n1644_n2088# 0.151236f
C60 drain_right.t4 a_n1644_n2088# 0.151236f
C61 drain_right.n37 a_n1644_n2088# 1.26408f
C62 drain_right.t13 a_n1644_n2088# 0.151236f
C63 drain_right.t6 a_n1644_n2088# 0.151236f
C64 drain_right.n38 a_n1644_n2088# 1.26132f
C65 drain_right.n39 a_n1644_n2088# 0.73341f
C66 drain_right.t10 a_n1644_n2088# 0.151236f
C67 drain_right.t2 a_n1644_n2088# 0.151236f
C68 drain_right.n40 a_n1644_n2088# 1.26132f
C69 drain_right.n41 a_n1644_n2088# 0.361662f
C70 drain_right.n42 a_n1644_n2088# 0.044834f
C71 drain_right.n43 a_n1644_n2088# 0.031897f
C72 drain_right.n44 a_n1644_n2088# 0.01714f
C73 drain_right.n45 a_n1644_n2088# 0.040513f
C74 drain_right.n46 a_n1644_n2088# 0.018148f
C75 drain_right.n47 a_n1644_n2088# 0.031897f
C76 drain_right.n48 a_n1644_n2088# 0.01714f
C77 drain_right.n49 a_n1644_n2088# 0.040513f
C78 drain_right.n50 a_n1644_n2088# 0.018148f
C79 drain_right.n51 a_n1644_n2088# 0.136497f
C80 drain_right.t1 a_n1644_n2088# 0.066031f
C81 drain_right.n52 a_n1644_n2088# 0.030385f
C82 drain_right.n53 a_n1644_n2088# 0.023931f
C83 drain_right.n54 a_n1644_n2088# 0.01714f
C84 drain_right.n55 a_n1644_n2088# 0.75896f
C85 drain_right.n56 a_n1644_n2088# 0.031897f
C86 drain_right.n57 a_n1644_n2088# 0.01714f
C87 drain_right.n58 a_n1644_n2088# 0.018148f
C88 drain_right.n59 a_n1644_n2088# 0.040513f
C89 drain_right.n60 a_n1644_n2088# 0.040513f
C90 drain_right.n61 a_n1644_n2088# 0.018148f
C91 drain_right.n62 a_n1644_n2088# 0.01714f
C92 drain_right.n63 a_n1644_n2088# 0.031897f
C93 drain_right.n64 a_n1644_n2088# 0.031897f
C94 drain_right.n65 a_n1644_n2088# 0.01714f
C95 drain_right.n66 a_n1644_n2088# 0.018148f
C96 drain_right.n67 a_n1644_n2088# 0.040513f
C97 drain_right.n68 a_n1644_n2088# 0.087704f
C98 drain_right.n69 a_n1644_n2088# 0.018148f
C99 drain_right.n70 a_n1644_n2088# 0.01714f
C100 drain_right.n71 a_n1644_n2088# 0.073729f
C101 drain_right.n72 a_n1644_n2088# 0.071098f
C102 drain_right.n73 a_n1644_n2088# 0.375491f
C103 minus.n0 a_n1644_n2088# 0.052568f
C104 minus.t12 a_n1644_n2088# 0.229668f
C105 minus.t3 a_n1644_n2088# 0.224662f
C106 minus.t11 a_n1644_n2088# 0.224662f
C107 minus.t0 a_n1644_n2088# 0.224662f
C108 minus.n1 a_n1644_n2088# 0.123263f
C109 minus.n2 a_n1644_n2088# 0.112519f
C110 minus.t7 a_n1644_n2088# 0.224662f
C111 minus.t1 a_n1644_n2088# 0.224662f
C112 minus.t9 a_n1644_n2088# 0.229668f
C113 minus.n3 a_n1644_n2088# 0.120596f
C114 minus.n4 a_n1644_n2088# 0.105824f
C115 minus.n5 a_n1644_n2088# 0.020031f
C116 minus.n6 a_n1644_n2088# 0.105824f
C117 minus.n7 a_n1644_n2088# 0.020031f
C118 minus.n8 a_n1644_n2088# 0.052568f
C119 minus.n9 a_n1644_n2088# 0.052568f
C120 minus.n10 a_n1644_n2088# 0.052568f
C121 minus.n11 a_n1644_n2088# 0.020031f
C122 minus.n12 a_n1644_n2088# 0.105824f
C123 minus.n13 a_n1644_n2088# 0.020031f
C124 minus.n14 a_n1644_n2088# 0.105824f
C125 minus.n15 a_n1644_n2088# 0.120526f
C126 minus.n16 a_n1644_n2088# 1.42404f
C127 minus.n17 a_n1644_n2088# 0.052568f
C128 minus.t6 a_n1644_n2088# 0.224662f
C129 minus.t13 a_n1644_n2088# 0.224662f
C130 minus.t2 a_n1644_n2088# 0.224662f
C131 minus.n18 a_n1644_n2088# 0.123263f
C132 minus.n19 a_n1644_n2088# 0.112519f
C133 minus.t5 a_n1644_n2088# 0.224662f
C134 minus.t10 a_n1644_n2088# 0.224662f
C135 minus.t8 a_n1644_n2088# 0.229668f
C136 minus.n20 a_n1644_n2088# 0.120596f
C137 minus.n21 a_n1644_n2088# 0.105824f
C138 minus.n22 a_n1644_n2088# 0.020031f
C139 minus.n23 a_n1644_n2088# 0.105824f
C140 minus.n24 a_n1644_n2088# 0.020031f
C141 minus.n25 a_n1644_n2088# 0.052568f
C142 minus.n26 a_n1644_n2088# 0.052568f
C143 minus.n27 a_n1644_n2088# 0.052568f
C144 minus.n28 a_n1644_n2088# 0.020031f
C145 minus.n29 a_n1644_n2088# 0.105824f
C146 minus.n30 a_n1644_n2088# 0.020031f
C147 minus.n31 a_n1644_n2088# 0.105824f
C148 minus.t4 a_n1644_n2088# 0.229668f
C149 minus.n32 a_n1644_n2088# 0.120526f
C150 minus.n33 a_n1644_n2088# 0.337624f
C151 minus.n34 a_n1644_n2088# 1.75733f
C152 source.n0 a_n1644_n2088# 0.048676f
C153 source.n1 a_n1644_n2088# 0.034631f
C154 source.n2 a_n1644_n2088# 0.018609f
C155 source.n3 a_n1644_n2088# 0.043985f
C156 source.n4 a_n1644_n2088# 0.019704f
C157 source.n5 a_n1644_n2088# 0.034631f
C158 source.n6 a_n1644_n2088# 0.018609f
C159 source.n7 a_n1644_n2088# 0.043985f
C160 source.n8 a_n1644_n2088# 0.019704f
C161 source.n9 a_n1644_n2088# 0.148195f
C162 source.t20 a_n1644_n2088# 0.07169f
C163 source.n10 a_n1644_n2088# 0.032989f
C164 source.n11 a_n1644_n2088# 0.025982f
C165 source.n12 a_n1644_n2088# 0.018609f
C166 source.n13 a_n1644_n2088# 0.824002f
C167 source.n14 a_n1644_n2088# 0.034631f
C168 source.n15 a_n1644_n2088# 0.018609f
C169 source.n16 a_n1644_n2088# 0.019704f
C170 source.n17 a_n1644_n2088# 0.043985f
C171 source.n18 a_n1644_n2088# 0.043985f
C172 source.n19 a_n1644_n2088# 0.019704f
C173 source.n20 a_n1644_n2088# 0.018609f
C174 source.n21 a_n1644_n2088# 0.034631f
C175 source.n22 a_n1644_n2088# 0.034631f
C176 source.n23 a_n1644_n2088# 0.018609f
C177 source.n24 a_n1644_n2088# 0.019704f
C178 source.n25 a_n1644_n2088# 0.043985f
C179 source.n26 a_n1644_n2088# 0.09522f
C180 source.n27 a_n1644_n2088# 0.019704f
C181 source.n28 a_n1644_n2088# 0.018609f
C182 source.n29 a_n1644_n2088# 0.080047f
C183 source.n30 a_n1644_n2088# 0.053279f
C184 source.n31 a_n1644_n2088# 0.830574f
C185 source.t19 a_n1644_n2088# 0.164197f
C186 source.t14 a_n1644_n2088# 0.164197f
C187 source.n32 a_n1644_n2088# 1.27878f
C188 source.n33 a_n1644_n2088# 0.436216f
C189 source.t18 a_n1644_n2088# 0.164197f
C190 source.t27 a_n1644_n2088# 0.164197f
C191 source.n34 a_n1644_n2088# 1.27878f
C192 source.n35 a_n1644_n2088# 0.436216f
C193 source.t24 a_n1644_n2088# 0.164197f
C194 source.t26 a_n1644_n2088# 0.164197f
C195 source.n36 a_n1644_n2088# 1.27878f
C196 source.n37 a_n1644_n2088# 0.460746f
C197 source.n38 a_n1644_n2088# 0.048676f
C198 source.n39 a_n1644_n2088# 0.034631f
C199 source.n40 a_n1644_n2088# 0.018609f
C200 source.n41 a_n1644_n2088# 0.043985f
C201 source.n42 a_n1644_n2088# 0.019704f
C202 source.n43 a_n1644_n2088# 0.034631f
C203 source.n44 a_n1644_n2088# 0.018609f
C204 source.n45 a_n1644_n2088# 0.043985f
C205 source.n46 a_n1644_n2088# 0.019704f
C206 source.n47 a_n1644_n2088# 0.148195f
C207 source.t11 a_n1644_n2088# 0.07169f
C208 source.n48 a_n1644_n2088# 0.032989f
C209 source.n49 a_n1644_n2088# 0.025982f
C210 source.n50 a_n1644_n2088# 0.018609f
C211 source.n51 a_n1644_n2088# 0.824002f
C212 source.n52 a_n1644_n2088# 0.034631f
C213 source.n53 a_n1644_n2088# 0.018609f
C214 source.n54 a_n1644_n2088# 0.019704f
C215 source.n55 a_n1644_n2088# 0.043985f
C216 source.n56 a_n1644_n2088# 0.043985f
C217 source.n57 a_n1644_n2088# 0.019704f
C218 source.n58 a_n1644_n2088# 0.018609f
C219 source.n59 a_n1644_n2088# 0.034631f
C220 source.n60 a_n1644_n2088# 0.034631f
C221 source.n61 a_n1644_n2088# 0.018609f
C222 source.n62 a_n1644_n2088# 0.019704f
C223 source.n63 a_n1644_n2088# 0.043985f
C224 source.n64 a_n1644_n2088# 0.09522f
C225 source.n65 a_n1644_n2088# 0.019704f
C226 source.n66 a_n1644_n2088# 0.018609f
C227 source.n67 a_n1644_n2088# 0.080047f
C228 source.n68 a_n1644_n2088# 0.053279f
C229 source.n69 a_n1644_n2088# 0.165695f
C230 source.t4 a_n1644_n2088# 0.164197f
C231 source.t10 a_n1644_n2088# 0.164197f
C232 source.n70 a_n1644_n2088# 1.27878f
C233 source.n71 a_n1644_n2088# 0.436216f
C234 source.t12 a_n1644_n2088# 0.164197f
C235 source.t7 a_n1644_n2088# 0.164197f
C236 source.n72 a_n1644_n2088# 1.27878f
C237 source.n73 a_n1644_n2088# 0.436216f
C238 source.t2 a_n1644_n2088# 0.164197f
C239 source.t6 a_n1644_n2088# 0.164197f
C240 source.n74 a_n1644_n2088# 1.27878f
C241 source.n75 a_n1644_n2088# 1.62588f
C242 source.t23 a_n1644_n2088# 0.164197f
C243 source.t21 a_n1644_n2088# 0.164197f
C244 source.n76 a_n1644_n2088# 1.27877f
C245 source.n77 a_n1644_n2088# 1.62589f
C246 source.t15 a_n1644_n2088# 0.164197f
C247 source.t16 a_n1644_n2088# 0.164197f
C248 source.n78 a_n1644_n2088# 1.27877f
C249 source.n79 a_n1644_n2088# 0.436225f
C250 source.t25 a_n1644_n2088# 0.164197f
C251 source.t22 a_n1644_n2088# 0.164197f
C252 source.n80 a_n1644_n2088# 1.27877f
C253 source.n81 a_n1644_n2088# 0.436225f
C254 source.n82 a_n1644_n2088# 0.048676f
C255 source.n83 a_n1644_n2088# 0.034631f
C256 source.n84 a_n1644_n2088# 0.018609f
C257 source.n85 a_n1644_n2088# 0.043985f
C258 source.n86 a_n1644_n2088# 0.019704f
C259 source.n87 a_n1644_n2088# 0.034631f
C260 source.n88 a_n1644_n2088# 0.018609f
C261 source.n89 a_n1644_n2088# 0.043985f
C262 source.n90 a_n1644_n2088# 0.019704f
C263 source.n91 a_n1644_n2088# 0.148195f
C264 source.t17 a_n1644_n2088# 0.07169f
C265 source.n92 a_n1644_n2088# 0.032989f
C266 source.n93 a_n1644_n2088# 0.025982f
C267 source.n94 a_n1644_n2088# 0.018609f
C268 source.n95 a_n1644_n2088# 0.824002f
C269 source.n96 a_n1644_n2088# 0.034631f
C270 source.n97 a_n1644_n2088# 0.018609f
C271 source.n98 a_n1644_n2088# 0.019704f
C272 source.n99 a_n1644_n2088# 0.043985f
C273 source.n100 a_n1644_n2088# 0.043985f
C274 source.n101 a_n1644_n2088# 0.019704f
C275 source.n102 a_n1644_n2088# 0.018609f
C276 source.n103 a_n1644_n2088# 0.034631f
C277 source.n104 a_n1644_n2088# 0.034631f
C278 source.n105 a_n1644_n2088# 0.018609f
C279 source.n106 a_n1644_n2088# 0.019704f
C280 source.n107 a_n1644_n2088# 0.043985f
C281 source.n108 a_n1644_n2088# 0.09522f
C282 source.n109 a_n1644_n2088# 0.019704f
C283 source.n110 a_n1644_n2088# 0.018609f
C284 source.n111 a_n1644_n2088# 0.080047f
C285 source.n112 a_n1644_n2088# 0.053279f
C286 source.n113 a_n1644_n2088# 0.165695f
C287 source.t9 a_n1644_n2088# 0.164197f
C288 source.t0 a_n1644_n2088# 0.164197f
C289 source.n114 a_n1644_n2088# 1.27877f
C290 source.n115 a_n1644_n2088# 0.460755f
C291 source.t8 a_n1644_n2088# 0.164197f
C292 source.t5 a_n1644_n2088# 0.164197f
C293 source.n116 a_n1644_n2088# 1.27877f
C294 source.n117 a_n1644_n2088# 0.436225f
C295 source.t1 a_n1644_n2088# 0.164197f
C296 source.t3 a_n1644_n2088# 0.164197f
C297 source.n118 a_n1644_n2088# 1.27877f
C298 source.n119 a_n1644_n2088# 0.436225f
C299 source.n120 a_n1644_n2088# 0.048676f
C300 source.n121 a_n1644_n2088# 0.034631f
C301 source.n122 a_n1644_n2088# 0.018609f
C302 source.n123 a_n1644_n2088# 0.043985f
C303 source.n124 a_n1644_n2088# 0.019704f
C304 source.n125 a_n1644_n2088# 0.034631f
C305 source.n126 a_n1644_n2088# 0.018609f
C306 source.n127 a_n1644_n2088# 0.043985f
C307 source.n128 a_n1644_n2088# 0.019704f
C308 source.n129 a_n1644_n2088# 0.148195f
C309 source.t13 a_n1644_n2088# 0.07169f
C310 source.n130 a_n1644_n2088# 0.032989f
C311 source.n131 a_n1644_n2088# 0.025982f
C312 source.n132 a_n1644_n2088# 0.018609f
C313 source.n133 a_n1644_n2088# 0.824002f
C314 source.n134 a_n1644_n2088# 0.034631f
C315 source.n135 a_n1644_n2088# 0.018609f
C316 source.n136 a_n1644_n2088# 0.019704f
C317 source.n137 a_n1644_n2088# 0.043985f
C318 source.n138 a_n1644_n2088# 0.043985f
C319 source.n139 a_n1644_n2088# 0.019704f
C320 source.n140 a_n1644_n2088# 0.018609f
C321 source.n141 a_n1644_n2088# 0.034631f
C322 source.n142 a_n1644_n2088# 0.034631f
C323 source.n143 a_n1644_n2088# 0.018609f
C324 source.n144 a_n1644_n2088# 0.019704f
C325 source.n145 a_n1644_n2088# 0.043985f
C326 source.n146 a_n1644_n2088# 0.09522f
C327 source.n147 a_n1644_n2088# 0.019704f
C328 source.n148 a_n1644_n2088# 0.018609f
C329 source.n149 a_n1644_n2088# 0.080047f
C330 source.n150 a_n1644_n2088# 0.053279f
C331 source.n151 a_n1644_n2088# 0.329437f
C332 source.n152 a_n1644_n2088# 1.41469f
C333 drain_left.n0 a_n1644_n2088# 0.04501f
C334 drain_left.n1 a_n1644_n2088# 0.032023f
C335 drain_left.n2 a_n1644_n2088# 0.017208f
C336 drain_left.n3 a_n1644_n2088# 0.040672f
C337 drain_left.n4 a_n1644_n2088# 0.01822f
C338 drain_left.n5 a_n1644_n2088# 0.032023f
C339 drain_left.n6 a_n1644_n2088# 0.017208f
C340 drain_left.n7 a_n1644_n2088# 0.040672f
C341 drain_left.n8 a_n1644_n2088# 0.01822f
C342 drain_left.n9 a_n1644_n2088# 0.137034f
C343 drain_left.t8 a_n1644_n2088# 0.066291f
C344 drain_left.n10 a_n1644_n2088# 0.030504f
C345 drain_left.n11 a_n1644_n2088# 0.024025f
C346 drain_left.n12 a_n1644_n2088# 0.017208f
C347 drain_left.n13 a_n1644_n2088# 0.761945f
C348 drain_left.n14 a_n1644_n2088# 0.032023f
C349 drain_left.n15 a_n1644_n2088# 0.017208f
C350 drain_left.n16 a_n1644_n2088# 0.01822f
C351 drain_left.n17 a_n1644_n2088# 0.040672f
C352 drain_left.n18 a_n1644_n2088# 0.040672f
C353 drain_left.n19 a_n1644_n2088# 0.01822f
C354 drain_left.n20 a_n1644_n2088# 0.017208f
C355 drain_left.n21 a_n1644_n2088# 0.032023f
C356 drain_left.n22 a_n1644_n2088# 0.032023f
C357 drain_left.n23 a_n1644_n2088# 0.017208f
C358 drain_left.n24 a_n1644_n2088# 0.01822f
C359 drain_left.n25 a_n1644_n2088# 0.040672f
C360 drain_left.n26 a_n1644_n2088# 0.088049f
C361 drain_left.n27 a_n1644_n2088# 0.01822f
C362 drain_left.n28 a_n1644_n2088# 0.017208f
C363 drain_left.n29 a_n1644_n2088# 0.074019f
C364 drain_left.n30 a_n1644_n2088# 0.072525f
C365 drain_left.t10 a_n1644_n2088# 0.151831f
C366 drain_left.t4 a_n1644_n2088# 0.151831f
C367 drain_left.n31 a_n1644_n2088# 1.26627f
C368 drain_left.n32 a_n1644_n2088# 0.45891f
C369 drain_left.t9 a_n1644_n2088# 0.151831f
C370 drain_left.t6 a_n1644_n2088# 0.151831f
C371 drain_left.n33 a_n1644_n2088# 1.26905f
C372 drain_left.t11 a_n1644_n2088# 0.151831f
C373 drain_left.t13 a_n1644_n2088# 0.151831f
C374 drain_left.n34 a_n1644_n2088# 1.26627f
C375 drain_left.n35 a_n1644_n2088# 0.702554f
C376 drain_left.n36 a_n1644_n2088# 1.07549f
C377 drain_left.n37 a_n1644_n2088# 0.04501f
C378 drain_left.n38 a_n1644_n2088# 0.032023f
C379 drain_left.n39 a_n1644_n2088# 0.017208f
C380 drain_left.n40 a_n1644_n2088# 0.040672f
C381 drain_left.n41 a_n1644_n2088# 0.01822f
C382 drain_left.n42 a_n1644_n2088# 0.032023f
C383 drain_left.n43 a_n1644_n2088# 0.017208f
C384 drain_left.n44 a_n1644_n2088# 0.040672f
C385 drain_left.n45 a_n1644_n2088# 0.01822f
C386 drain_left.n46 a_n1644_n2088# 0.137034f
C387 drain_left.t7 a_n1644_n2088# 0.066291f
C388 drain_left.n47 a_n1644_n2088# 0.030504f
C389 drain_left.n48 a_n1644_n2088# 0.024025f
C390 drain_left.n49 a_n1644_n2088# 0.017208f
C391 drain_left.n50 a_n1644_n2088# 0.761945f
C392 drain_left.n51 a_n1644_n2088# 0.032023f
C393 drain_left.n52 a_n1644_n2088# 0.017208f
C394 drain_left.n53 a_n1644_n2088# 0.01822f
C395 drain_left.n54 a_n1644_n2088# 0.040672f
C396 drain_left.n55 a_n1644_n2088# 0.040672f
C397 drain_left.n56 a_n1644_n2088# 0.01822f
C398 drain_left.n57 a_n1644_n2088# 0.017208f
C399 drain_left.n58 a_n1644_n2088# 0.032023f
C400 drain_left.n59 a_n1644_n2088# 0.032023f
C401 drain_left.n60 a_n1644_n2088# 0.017208f
C402 drain_left.n61 a_n1644_n2088# 0.01822f
C403 drain_left.n62 a_n1644_n2088# 0.040672f
C404 drain_left.n63 a_n1644_n2088# 0.088049f
C405 drain_left.n64 a_n1644_n2088# 0.01822f
C406 drain_left.n65 a_n1644_n2088# 0.017208f
C407 drain_left.n66 a_n1644_n2088# 0.074019f
C408 drain_left.n67 a_n1644_n2088# 0.072525f
C409 drain_left.t2 a_n1644_n2088# 0.151831f
C410 drain_left.t1 a_n1644_n2088# 0.151831f
C411 drain_left.n68 a_n1644_n2088# 1.26628f
C412 drain_left.n69 a_n1644_n2088# 0.47519f
C413 drain_left.t12 a_n1644_n2088# 0.151831f
C414 drain_left.t3 a_n1644_n2088# 0.151831f
C415 drain_left.n70 a_n1644_n2088# 1.26628f
C416 drain_left.n71 a_n1644_n2088# 0.363084f
C417 drain_left.t5 a_n1644_n2088# 0.151831f
C418 drain_left.t0 a_n1644_n2088# 0.151831f
C419 drain_left.n72 a_n1644_n2088# 1.26627f
C420 drain_left.n73 a_n1644_n2088# 0.627414f
C421 plus.n0 a_n1644_n2088# 0.054358f
C422 plus.t13 a_n1644_n2088# 0.232314f
C423 plus.t8 a_n1644_n2088# 0.232314f
C424 plus.t0 a_n1644_n2088# 0.232314f
C425 plus.n1 a_n1644_n2088# 0.127461f
C426 plus.n2 a_n1644_n2088# 0.116352f
C427 plus.t9 a_n1644_n2088# 0.232314f
C428 plus.t1 a_n1644_n2088# 0.232314f
C429 plus.t3 a_n1644_n2088# 0.23749f
C430 plus.n3 a_n1644_n2088# 0.124703f
C431 plus.n4 a_n1644_n2088# 0.109429f
C432 plus.n5 a_n1644_n2088# 0.020713f
C433 plus.n6 a_n1644_n2088# 0.109429f
C434 plus.n7 a_n1644_n2088# 0.020713f
C435 plus.n8 a_n1644_n2088# 0.054358f
C436 plus.n9 a_n1644_n2088# 0.054358f
C437 plus.n10 a_n1644_n2088# 0.054358f
C438 plus.n11 a_n1644_n2088# 0.020713f
C439 plus.n12 a_n1644_n2088# 0.109429f
C440 plus.n13 a_n1644_n2088# 0.020713f
C441 plus.n14 a_n1644_n2088# 0.109429f
C442 plus.t7 a_n1644_n2088# 0.23749f
C443 plus.n15 a_n1644_n2088# 0.124631f
C444 plus.n16 a_n1644_n2088# 0.45927f
C445 plus.n17 a_n1644_n2088# 0.054358f
C446 plus.t4 a_n1644_n2088# 0.23749f
C447 plus.t6 a_n1644_n2088# 0.232314f
C448 plus.t12 a_n1644_n2088# 0.232314f
C449 plus.t11 a_n1644_n2088# 0.232314f
C450 plus.n18 a_n1644_n2088# 0.127461f
C451 plus.n19 a_n1644_n2088# 0.116352f
C452 plus.t2 a_n1644_n2088# 0.232314f
C453 plus.t5 a_n1644_n2088# 0.232314f
C454 plus.t10 a_n1644_n2088# 0.23749f
C455 plus.n20 a_n1644_n2088# 0.124703f
C456 plus.n21 a_n1644_n2088# 0.109429f
C457 plus.n22 a_n1644_n2088# 0.020713f
C458 plus.n23 a_n1644_n2088# 0.109429f
C459 plus.n24 a_n1644_n2088# 0.020713f
C460 plus.n25 a_n1644_n2088# 0.054358f
C461 plus.n26 a_n1644_n2088# 0.054358f
C462 plus.n27 a_n1644_n2088# 0.054358f
C463 plus.n28 a_n1644_n2088# 0.020713f
C464 plus.n29 a_n1644_n2088# 0.109429f
C465 plus.n30 a_n1644_n2088# 0.020713f
C466 plus.n31 a_n1644_n2088# 0.109429f
C467 plus.n32 a_n1644_n2088# 0.124631f
C468 plus.n33 a_n1644_n2088# 1.32989f
.ends

