* NGSPICE file created from diffpair368.ext - technology: sky130A

.subckt diffpair368 minus drain_right drain_left source plus
X0 drain_right.t19 minus.t0 source.t24 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X1 source.t37 minus.t1 drain_right.t18 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X2 drain_left.t19 plus.t0 source.t9 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 drain_left.t18 plus.t1 source.t13 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 source.t35 minus.t2 drain_right.t17 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X5 source.t7 plus.t2 drain_left.t17 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X6 drain_right.t16 minus.t3 source.t33 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X7 source.t8 plus.t3 drain_left.t16 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X8 source.t23 minus.t4 drain_right.t15 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X9 drain_left.t15 plus.t4 source.t19 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X10 source.t10 plus.t5 drain_left.t14 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X11 drain_right.t14 minus.t5 source.t26 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X12 source.t3 plus.t6 drain_left.t13 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X13 drain_right.t13 minus.t6 source.t38 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X14 drain_right.t12 minus.t7 source.t29 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X15 source.t31 minus.t8 drain_right.t11 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X16 a_n2542_n2688# a_n2542_n2688# a_n2542_n2688# a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.5
X17 drain_left.t12 plus.t7 source.t5 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X18 a_n2542_n2688# a_n2542_n2688# a_n2542_n2688# a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X19 source.t21 minus.t9 drain_right.t10 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X20 drain_right.t9 minus.t10 source.t32 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X21 source.t11 plus.t8 drain_left.t11 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X22 source.t25 minus.t11 drain_right.t8 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X23 source.t36 minus.t12 drain_right.t7 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X24 drain_right.t6 minus.t13 source.t27 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X25 drain_left.t10 plus.t9 source.t14 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X26 drain_right.t5 minus.t14 source.t22 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X27 drain_left.t9 plus.t10 source.t0 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X28 drain_right.t4 minus.t15 source.t20 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X29 drain_left.t8 plus.t11 source.t16 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X30 source.t2 plus.t12 drain_left.t7 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X31 source.t28 minus.t16 drain_right.t3 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X32 a_n2542_n2688# a_n2542_n2688# a_n2542_n2688# a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X33 source.t1 plus.t13 drain_left.t6 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X34 source.t39 minus.t17 drain_right.t2 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X35 source.t18 plus.t14 drain_left.t5 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X36 source.t4 plus.t15 drain_left.t4 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X37 drain_left.t3 plus.t16 source.t17 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X38 drain_left.t2 plus.t17 source.t6 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X39 source.t12 plus.t18 drain_left.t1 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X40 a_n2542_n2688# a_n2542_n2688# a_n2542_n2688# a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X41 drain_right.t1 minus.t18 source.t34 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X42 source.t30 minus.t19 drain_right.t0 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X43 drain_left.t0 plus.t19 source.t15 a_n2542_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 minus.n6 minus.t14 533.348
R1 minus.n34 minus.t19 533.348
R2 minus.n7 minus.t2 512.366
R3 minus.n5 minus.t7 512.366
R4 minus.n13 minus.t16 512.366
R5 minus.n14 minus.t5 512.366
R6 minus.n18 minus.t11 512.366
R7 minus.n19 minus.t0 512.366
R8 minus.n1 minus.t12 512.366
R9 minus.n25 minus.t15 512.366
R10 minus.n26 minus.t4 512.366
R11 minus.n35 minus.t18 512.366
R12 minus.n33 minus.t8 512.366
R13 minus.n41 minus.t6 512.366
R14 minus.n42 minus.t1 512.366
R15 minus.n46 minus.t10 512.366
R16 minus.n47 minus.t9 512.366
R17 minus.n29 minus.t3 512.366
R18 minus.n53 minus.t17 512.366
R19 minus.n54 minus.t13 512.366
R20 minus.n27 minus.n26 161.3
R21 minus.n25 minus.n0 161.3
R22 minus.n24 minus.n23 161.3
R23 minus.n22 minus.n1 161.3
R24 minus.n21 minus.n20 161.3
R25 minus.n19 minus.n2 161.3
R26 minus.n18 minus.n17 161.3
R27 minus.n16 minus.n3 161.3
R28 minus.n15 minus.n14 161.3
R29 minus.n13 minus.n4 161.3
R30 minus.n12 minus.n11 161.3
R31 minus.n10 minus.n5 161.3
R32 minus.n9 minus.n8 161.3
R33 minus.n55 minus.n54 161.3
R34 minus.n53 minus.n28 161.3
R35 minus.n52 minus.n51 161.3
R36 minus.n50 minus.n29 161.3
R37 minus.n49 minus.n48 161.3
R38 minus.n47 minus.n30 161.3
R39 minus.n46 minus.n45 161.3
R40 minus.n44 minus.n31 161.3
R41 minus.n43 minus.n42 161.3
R42 minus.n41 minus.n32 161.3
R43 minus.n40 minus.n39 161.3
R44 minus.n38 minus.n33 161.3
R45 minus.n37 minus.n36 161.3
R46 minus.n9 minus.n6 70.4033
R47 minus.n37 minus.n34 70.4033
R48 minus.n14 minus.n13 48.2005
R49 minus.n19 minus.n18 48.2005
R50 minus.n26 minus.n25 48.2005
R51 minus.n42 minus.n41 48.2005
R52 minus.n47 minus.n46 48.2005
R53 minus.n54 minus.n53 48.2005
R54 minus.n12 minus.n5 47.4702
R55 minus.n20 minus.n1 47.4702
R56 minus.n40 minus.n33 47.4702
R57 minus.n48 minus.n29 47.4702
R58 minus.n56 minus.n27 36.5687
R59 minus.n8 minus.n5 25.5611
R60 minus.n24 minus.n1 25.5611
R61 minus.n36 minus.n33 25.5611
R62 minus.n52 minus.n29 25.5611
R63 minus.n18 minus.n3 24.1005
R64 minus.n14 minus.n3 24.1005
R65 minus.n42 minus.n31 24.1005
R66 minus.n46 minus.n31 24.1005
R67 minus.n8 minus.n7 22.6399
R68 minus.n25 minus.n24 22.6399
R69 minus.n36 minus.n35 22.6399
R70 minus.n53 minus.n52 22.6399
R71 minus.n7 minus.n6 20.9576
R72 minus.n35 minus.n34 20.9576
R73 minus.n56 minus.n55 6.59141
R74 minus.n13 minus.n12 0.730803
R75 minus.n20 minus.n19 0.730803
R76 minus.n41 minus.n40 0.730803
R77 minus.n48 minus.n47 0.730803
R78 minus.n27 minus.n0 0.189894
R79 minus.n23 minus.n0 0.189894
R80 minus.n23 minus.n22 0.189894
R81 minus.n22 minus.n21 0.189894
R82 minus.n21 minus.n2 0.189894
R83 minus.n17 minus.n2 0.189894
R84 minus.n17 minus.n16 0.189894
R85 minus.n16 minus.n15 0.189894
R86 minus.n15 minus.n4 0.189894
R87 minus.n11 minus.n4 0.189894
R88 minus.n11 minus.n10 0.189894
R89 minus.n10 minus.n9 0.189894
R90 minus.n38 minus.n37 0.189894
R91 minus.n39 minus.n38 0.189894
R92 minus.n39 minus.n32 0.189894
R93 minus.n43 minus.n32 0.189894
R94 minus.n44 minus.n43 0.189894
R95 minus.n45 minus.n44 0.189894
R96 minus.n45 minus.n30 0.189894
R97 minus.n49 minus.n30 0.189894
R98 minus.n50 minus.n49 0.189894
R99 minus.n51 minus.n50 0.189894
R100 minus.n51 minus.n28 0.189894
R101 minus.n55 minus.n28 0.189894
R102 minus minus.n56 0.188
R103 source.n9 source.t8 51.0588
R104 source.n10 source.t22 51.0588
R105 source.n19 source.t23 51.0588
R106 source.n39 source.t27 51.0586
R107 source.n30 source.t30 51.0586
R108 source.n29 source.t16 51.0586
R109 source.n20 source.t10 51.0586
R110 source.n0 source.t14 51.0586
R111 source.n2 source.n1 48.8588
R112 source.n4 source.n3 48.8588
R113 source.n6 source.n5 48.8588
R114 source.n8 source.n7 48.8588
R115 source.n12 source.n11 48.8588
R116 source.n14 source.n13 48.8588
R117 source.n16 source.n15 48.8588
R118 source.n18 source.n17 48.8588
R119 source.n38 source.n37 48.8586
R120 source.n36 source.n35 48.8586
R121 source.n34 source.n33 48.8586
R122 source.n32 source.n31 48.8586
R123 source.n28 source.n27 48.8586
R124 source.n26 source.n25 48.8586
R125 source.n24 source.n23 48.8586
R126 source.n22 source.n21 48.8586
R127 source.n20 source.n19 19.7305
R128 source.n40 source.n0 14.1098
R129 source.n40 source.n39 5.62119
R130 source.n37 source.t33 2.2005
R131 source.n37 source.t39 2.2005
R132 source.n35 source.t32 2.2005
R133 source.n35 source.t21 2.2005
R134 source.n33 source.t38 2.2005
R135 source.n33 source.t37 2.2005
R136 source.n31 source.t34 2.2005
R137 source.n31 source.t31 2.2005
R138 source.n27 source.t13 2.2005
R139 source.n27 source.t2 2.2005
R140 source.n25 source.t17 2.2005
R141 source.n25 source.t4 2.2005
R142 source.n23 source.t9 2.2005
R143 source.n23 source.t3 2.2005
R144 source.n21 source.t19 2.2005
R145 source.n21 source.t1 2.2005
R146 source.n1 source.t6 2.2005
R147 source.n1 source.t7 2.2005
R148 source.n3 source.t15 2.2005
R149 source.n3 source.t11 2.2005
R150 source.n5 source.t5 2.2005
R151 source.n5 source.t18 2.2005
R152 source.n7 source.t0 2.2005
R153 source.n7 source.t12 2.2005
R154 source.n11 source.t29 2.2005
R155 source.n11 source.t35 2.2005
R156 source.n13 source.t26 2.2005
R157 source.n13 source.t28 2.2005
R158 source.n15 source.t24 2.2005
R159 source.n15 source.t25 2.2005
R160 source.n17 source.t20 2.2005
R161 source.n17 source.t36 2.2005
R162 source.n19 source.n18 0.716017
R163 source.n18 source.n16 0.716017
R164 source.n16 source.n14 0.716017
R165 source.n14 source.n12 0.716017
R166 source.n12 source.n10 0.716017
R167 source.n9 source.n8 0.716017
R168 source.n8 source.n6 0.716017
R169 source.n6 source.n4 0.716017
R170 source.n4 source.n2 0.716017
R171 source.n2 source.n0 0.716017
R172 source.n22 source.n20 0.716017
R173 source.n24 source.n22 0.716017
R174 source.n26 source.n24 0.716017
R175 source.n28 source.n26 0.716017
R176 source.n29 source.n28 0.716017
R177 source.n32 source.n30 0.716017
R178 source.n34 source.n32 0.716017
R179 source.n36 source.n34 0.716017
R180 source.n38 source.n36 0.716017
R181 source.n39 source.n38 0.716017
R182 source.n10 source.n9 0.470328
R183 source.n30 source.n29 0.470328
R184 source source.n40 0.188
R185 drain_right.n10 drain_right.n8 66.2529
R186 drain_right.n6 drain_right.n4 66.2529
R187 drain_right.n2 drain_right.n0 66.2529
R188 drain_right.n10 drain_right.n9 65.5376
R189 drain_right.n12 drain_right.n11 65.5376
R190 drain_right.n14 drain_right.n13 65.5376
R191 drain_right.n16 drain_right.n15 65.5376
R192 drain_right.n7 drain_right.n3 65.5373
R193 drain_right.n6 drain_right.n5 65.5373
R194 drain_right.n2 drain_right.n1 65.5373
R195 drain_right drain_right.n7 30.2653
R196 drain_right drain_right.n16 6.36873
R197 drain_right.n3 drain_right.t18 2.2005
R198 drain_right.n3 drain_right.t9 2.2005
R199 drain_right.n4 drain_right.t2 2.2005
R200 drain_right.n4 drain_right.t6 2.2005
R201 drain_right.n5 drain_right.t10 2.2005
R202 drain_right.n5 drain_right.t16 2.2005
R203 drain_right.n1 drain_right.t11 2.2005
R204 drain_right.n1 drain_right.t13 2.2005
R205 drain_right.n0 drain_right.t0 2.2005
R206 drain_right.n0 drain_right.t1 2.2005
R207 drain_right.n8 drain_right.t17 2.2005
R208 drain_right.n8 drain_right.t5 2.2005
R209 drain_right.n9 drain_right.t3 2.2005
R210 drain_right.n9 drain_right.t12 2.2005
R211 drain_right.n11 drain_right.t8 2.2005
R212 drain_right.n11 drain_right.t14 2.2005
R213 drain_right.n13 drain_right.t7 2.2005
R214 drain_right.n13 drain_right.t19 2.2005
R215 drain_right.n15 drain_right.t15 2.2005
R216 drain_right.n15 drain_right.t4 2.2005
R217 drain_right.n16 drain_right.n14 0.716017
R218 drain_right.n14 drain_right.n12 0.716017
R219 drain_right.n12 drain_right.n10 0.716017
R220 drain_right.n7 drain_right.n6 0.660671
R221 drain_right.n7 drain_right.n2 0.660671
R222 plus.n8 plus.t3 533.348
R223 plus.n36 plus.t11 533.348
R224 plus.n26 plus.t9 512.366
R225 plus.n25 plus.t2 512.366
R226 plus.n1 plus.t17 512.366
R227 plus.n19 plus.t8 512.366
R228 plus.n18 plus.t19 512.366
R229 plus.n4 plus.t14 512.366
R230 plus.n13 plus.t7 512.366
R231 plus.n11 plus.t18 512.366
R232 plus.n7 plus.t10 512.366
R233 plus.n54 plus.t5 512.366
R234 plus.n53 plus.t4 512.366
R235 plus.n29 plus.t13 512.366
R236 plus.n47 plus.t0 512.366
R237 plus.n46 plus.t6 512.366
R238 plus.n32 plus.t16 512.366
R239 plus.n41 plus.t15 512.366
R240 plus.n39 plus.t1 512.366
R241 plus.n35 plus.t12 512.366
R242 plus.n10 plus.n9 161.3
R243 plus.n11 plus.n6 161.3
R244 plus.n12 plus.n5 161.3
R245 plus.n14 plus.n13 161.3
R246 plus.n15 plus.n4 161.3
R247 plus.n17 plus.n16 161.3
R248 plus.n18 plus.n3 161.3
R249 plus.n19 plus.n2 161.3
R250 plus.n21 plus.n20 161.3
R251 plus.n22 plus.n1 161.3
R252 plus.n24 plus.n23 161.3
R253 plus.n25 plus.n0 161.3
R254 plus.n27 plus.n26 161.3
R255 plus.n38 plus.n37 161.3
R256 plus.n39 plus.n34 161.3
R257 plus.n40 plus.n33 161.3
R258 plus.n42 plus.n41 161.3
R259 plus.n43 plus.n32 161.3
R260 plus.n45 plus.n44 161.3
R261 plus.n46 plus.n31 161.3
R262 plus.n47 plus.n30 161.3
R263 plus.n49 plus.n48 161.3
R264 plus.n50 plus.n29 161.3
R265 plus.n52 plus.n51 161.3
R266 plus.n53 plus.n28 161.3
R267 plus.n55 plus.n54 161.3
R268 plus.n9 plus.n8 70.4033
R269 plus.n37 plus.n36 70.4033
R270 plus.n26 plus.n25 48.2005
R271 plus.n19 plus.n18 48.2005
R272 plus.n13 plus.n4 48.2005
R273 plus.n54 plus.n53 48.2005
R274 plus.n47 plus.n46 48.2005
R275 plus.n41 plus.n32 48.2005
R276 plus.n20 plus.n1 47.4702
R277 plus.n12 plus.n11 47.4702
R278 plus.n48 plus.n29 47.4702
R279 plus.n40 plus.n39 47.4702
R280 plus plus.n55 31.5861
R281 plus.n24 plus.n1 25.5611
R282 plus.n11 plus.n10 25.5611
R283 plus.n52 plus.n29 25.5611
R284 plus.n39 plus.n38 25.5611
R285 plus.n17 plus.n4 24.1005
R286 plus.n18 plus.n17 24.1005
R287 plus.n46 plus.n45 24.1005
R288 plus.n45 plus.n32 24.1005
R289 plus.n25 plus.n24 22.6399
R290 plus.n10 plus.n7 22.6399
R291 plus.n53 plus.n52 22.6399
R292 plus.n38 plus.n35 22.6399
R293 plus.n8 plus.n7 20.9576
R294 plus.n36 plus.n35 20.9576
R295 plus plus.n27 11.099
R296 plus.n20 plus.n19 0.730803
R297 plus.n13 plus.n12 0.730803
R298 plus.n48 plus.n47 0.730803
R299 plus.n41 plus.n40 0.730803
R300 plus.n9 plus.n6 0.189894
R301 plus.n6 plus.n5 0.189894
R302 plus.n14 plus.n5 0.189894
R303 plus.n15 plus.n14 0.189894
R304 plus.n16 plus.n15 0.189894
R305 plus.n16 plus.n3 0.189894
R306 plus.n3 plus.n2 0.189894
R307 plus.n21 plus.n2 0.189894
R308 plus.n22 plus.n21 0.189894
R309 plus.n23 plus.n22 0.189894
R310 plus.n23 plus.n0 0.189894
R311 plus.n27 plus.n0 0.189894
R312 plus.n55 plus.n28 0.189894
R313 plus.n51 plus.n28 0.189894
R314 plus.n51 plus.n50 0.189894
R315 plus.n50 plus.n49 0.189894
R316 plus.n49 plus.n30 0.189894
R317 plus.n31 plus.n30 0.189894
R318 plus.n44 plus.n31 0.189894
R319 plus.n44 plus.n43 0.189894
R320 plus.n43 plus.n42 0.189894
R321 plus.n42 plus.n33 0.189894
R322 plus.n34 plus.n33 0.189894
R323 plus.n37 plus.n34 0.189894
R324 drain_left.n10 drain_left.n8 66.2531
R325 drain_left.n6 drain_left.n4 66.2529
R326 drain_left.n2 drain_left.n0 66.2529
R327 drain_left.n14 drain_left.n13 65.5376
R328 drain_left.n12 drain_left.n11 65.5376
R329 drain_left.n10 drain_left.n9 65.5376
R330 drain_left.n16 drain_left.n15 65.5374
R331 drain_left.n7 drain_left.n3 65.5373
R332 drain_left.n6 drain_left.n5 65.5373
R333 drain_left.n2 drain_left.n1 65.5373
R334 drain_left drain_left.n7 30.8185
R335 drain_left drain_left.n16 6.36873
R336 drain_left.n3 drain_left.t13 2.2005
R337 drain_left.n3 drain_left.t3 2.2005
R338 drain_left.n4 drain_left.t7 2.2005
R339 drain_left.n4 drain_left.t8 2.2005
R340 drain_left.n5 drain_left.t4 2.2005
R341 drain_left.n5 drain_left.t18 2.2005
R342 drain_left.n1 drain_left.t6 2.2005
R343 drain_left.n1 drain_left.t19 2.2005
R344 drain_left.n0 drain_left.t14 2.2005
R345 drain_left.n0 drain_left.t15 2.2005
R346 drain_left.n15 drain_left.t17 2.2005
R347 drain_left.n15 drain_left.t10 2.2005
R348 drain_left.n13 drain_left.t11 2.2005
R349 drain_left.n13 drain_left.t2 2.2005
R350 drain_left.n11 drain_left.t5 2.2005
R351 drain_left.n11 drain_left.t0 2.2005
R352 drain_left.n9 drain_left.t1 2.2005
R353 drain_left.n9 drain_left.t12 2.2005
R354 drain_left.n8 drain_left.t16 2.2005
R355 drain_left.n8 drain_left.t9 2.2005
R356 drain_left.n12 drain_left.n10 0.716017
R357 drain_left.n14 drain_left.n12 0.716017
R358 drain_left.n16 drain_left.n14 0.716017
R359 drain_left.n7 drain_left.n6 0.660671
R360 drain_left.n7 drain_left.n2 0.660671
C0 drain_right minus 7.841701f
C1 drain_right plus 0.40825f
C2 drain_right drain_left 1.35855f
C3 drain_right source 22.4794f
C4 plus minus 5.76443f
C5 minus drain_left 0.173163f
C6 minus source 7.93556f
C7 plus drain_left 8.09345f
C8 plus source 7.9496f
C9 source drain_left 22.4781f
C10 drain_right a_n2542_n2688# 6.434259f
C11 drain_left a_n2542_n2688# 6.80727f
C12 source a_n2542_n2688# 7.482327f
C13 minus a_n2542_n2688# 9.917062f
C14 plus a_n2542_n2688# 11.664531f
C15 drain_left.t14 a_n2542_n2688# 0.208951f
C16 drain_left.t15 a_n2542_n2688# 0.208951f
C17 drain_left.n0 a_n2542_n2688# 1.83176f
C18 drain_left.t6 a_n2542_n2688# 0.208951f
C19 drain_left.t19 a_n2542_n2688# 0.208951f
C20 drain_left.n1 a_n2542_n2688# 1.82763f
C21 drain_left.n2 a_n2542_n2688# 0.745112f
C22 drain_left.t13 a_n2542_n2688# 0.208951f
C23 drain_left.t3 a_n2542_n2688# 0.208951f
C24 drain_left.n3 a_n2542_n2688# 1.82763f
C25 drain_left.t7 a_n2542_n2688# 0.208951f
C26 drain_left.t8 a_n2542_n2688# 0.208951f
C27 drain_left.n4 a_n2542_n2688# 1.83176f
C28 drain_left.t4 a_n2542_n2688# 0.208951f
C29 drain_left.t18 a_n2542_n2688# 0.208951f
C30 drain_left.n5 a_n2542_n2688# 1.82763f
C31 drain_left.n6 a_n2542_n2688# 0.745112f
C32 drain_left.n7 a_n2542_n2688# 1.77124f
C33 drain_left.t16 a_n2542_n2688# 0.208951f
C34 drain_left.t9 a_n2542_n2688# 0.208951f
C35 drain_left.n8 a_n2542_n2688# 1.83176f
C36 drain_left.t1 a_n2542_n2688# 0.208951f
C37 drain_left.t12 a_n2542_n2688# 0.208951f
C38 drain_left.n9 a_n2542_n2688# 1.82763f
C39 drain_left.n10 a_n2542_n2688# 0.749313f
C40 drain_left.t5 a_n2542_n2688# 0.208951f
C41 drain_left.t0 a_n2542_n2688# 0.208951f
C42 drain_left.n11 a_n2542_n2688# 1.82763f
C43 drain_left.n12 a_n2542_n2688# 0.370806f
C44 drain_left.t11 a_n2542_n2688# 0.208951f
C45 drain_left.t2 a_n2542_n2688# 0.208951f
C46 drain_left.n13 a_n2542_n2688# 1.82763f
C47 drain_left.n14 a_n2542_n2688# 0.370806f
C48 drain_left.t17 a_n2542_n2688# 0.208951f
C49 drain_left.t10 a_n2542_n2688# 0.208951f
C50 drain_left.n15 a_n2542_n2688# 1.82762f
C51 drain_left.n16 a_n2542_n2688# 0.623227f
C52 plus.n0 a_n2542_n2688# 0.044935f
C53 plus.t9 a_n2542_n2688# 0.579907f
C54 plus.t2 a_n2542_n2688# 0.579907f
C55 plus.t17 a_n2542_n2688# 0.579907f
C56 plus.n1 a_n2542_n2688# 0.251864f
C57 plus.n2 a_n2542_n2688# 0.044935f
C58 plus.t8 a_n2542_n2688# 0.579907f
C59 plus.t19 a_n2542_n2688# 0.579907f
C60 plus.n3 a_n2542_n2688# 0.044935f
C61 plus.t14 a_n2542_n2688# 0.579907f
C62 plus.n4 a_n2542_n2688# 0.251726f
C63 plus.n5 a_n2542_n2688# 0.044935f
C64 plus.t7 a_n2542_n2688# 0.579907f
C65 plus.t18 a_n2542_n2688# 0.579907f
C66 plus.n6 a_n2542_n2688# 0.044935f
C67 plus.t10 a_n2542_n2688# 0.579907f
C68 plus.n7 a_n2542_n2688# 0.251449f
C69 plus.t3 a_n2542_n2688# 0.589632f
C70 plus.n8 a_n2542_n2688# 0.237774f
C71 plus.n9 a_n2542_n2688# 0.147482f
C72 plus.n10 a_n2542_n2688# 0.010197f
C73 plus.n11 a_n2542_n2688# 0.251864f
C74 plus.n12 a_n2542_n2688# 0.010197f
C75 plus.n13 a_n2542_n2688# 0.247293f
C76 plus.n14 a_n2542_n2688# 0.044935f
C77 plus.n15 a_n2542_n2688# 0.044935f
C78 plus.n16 a_n2542_n2688# 0.044935f
C79 plus.n17 a_n2542_n2688# 0.010197f
C80 plus.n18 a_n2542_n2688# 0.251726f
C81 plus.n19 a_n2542_n2688# 0.247293f
C82 plus.n20 a_n2542_n2688# 0.010197f
C83 plus.n21 a_n2542_n2688# 0.044935f
C84 plus.n22 a_n2542_n2688# 0.044935f
C85 plus.n23 a_n2542_n2688# 0.044935f
C86 plus.n24 a_n2542_n2688# 0.010197f
C87 plus.n25 a_n2542_n2688# 0.251449f
C88 plus.n26 a_n2542_n2688# 0.247155f
C89 plus.n27 a_n2542_n2688# 0.451335f
C90 plus.n28 a_n2542_n2688# 0.044935f
C91 plus.t5 a_n2542_n2688# 0.579907f
C92 plus.t4 a_n2542_n2688# 0.579907f
C93 plus.t13 a_n2542_n2688# 0.579907f
C94 plus.n29 a_n2542_n2688# 0.251864f
C95 plus.n30 a_n2542_n2688# 0.044935f
C96 plus.t0 a_n2542_n2688# 0.579907f
C97 plus.n31 a_n2542_n2688# 0.044935f
C98 plus.t6 a_n2542_n2688# 0.579907f
C99 plus.t16 a_n2542_n2688# 0.579907f
C100 plus.n32 a_n2542_n2688# 0.251726f
C101 plus.n33 a_n2542_n2688# 0.044935f
C102 plus.t15 a_n2542_n2688# 0.579907f
C103 plus.n34 a_n2542_n2688# 0.044935f
C104 plus.t1 a_n2542_n2688# 0.579907f
C105 plus.t12 a_n2542_n2688# 0.579907f
C106 plus.n35 a_n2542_n2688# 0.251449f
C107 plus.t11 a_n2542_n2688# 0.589632f
C108 plus.n36 a_n2542_n2688# 0.237774f
C109 plus.n37 a_n2542_n2688# 0.147482f
C110 plus.n38 a_n2542_n2688# 0.010197f
C111 plus.n39 a_n2542_n2688# 0.251864f
C112 plus.n40 a_n2542_n2688# 0.010197f
C113 plus.n41 a_n2542_n2688# 0.247293f
C114 plus.n42 a_n2542_n2688# 0.044935f
C115 plus.n43 a_n2542_n2688# 0.044935f
C116 plus.n44 a_n2542_n2688# 0.044935f
C117 plus.n45 a_n2542_n2688# 0.010197f
C118 plus.n46 a_n2542_n2688# 0.251726f
C119 plus.n47 a_n2542_n2688# 0.247293f
C120 plus.n48 a_n2542_n2688# 0.010197f
C121 plus.n49 a_n2542_n2688# 0.044935f
C122 plus.n50 a_n2542_n2688# 0.044935f
C123 plus.n51 a_n2542_n2688# 0.044935f
C124 plus.n52 a_n2542_n2688# 0.010197f
C125 plus.n53 a_n2542_n2688# 0.251449f
C126 plus.n54 a_n2542_n2688# 0.247155f
C127 plus.n55 a_n2542_n2688# 1.41711f
C128 drain_right.t0 a_n2542_n2688# 0.207683f
C129 drain_right.t1 a_n2542_n2688# 0.207683f
C130 drain_right.n0 a_n2542_n2688# 1.82064f
C131 drain_right.t11 a_n2542_n2688# 0.207683f
C132 drain_right.t13 a_n2542_n2688# 0.207683f
C133 drain_right.n1 a_n2542_n2688# 1.81653f
C134 drain_right.n2 a_n2542_n2688# 0.740588f
C135 drain_right.t18 a_n2542_n2688# 0.207683f
C136 drain_right.t9 a_n2542_n2688# 0.207683f
C137 drain_right.n3 a_n2542_n2688# 1.81653f
C138 drain_right.t2 a_n2542_n2688# 0.207683f
C139 drain_right.t6 a_n2542_n2688# 0.207683f
C140 drain_right.n4 a_n2542_n2688# 1.82064f
C141 drain_right.t10 a_n2542_n2688# 0.207683f
C142 drain_right.t16 a_n2542_n2688# 0.207683f
C143 drain_right.n5 a_n2542_n2688# 1.81653f
C144 drain_right.n6 a_n2542_n2688# 0.740588f
C145 drain_right.n7 a_n2542_n2688# 1.70107f
C146 drain_right.t17 a_n2542_n2688# 0.207683f
C147 drain_right.t5 a_n2542_n2688# 0.207683f
C148 drain_right.n8 a_n2542_n2688# 1.82064f
C149 drain_right.t3 a_n2542_n2688# 0.207683f
C150 drain_right.t12 a_n2542_n2688# 0.207683f
C151 drain_right.n9 a_n2542_n2688# 1.81654f
C152 drain_right.n10 a_n2542_n2688# 0.744771f
C153 drain_right.t8 a_n2542_n2688# 0.207683f
C154 drain_right.t14 a_n2542_n2688# 0.207683f
C155 drain_right.n11 a_n2542_n2688# 1.81654f
C156 drain_right.n12 a_n2542_n2688# 0.368555f
C157 drain_right.t7 a_n2542_n2688# 0.207683f
C158 drain_right.t19 a_n2542_n2688# 0.207683f
C159 drain_right.n13 a_n2542_n2688# 1.81654f
C160 drain_right.n14 a_n2542_n2688# 0.368555f
C161 drain_right.t15 a_n2542_n2688# 0.207683f
C162 drain_right.t4 a_n2542_n2688# 0.207683f
C163 drain_right.n15 a_n2542_n2688# 1.81654f
C164 drain_right.n16 a_n2542_n2688# 0.619436f
C165 source.t14 a_n2542_n2688# 1.99255f
C166 source.n0 a_n2542_n2688# 1.17019f
C167 source.t6 a_n2542_n2688# 0.186857f
C168 source.t7 a_n2542_n2688# 0.186857f
C169 source.n1 a_n2542_n2688# 1.56425f
C170 source.n2 a_n2542_n2688# 0.36602f
C171 source.t15 a_n2542_n2688# 0.186857f
C172 source.t11 a_n2542_n2688# 0.186857f
C173 source.n3 a_n2542_n2688# 1.56425f
C174 source.n4 a_n2542_n2688# 0.36602f
C175 source.t5 a_n2542_n2688# 0.186857f
C176 source.t18 a_n2542_n2688# 0.186857f
C177 source.n5 a_n2542_n2688# 1.56425f
C178 source.n6 a_n2542_n2688# 0.36602f
C179 source.t0 a_n2542_n2688# 0.186857f
C180 source.t12 a_n2542_n2688# 0.186857f
C181 source.n7 a_n2542_n2688# 1.56425f
C182 source.n8 a_n2542_n2688# 0.36602f
C183 source.t8 a_n2542_n2688# 1.99255f
C184 source.n9 a_n2542_n2688# 0.426528f
C185 source.t22 a_n2542_n2688# 1.99255f
C186 source.n10 a_n2542_n2688# 0.426528f
C187 source.t29 a_n2542_n2688# 0.186857f
C188 source.t35 a_n2542_n2688# 0.186857f
C189 source.n11 a_n2542_n2688# 1.56425f
C190 source.n12 a_n2542_n2688# 0.36602f
C191 source.t26 a_n2542_n2688# 0.186857f
C192 source.t28 a_n2542_n2688# 0.186857f
C193 source.n13 a_n2542_n2688# 1.56425f
C194 source.n14 a_n2542_n2688# 0.36602f
C195 source.t24 a_n2542_n2688# 0.186857f
C196 source.t25 a_n2542_n2688# 0.186857f
C197 source.n15 a_n2542_n2688# 1.56425f
C198 source.n16 a_n2542_n2688# 0.36602f
C199 source.t20 a_n2542_n2688# 0.186857f
C200 source.t36 a_n2542_n2688# 0.186857f
C201 source.n17 a_n2542_n2688# 1.56425f
C202 source.n18 a_n2542_n2688# 0.36602f
C203 source.t23 a_n2542_n2688# 1.99255f
C204 source.n19 a_n2542_n2688# 1.55671f
C205 source.t10 a_n2542_n2688# 1.99255f
C206 source.n20 a_n2542_n2688# 1.55671f
C207 source.t19 a_n2542_n2688# 0.186857f
C208 source.t1 a_n2542_n2688# 0.186857f
C209 source.n21 a_n2542_n2688# 1.56424f
C210 source.n22 a_n2542_n2688# 0.366025f
C211 source.t9 a_n2542_n2688# 0.186857f
C212 source.t3 a_n2542_n2688# 0.186857f
C213 source.n23 a_n2542_n2688# 1.56424f
C214 source.n24 a_n2542_n2688# 0.366025f
C215 source.t17 a_n2542_n2688# 0.186857f
C216 source.t4 a_n2542_n2688# 0.186857f
C217 source.n25 a_n2542_n2688# 1.56424f
C218 source.n26 a_n2542_n2688# 0.366025f
C219 source.t13 a_n2542_n2688# 0.186857f
C220 source.t2 a_n2542_n2688# 0.186857f
C221 source.n27 a_n2542_n2688# 1.56424f
C222 source.n28 a_n2542_n2688# 0.366025f
C223 source.t16 a_n2542_n2688# 1.99255f
C224 source.n29 a_n2542_n2688# 0.426533f
C225 source.t30 a_n2542_n2688# 1.99255f
C226 source.n30 a_n2542_n2688# 0.426533f
C227 source.t34 a_n2542_n2688# 0.186857f
C228 source.t31 a_n2542_n2688# 0.186857f
C229 source.n31 a_n2542_n2688# 1.56424f
C230 source.n32 a_n2542_n2688# 0.366025f
C231 source.t38 a_n2542_n2688# 0.186857f
C232 source.t37 a_n2542_n2688# 0.186857f
C233 source.n33 a_n2542_n2688# 1.56424f
C234 source.n34 a_n2542_n2688# 0.366025f
C235 source.t32 a_n2542_n2688# 0.186857f
C236 source.t21 a_n2542_n2688# 0.186857f
C237 source.n35 a_n2542_n2688# 1.56424f
C238 source.n36 a_n2542_n2688# 0.366025f
C239 source.t33 a_n2542_n2688# 0.186857f
C240 source.t39 a_n2542_n2688# 0.186857f
C241 source.n37 a_n2542_n2688# 1.56424f
C242 source.n38 a_n2542_n2688# 0.366025f
C243 source.t27 a_n2542_n2688# 1.99255f
C244 source.n39 a_n2542_n2688# 0.586445f
C245 source.n40 a_n2542_n2688# 1.37548f
C246 minus.n0 a_n2542_n2688# 0.044133f
C247 minus.t12 a_n2542_n2688# 0.569552f
C248 minus.n1 a_n2542_n2688# 0.247367f
C249 minus.n2 a_n2542_n2688# 0.044133f
C250 minus.n3 a_n2542_n2688# 0.010015f
C251 minus.t11 a_n2542_n2688# 0.569552f
C252 minus.n4 a_n2542_n2688# 0.044133f
C253 minus.t7 a_n2542_n2688# 0.569552f
C254 minus.n5 a_n2542_n2688# 0.247367f
C255 minus.t14 a_n2542_n2688# 0.579104f
C256 minus.n6 a_n2542_n2688# 0.233528f
C257 minus.t2 a_n2542_n2688# 0.569552f
C258 minus.n7 a_n2542_n2688# 0.246959f
C259 minus.n8 a_n2542_n2688# 0.010015f
C260 minus.n9 a_n2542_n2688# 0.144849f
C261 minus.n10 a_n2542_n2688# 0.044133f
C262 minus.n11 a_n2542_n2688# 0.044133f
C263 minus.n12 a_n2542_n2688# 0.010015f
C264 minus.t16 a_n2542_n2688# 0.569552f
C265 minus.n13 a_n2542_n2688# 0.242878f
C266 minus.t5 a_n2542_n2688# 0.569552f
C267 minus.n14 a_n2542_n2688# 0.247231f
C268 minus.n15 a_n2542_n2688# 0.044133f
C269 minus.n16 a_n2542_n2688# 0.044133f
C270 minus.n17 a_n2542_n2688# 0.044133f
C271 minus.n18 a_n2542_n2688# 0.247231f
C272 minus.t0 a_n2542_n2688# 0.569552f
C273 minus.n19 a_n2542_n2688# 0.242878f
C274 minus.n20 a_n2542_n2688# 0.010015f
C275 minus.n21 a_n2542_n2688# 0.044133f
C276 minus.n22 a_n2542_n2688# 0.044133f
C277 minus.n23 a_n2542_n2688# 0.044133f
C278 minus.n24 a_n2542_n2688# 0.010015f
C279 minus.t15 a_n2542_n2688# 0.569552f
C280 minus.n25 a_n2542_n2688# 0.246959f
C281 minus.t4 a_n2542_n2688# 0.569552f
C282 minus.n26 a_n2542_n2688# 0.242742f
C283 minus.n27 a_n2542_n2688# 1.58806f
C284 minus.n28 a_n2542_n2688# 0.044133f
C285 minus.t3 a_n2542_n2688# 0.569552f
C286 minus.n29 a_n2542_n2688# 0.247367f
C287 minus.n30 a_n2542_n2688# 0.044133f
C288 minus.n31 a_n2542_n2688# 0.010015f
C289 minus.n32 a_n2542_n2688# 0.044133f
C290 minus.t8 a_n2542_n2688# 0.569552f
C291 minus.n33 a_n2542_n2688# 0.247367f
C292 minus.t19 a_n2542_n2688# 0.579104f
C293 minus.n34 a_n2542_n2688# 0.233528f
C294 minus.t18 a_n2542_n2688# 0.569552f
C295 minus.n35 a_n2542_n2688# 0.246959f
C296 minus.n36 a_n2542_n2688# 0.010015f
C297 minus.n37 a_n2542_n2688# 0.144849f
C298 minus.n38 a_n2542_n2688# 0.044133f
C299 minus.n39 a_n2542_n2688# 0.044133f
C300 minus.n40 a_n2542_n2688# 0.010015f
C301 minus.t6 a_n2542_n2688# 0.569552f
C302 minus.n41 a_n2542_n2688# 0.242878f
C303 minus.t1 a_n2542_n2688# 0.569552f
C304 minus.n42 a_n2542_n2688# 0.247231f
C305 minus.n43 a_n2542_n2688# 0.044133f
C306 minus.n44 a_n2542_n2688# 0.044133f
C307 minus.n45 a_n2542_n2688# 0.044133f
C308 minus.t10 a_n2542_n2688# 0.569552f
C309 minus.n46 a_n2542_n2688# 0.247231f
C310 minus.t9 a_n2542_n2688# 0.569552f
C311 minus.n47 a_n2542_n2688# 0.242878f
C312 minus.n48 a_n2542_n2688# 0.010015f
C313 minus.n49 a_n2542_n2688# 0.044133f
C314 minus.n50 a_n2542_n2688# 0.044133f
C315 minus.n51 a_n2542_n2688# 0.044133f
C316 minus.n52 a_n2542_n2688# 0.010015f
C317 minus.t17 a_n2542_n2688# 0.569552f
C318 minus.n53 a_n2542_n2688# 0.246959f
C319 minus.t13 a_n2542_n2688# 0.569552f
C320 minus.n54 a_n2542_n2688# 0.242742f
C321 minus.n55 a_n2542_n2688# 0.297993f
C322 minus.n56 a_n2542_n2688# 1.92377f
.ends

