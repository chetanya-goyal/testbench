* NGSPICE file created from diffpair37.ext - technology: sky130A

.subckt diffpair37 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t26 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X1 drain_left.t14 plus.t1 source.t21 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X2 source.t12 minus.t0 drain_right.t15 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X3 drain_right.t14 minus.t1 source.t6 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X4 a_n1850_n1088# a_n1850_n1088# a_n1850_n1088# a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.3
X5 source.t14 minus.t2 drain_right.t13 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X6 source.t28 plus.t2 drain_left.t13 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X7 source.t27 plus.t3 drain_left.t12 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X8 source.t17 plus.t4 drain_left.t11 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X9 drain_right.t12 minus.t3 source.t15 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X10 drain_right.t11 minus.t4 source.t11 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X11 drain_left.t10 plus.t5 source.t30 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X12 drain_right.t10 minus.t5 source.t2 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X13 source.t3 minus.t6 drain_right.t9 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X14 source.t20 plus.t6 drain_left.t9 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X15 source.t18 plus.t7 drain_left.t8 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X16 a_n1850_n1088# a_n1850_n1088# a_n1850_n1088# a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X17 drain_left.t7 plus.t8 source.t23 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X18 drain_left.t6 plus.t9 source.t24 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X19 source.t5 minus.t7 drain_right.t8 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X20 drain_right.t7 minus.t8 source.t8 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X21 source.t10 minus.t9 drain_right.t6 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X22 drain_left.t5 plus.t10 source.t16 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X23 a_n1850_n1088# a_n1850_n1088# a_n1850_n1088# a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X24 a_n1850_n1088# a_n1850_n1088# a_n1850_n1088# a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.3
X25 source.t25 plus.t11 drain_left.t4 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X26 source.t29 plus.t12 drain_left.t3 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X27 drain_right.t5 minus.t10 source.t0 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X28 drain_left.t2 plus.t13 source.t31 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X29 drain_right.t4 minus.t11 source.t1 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X30 drain_right.t3 minus.t12 source.t4 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.3
X31 source.t7 minus.t13 drain_right.t2 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X32 source.t9 minus.t14 drain_right.t1 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.3
X33 source.t13 minus.t15 drain_right.t0 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X34 source.t19 plus.t14 drain_left.t1 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
X35 drain_left.t0 plus.t15 source.t22 a_n1850_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.3
R0 plus.n5 plus.t4 214.709
R1 plus.n21 plus.t1 214.709
R2 plus.n28 plus.t9 214.709
R3 plus.n44 plus.t6 214.709
R4 plus.n6 plus.t8 184.768
R5 plus.n3 plus.t12 184.768
R6 plus.n12 plus.t15 184.768
R7 plus.n14 plus.t7 184.768
R8 plus.n1 plus.t10 184.768
R9 plus.n20 plus.t14 184.768
R10 plus.n29 plus.t2 184.768
R11 plus.n26 plus.t0 184.768
R12 plus.n35 plus.t11 184.768
R13 plus.n37 plus.t5 184.768
R14 plus.n24 plus.t3 184.768
R15 plus.n43 plus.t13 184.768
R16 plus.n5 plus.n4 161.489
R17 plus.n28 plus.n27 161.489
R18 plus.n7 plus.n4 161.3
R19 plus.n9 plus.n8 161.3
R20 plus.n11 plus.n10 161.3
R21 plus.n13 plus.n2 161.3
R22 plus.n16 plus.n15 161.3
R23 plus.n18 plus.n17 161.3
R24 plus.n19 plus.n0 161.3
R25 plus.n22 plus.n21 161.3
R26 plus.n30 plus.n27 161.3
R27 plus.n32 plus.n31 161.3
R28 plus.n34 plus.n33 161.3
R29 plus.n36 plus.n25 161.3
R30 plus.n39 plus.n38 161.3
R31 plus.n41 plus.n40 161.3
R32 plus.n42 plus.n23 161.3
R33 plus.n45 plus.n44 161.3
R34 plus.n8 plus.n7 73.0308
R35 plus.n19 plus.n18 73.0308
R36 plus.n42 plus.n41 73.0308
R37 plus.n31 plus.n30 73.0308
R38 plus.n11 plus.n3 64.9975
R39 plus.n15 plus.n1 64.9975
R40 plus.n38 plus.n24 64.9975
R41 plus.n34 plus.n26 64.9975
R42 plus.n6 plus.n5 62.0763
R43 plus.n21 plus.n20 62.0763
R44 plus.n44 plus.n43 62.0763
R45 plus.n29 plus.n28 62.0763
R46 plus.n13 plus.n12 46.0096
R47 plus.n14 plus.n13 46.0096
R48 plus.n37 plus.n36 46.0096
R49 plus.n36 plus.n35 46.0096
R50 plus.n12 plus.n11 27.0217
R51 plus.n15 plus.n14 27.0217
R52 plus.n38 plus.n37 27.0217
R53 plus.n35 plus.n34 27.0217
R54 plus plus.n45 25.8096
R55 plus.n7 plus.n6 10.955
R56 plus.n20 plus.n19 10.955
R57 plus.n43 plus.n42 10.955
R58 plus.n30 plus.n29 10.955
R59 plus.n8 plus.n3 8.03383
R60 plus.n18 plus.n1 8.03383
R61 plus.n41 plus.n24 8.03383
R62 plus.n31 plus.n26 8.03383
R63 plus plus.n22 7.94368
R64 plus.n9 plus.n4 0.189894
R65 plus.n10 plus.n9 0.189894
R66 plus.n10 plus.n2 0.189894
R67 plus.n16 plus.n2 0.189894
R68 plus.n17 plus.n16 0.189894
R69 plus.n17 plus.n0 0.189894
R70 plus.n22 plus.n0 0.189894
R71 plus.n45 plus.n23 0.189894
R72 plus.n40 plus.n23 0.189894
R73 plus.n40 plus.n39 0.189894
R74 plus.n39 plus.n25 0.189894
R75 plus.n33 plus.n25 0.189894
R76 plus.n33 plus.n32 0.189894
R77 plus.n32 plus.n27 0.189894
R78 source.n0 source.t21 243.255
R79 source.n7 source.t17 243.255
R80 source.n8 source.t8 243.255
R81 source.n15 source.t9 243.255
R82 source.n31 source.t4 243.254
R83 source.n24 source.t10 243.254
R84 source.n23 source.t24 243.254
R85 source.n16 source.t20 243.254
R86 source.n2 source.n1 223.454
R87 source.n4 source.n3 223.454
R88 source.n6 source.n5 223.454
R89 source.n10 source.n9 223.454
R90 source.n12 source.n11 223.454
R91 source.n14 source.n13 223.454
R92 source.n30 source.n29 223.453
R93 source.n28 source.n27 223.453
R94 source.n26 source.n25 223.453
R95 source.n22 source.n21 223.453
R96 source.n20 source.n19 223.453
R97 source.n18 source.n17 223.453
R98 source.n29 source.t11 19.8005
R99 source.n29 source.t13 19.8005
R100 source.n27 source.t0 19.8005
R101 source.n27 source.t3 19.8005
R102 source.n25 source.t15 19.8005
R103 source.n25 source.t14 19.8005
R104 source.n21 source.t26 19.8005
R105 source.n21 source.t28 19.8005
R106 source.n19 source.t30 19.8005
R107 source.n19 source.t25 19.8005
R108 source.n17 source.t31 19.8005
R109 source.n17 source.t27 19.8005
R110 source.n1 source.t16 19.8005
R111 source.n1 source.t19 19.8005
R112 source.n3 source.t22 19.8005
R113 source.n3 source.t18 19.8005
R114 source.n5 source.t23 19.8005
R115 source.n5 source.t29 19.8005
R116 source.n9 source.t6 19.8005
R117 source.n9 source.t7 19.8005
R118 source.n11 source.t1 19.8005
R119 source.n11 source.t5 19.8005
R120 source.n13 source.t2 19.8005
R121 source.n13 source.t12 19.8005
R122 source.n16 source.n15 13.4975
R123 source.n32 source.n0 7.96301
R124 source.n32 source.n31 5.53498
R125 source.n15 source.n14 0.543603
R126 source.n14 source.n12 0.543603
R127 source.n12 source.n10 0.543603
R128 source.n10 source.n8 0.543603
R129 source.n7 source.n6 0.543603
R130 source.n6 source.n4 0.543603
R131 source.n4 source.n2 0.543603
R132 source.n2 source.n0 0.543603
R133 source.n18 source.n16 0.543603
R134 source.n20 source.n18 0.543603
R135 source.n22 source.n20 0.543603
R136 source.n23 source.n22 0.543603
R137 source.n26 source.n24 0.543603
R138 source.n28 source.n26 0.543603
R139 source.n30 source.n28 0.543603
R140 source.n31 source.n30 0.543603
R141 source.n8 source.n7 0.470328
R142 source.n24 source.n23 0.470328
R143 source source.n32 0.188
R144 drain_left.n9 drain_left.n7 240.675
R145 drain_left.n5 drain_left.n3 240.674
R146 drain_left.n2 drain_left.n0 240.674
R147 drain_left.n13 drain_left.n12 240.132
R148 drain_left.n11 drain_left.n10 240.132
R149 drain_left.n9 drain_left.n8 240.132
R150 drain_left.n5 drain_left.n4 240.131
R151 drain_left.n2 drain_left.n1 240.131
R152 drain_left drain_left.n6 22.5639
R153 drain_left.n3 drain_left.t13 19.8005
R154 drain_left.n3 drain_left.t6 19.8005
R155 drain_left.n4 drain_left.t4 19.8005
R156 drain_left.n4 drain_left.t15 19.8005
R157 drain_left.n1 drain_left.t12 19.8005
R158 drain_left.n1 drain_left.t10 19.8005
R159 drain_left.n0 drain_left.t9 19.8005
R160 drain_left.n0 drain_left.t2 19.8005
R161 drain_left.n12 drain_left.t1 19.8005
R162 drain_left.n12 drain_left.t14 19.8005
R163 drain_left.n10 drain_left.t8 19.8005
R164 drain_left.n10 drain_left.t5 19.8005
R165 drain_left.n8 drain_left.t3 19.8005
R166 drain_left.n8 drain_left.t0 19.8005
R167 drain_left.n7 drain_left.t11 19.8005
R168 drain_left.n7 drain_left.t7 19.8005
R169 drain_left drain_left.n13 6.19632
R170 drain_left.n11 drain_left.n9 0.543603
R171 drain_left.n13 drain_left.n11 0.543603
R172 drain_left.n6 drain_left.n5 0.216706
R173 drain_left.n6 drain_left.n2 0.216706
R174 minus.n21 minus.t14 214.709
R175 minus.n5 minus.t8 214.709
R176 minus.n44 minus.t12 214.709
R177 minus.n28 minus.t9 214.709
R178 minus.n20 minus.t5 184.768
R179 minus.n1 minus.t0 184.768
R180 minus.n14 minus.t11 184.768
R181 minus.n12 minus.t7 184.768
R182 minus.n3 minus.t1 184.768
R183 minus.n6 minus.t13 184.768
R184 minus.n43 minus.t15 184.768
R185 minus.n24 minus.t4 184.768
R186 minus.n37 minus.t6 184.768
R187 minus.n35 minus.t10 184.768
R188 minus.n26 minus.t2 184.768
R189 minus.n29 minus.t3 184.768
R190 minus.n5 minus.n4 161.489
R191 minus.n28 minus.n27 161.489
R192 minus.n22 minus.n21 161.3
R193 minus.n19 minus.n0 161.3
R194 minus.n18 minus.n17 161.3
R195 minus.n16 minus.n15 161.3
R196 minus.n13 minus.n2 161.3
R197 minus.n11 minus.n10 161.3
R198 minus.n9 minus.n8 161.3
R199 minus.n7 minus.n4 161.3
R200 minus.n45 minus.n44 161.3
R201 minus.n42 minus.n23 161.3
R202 minus.n41 minus.n40 161.3
R203 minus.n39 minus.n38 161.3
R204 minus.n36 minus.n25 161.3
R205 minus.n34 minus.n33 161.3
R206 minus.n32 minus.n31 161.3
R207 minus.n30 minus.n27 161.3
R208 minus.n19 minus.n18 73.0308
R209 minus.n8 minus.n7 73.0308
R210 minus.n31 minus.n30 73.0308
R211 minus.n42 minus.n41 73.0308
R212 minus.n15 minus.n1 64.9975
R213 minus.n11 minus.n3 64.9975
R214 minus.n34 minus.n26 64.9975
R215 minus.n38 minus.n24 64.9975
R216 minus.n21 minus.n20 62.0763
R217 minus.n6 minus.n5 62.0763
R218 minus.n29 minus.n28 62.0763
R219 minus.n44 minus.n43 62.0763
R220 minus.n14 minus.n13 46.0096
R221 minus.n13 minus.n12 46.0096
R222 minus.n36 minus.n35 46.0096
R223 minus.n37 minus.n36 46.0096
R224 minus.n46 minus.n22 27.7619
R225 minus.n15 minus.n14 27.0217
R226 minus.n12 minus.n11 27.0217
R227 minus.n35 minus.n34 27.0217
R228 minus.n38 minus.n37 27.0217
R229 minus.n20 minus.n19 10.955
R230 minus.n7 minus.n6 10.955
R231 minus.n30 minus.n29 10.955
R232 minus.n43 minus.n42 10.955
R233 minus.n18 minus.n1 8.03383
R234 minus.n8 minus.n3 8.03383
R235 minus.n31 minus.n26 8.03383
R236 minus.n41 minus.n24 8.03383
R237 minus.n46 minus.n45 6.46641
R238 minus.n22 minus.n0 0.189894
R239 minus.n17 minus.n0 0.189894
R240 minus.n17 minus.n16 0.189894
R241 minus.n16 minus.n2 0.189894
R242 minus.n10 minus.n2 0.189894
R243 minus.n10 minus.n9 0.189894
R244 minus.n9 minus.n4 0.189894
R245 minus.n32 minus.n27 0.189894
R246 minus.n33 minus.n32 0.189894
R247 minus.n33 minus.n25 0.189894
R248 minus.n39 minus.n25 0.189894
R249 minus.n40 minus.n39 0.189894
R250 minus.n40 minus.n23 0.189894
R251 minus.n45 minus.n23 0.189894
R252 minus minus.n46 0.188
R253 drain_right.n9 drain_right.n7 240.675
R254 drain_right.n5 drain_right.n3 240.674
R255 drain_right.n2 drain_right.n0 240.674
R256 drain_right.n9 drain_right.n8 240.132
R257 drain_right.n11 drain_right.n10 240.132
R258 drain_right.n13 drain_right.n12 240.132
R259 drain_right.n5 drain_right.n4 240.131
R260 drain_right.n2 drain_right.n1 240.131
R261 drain_right drain_right.n6 22.0107
R262 drain_right.n3 drain_right.t0 19.8005
R263 drain_right.n3 drain_right.t3 19.8005
R264 drain_right.n4 drain_right.t9 19.8005
R265 drain_right.n4 drain_right.t11 19.8005
R266 drain_right.n1 drain_right.t13 19.8005
R267 drain_right.n1 drain_right.t5 19.8005
R268 drain_right.n0 drain_right.t6 19.8005
R269 drain_right.n0 drain_right.t12 19.8005
R270 drain_right.n7 drain_right.t2 19.8005
R271 drain_right.n7 drain_right.t7 19.8005
R272 drain_right.n8 drain_right.t8 19.8005
R273 drain_right.n8 drain_right.t14 19.8005
R274 drain_right.n10 drain_right.t15 19.8005
R275 drain_right.n10 drain_right.t4 19.8005
R276 drain_right.n12 drain_right.t1 19.8005
R277 drain_right.n12 drain_right.t10 19.8005
R278 drain_right drain_right.n13 6.19632
R279 drain_right.n13 drain_right.n11 0.543603
R280 drain_right.n11 drain_right.n9 0.543603
R281 drain_right.n6 drain_right.n5 0.216706
R282 drain_right.n6 drain_right.n2 0.216706
C0 plus source 1.28f
C1 minus source 1.26614f
C2 drain_right plus 0.342764f
C3 drain_left source 5.12185f
C4 drain_right minus 0.964167f
C5 drain_right drain_left 0.948789f
C6 plus minus 3.43566f
C7 plus drain_left 1.1438f
C8 drain_left minus 0.178898f
C9 drain_right source 5.12208f
C10 drain_right a_n1850_n1088# 3.67031f
C11 drain_left a_n1850_n1088# 3.91657f
C12 source a_n1850_n1088# 2.524018f
C13 minus a_n1850_n1088# 6.333418f
C14 plus a_n1850_n1088# 6.985127f
C15 drain_right.t6 a_n1850_n1088# 0.019855f
C16 drain_right.t12 a_n1850_n1088# 0.019855f
C17 drain_right.n0 a_n1850_n1088# 0.077768f
C18 drain_right.t13 a_n1850_n1088# 0.019855f
C19 drain_right.t5 a_n1850_n1088# 0.019855f
C20 drain_right.n1 a_n1850_n1088# 0.07715f
C21 drain_right.n2 a_n1850_n1088# 0.51302f
C22 drain_right.t0 a_n1850_n1088# 0.019855f
C23 drain_right.t3 a_n1850_n1088# 0.019855f
C24 drain_right.n3 a_n1850_n1088# 0.077768f
C25 drain_right.t9 a_n1850_n1088# 0.019855f
C26 drain_right.t11 a_n1850_n1088# 0.019855f
C27 drain_right.n4 a_n1850_n1088# 0.07715f
C28 drain_right.n5 a_n1850_n1088# 0.51302f
C29 drain_right.n6 a_n1850_n1088# 0.628292f
C30 drain_right.t2 a_n1850_n1088# 0.019855f
C31 drain_right.t7 a_n1850_n1088# 0.019855f
C32 drain_right.n7 a_n1850_n1088# 0.077768f
C33 drain_right.t8 a_n1850_n1088# 0.019855f
C34 drain_right.t14 a_n1850_n1088# 0.019855f
C35 drain_right.n8 a_n1850_n1088# 0.077151f
C36 drain_right.n9 a_n1850_n1088# 0.536791f
C37 drain_right.t15 a_n1850_n1088# 0.019855f
C38 drain_right.t4 a_n1850_n1088# 0.019855f
C39 drain_right.n10 a_n1850_n1088# 0.077151f
C40 drain_right.n11 a_n1850_n1088# 0.263645f
C41 drain_right.t1 a_n1850_n1088# 0.019855f
C42 drain_right.t10 a_n1850_n1088# 0.019855f
C43 drain_right.n12 a_n1850_n1088# 0.077151f
C44 drain_right.n13 a_n1850_n1088# 0.472779f
C45 minus.n0 a_n1850_n1088# 0.030544f
C46 minus.t14 a_n1850_n1088# 0.03232f
C47 minus.t5 a_n1850_n1088# 0.028248f
C48 minus.t0 a_n1850_n1088# 0.028248f
C49 minus.n1 a_n1850_n1088# 0.029104f
C50 minus.n2 a_n1850_n1088# 0.030544f
C51 minus.t11 a_n1850_n1088# 0.028248f
C52 minus.t7 a_n1850_n1088# 0.028248f
C53 minus.t1 a_n1850_n1088# 0.028248f
C54 minus.n3 a_n1850_n1088# 0.029104f
C55 minus.n4 a_n1850_n1088# 0.065003f
C56 minus.t13 a_n1850_n1088# 0.028248f
C57 minus.t8 a_n1850_n1088# 0.03232f
C58 minus.n5 a_n1850_n1088# 0.037747f
C59 minus.n6 a_n1850_n1088# 0.029104f
C60 minus.n7 a_n1850_n1088# 0.011545f
C61 minus.n8 a_n1850_n1088# 0.011168f
C62 minus.n9 a_n1850_n1088# 0.030544f
C63 minus.n10 a_n1850_n1088# 0.030544f
C64 minus.n11 a_n1850_n1088# 0.012581f
C65 minus.n12 a_n1850_n1088# 0.029104f
C66 minus.n13 a_n1850_n1088# 0.012581f
C67 minus.n14 a_n1850_n1088# 0.029104f
C68 minus.n15 a_n1850_n1088# 0.012581f
C69 minus.n16 a_n1850_n1088# 0.030544f
C70 minus.n17 a_n1850_n1088# 0.030544f
C71 minus.n18 a_n1850_n1088# 0.011168f
C72 minus.n19 a_n1850_n1088# 0.011545f
C73 minus.n20 a_n1850_n1088# 0.029104f
C74 minus.n21 a_n1850_n1088# 0.037707f
C75 minus.n22 a_n1850_n1088# 0.693141f
C76 minus.n23 a_n1850_n1088# 0.030544f
C77 minus.t15 a_n1850_n1088# 0.028248f
C78 minus.t4 a_n1850_n1088# 0.028248f
C79 minus.n24 a_n1850_n1088# 0.029104f
C80 minus.n25 a_n1850_n1088# 0.030544f
C81 minus.t6 a_n1850_n1088# 0.028248f
C82 minus.t10 a_n1850_n1088# 0.028248f
C83 minus.t2 a_n1850_n1088# 0.028248f
C84 minus.n26 a_n1850_n1088# 0.029104f
C85 minus.n27 a_n1850_n1088# 0.065003f
C86 minus.t3 a_n1850_n1088# 0.028248f
C87 minus.t9 a_n1850_n1088# 0.03232f
C88 minus.n28 a_n1850_n1088# 0.037747f
C89 minus.n29 a_n1850_n1088# 0.029104f
C90 minus.n30 a_n1850_n1088# 0.011545f
C91 minus.n31 a_n1850_n1088# 0.011168f
C92 minus.n32 a_n1850_n1088# 0.030544f
C93 minus.n33 a_n1850_n1088# 0.030544f
C94 minus.n34 a_n1850_n1088# 0.012581f
C95 minus.n35 a_n1850_n1088# 0.029104f
C96 minus.n36 a_n1850_n1088# 0.012581f
C97 minus.n37 a_n1850_n1088# 0.029104f
C98 minus.n38 a_n1850_n1088# 0.012581f
C99 minus.n39 a_n1850_n1088# 0.030544f
C100 minus.n40 a_n1850_n1088# 0.030544f
C101 minus.n41 a_n1850_n1088# 0.011168f
C102 minus.n42 a_n1850_n1088# 0.011545f
C103 minus.n43 a_n1850_n1088# 0.029104f
C104 minus.t12 a_n1850_n1088# 0.03232f
C105 minus.n44 a_n1850_n1088# 0.037707f
C106 minus.n45 a_n1850_n1088# 0.19727f
C107 minus.n46 a_n1850_n1088# 0.858249f
C108 drain_left.t9 a_n1850_n1088# 0.01948f
C109 drain_left.t2 a_n1850_n1088# 0.01948f
C110 drain_left.n0 a_n1850_n1088# 0.076298f
C111 drain_left.t12 a_n1850_n1088# 0.01948f
C112 drain_left.t10 a_n1850_n1088# 0.01948f
C113 drain_left.n1 a_n1850_n1088# 0.075692f
C114 drain_left.n2 a_n1850_n1088# 0.50332f
C115 drain_left.t13 a_n1850_n1088# 0.01948f
C116 drain_left.t6 a_n1850_n1088# 0.01948f
C117 drain_left.n3 a_n1850_n1088# 0.076298f
C118 drain_left.t4 a_n1850_n1088# 0.01948f
C119 drain_left.t15 a_n1850_n1088# 0.01948f
C120 drain_left.n4 a_n1850_n1088# 0.075692f
C121 drain_left.n5 a_n1850_n1088# 0.50332f
C122 drain_left.n6 a_n1850_n1088# 0.664054f
C123 drain_left.t11 a_n1850_n1088# 0.01948f
C124 drain_left.t7 a_n1850_n1088# 0.01948f
C125 drain_left.n7 a_n1850_n1088# 0.076298f
C126 drain_left.t3 a_n1850_n1088# 0.01948f
C127 drain_left.t0 a_n1850_n1088# 0.01948f
C128 drain_left.n8 a_n1850_n1088# 0.075692f
C129 drain_left.n9 a_n1850_n1088# 0.526642f
C130 drain_left.t8 a_n1850_n1088# 0.01948f
C131 drain_left.t5 a_n1850_n1088# 0.01948f
C132 drain_left.n10 a_n1850_n1088# 0.075692f
C133 drain_left.n11 a_n1850_n1088# 0.25866f
C134 drain_left.t1 a_n1850_n1088# 0.01948f
C135 drain_left.t14 a_n1850_n1088# 0.01948f
C136 drain_left.n12 a_n1850_n1088# 0.075692f
C137 drain_left.n13 a_n1850_n1088# 0.46384f
C138 source.t21 a_n1850_n1088# 0.128364f
C139 source.n0 a_n1850_n1088# 0.551175f
C140 source.t16 a_n1850_n1088# 0.023063f
C141 source.t19 a_n1850_n1088# 0.023063f
C142 source.n1 a_n1850_n1088# 0.074796f
C143 source.n2 a_n1850_n1088# 0.281391f
C144 source.t22 a_n1850_n1088# 0.023063f
C145 source.t18 a_n1850_n1088# 0.023063f
C146 source.n3 a_n1850_n1088# 0.074796f
C147 source.n4 a_n1850_n1088# 0.281391f
C148 source.t23 a_n1850_n1088# 0.023063f
C149 source.t29 a_n1850_n1088# 0.023063f
C150 source.n5 a_n1850_n1088# 0.074796f
C151 source.n6 a_n1850_n1088# 0.281391f
C152 source.t17 a_n1850_n1088# 0.128364f
C153 source.n7 a_n1850_n1088# 0.28383f
C154 source.t8 a_n1850_n1088# 0.128364f
C155 source.n8 a_n1850_n1088# 0.28383f
C156 source.t6 a_n1850_n1088# 0.023063f
C157 source.t7 a_n1850_n1088# 0.023063f
C158 source.n9 a_n1850_n1088# 0.074796f
C159 source.n10 a_n1850_n1088# 0.281391f
C160 source.t1 a_n1850_n1088# 0.023063f
C161 source.t5 a_n1850_n1088# 0.023063f
C162 source.n11 a_n1850_n1088# 0.074796f
C163 source.n12 a_n1850_n1088# 0.281391f
C164 source.t2 a_n1850_n1088# 0.023063f
C165 source.t12 a_n1850_n1088# 0.023063f
C166 source.n13 a_n1850_n1088# 0.074796f
C167 source.n14 a_n1850_n1088# 0.281391f
C168 source.t9 a_n1850_n1088# 0.128364f
C169 source.n15 a_n1850_n1088# 0.785033f
C170 source.t20 a_n1850_n1088# 0.128364f
C171 source.n16 a_n1850_n1088# 0.785033f
C172 source.t31 a_n1850_n1088# 0.023063f
C173 source.t27 a_n1850_n1088# 0.023063f
C174 source.n17 a_n1850_n1088# 0.074796f
C175 source.n18 a_n1850_n1088# 0.281391f
C176 source.t30 a_n1850_n1088# 0.023063f
C177 source.t25 a_n1850_n1088# 0.023063f
C178 source.n19 a_n1850_n1088# 0.074796f
C179 source.n20 a_n1850_n1088# 0.281391f
C180 source.t26 a_n1850_n1088# 0.023063f
C181 source.t28 a_n1850_n1088# 0.023063f
C182 source.n21 a_n1850_n1088# 0.074796f
C183 source.n22 a_n1850_n1088# 0.281391f
C184 source.t24 a_n1850_n1088# 0.128364f
C185 source.n23 a_n1850_n1088# 0.283831f
C186 source.t10 a_n1850_n1088# 0.128364f
C187 source.n24 a_n1850_n1088# 0.283831f
C188 source.t15 a_n1850_n1088# 0.023063f
C189 source.t14 a_n1850_n1088# 0.023063f
C190 source.n25 a_n1850_n1088# 0.074796f
C191 source.n26 a_n1850_n1088# 0.281391f
C192 source.t0 a_n1850_n1088# 0.023063f
C193 source.t3 a_n1850_n1088# 0.023063f
C194 source.n27 a_n1850_n1088# 0.074796f
C195 source.n28 a_n1850_n1088# 0.281391f
C196 source.t11 a_n1850_n1088# 0.023063f
C197 source.t13 a_n1850_n1088# 0.023063f
C198 source.n29 a_n1850_n1088# 0.074796f
C199 source.n30 a_n1850_n1088# 0.281391f
C200 source.t4 a_n1850_n1088# 0.128364f
C201 source.n31 a_n1850_n1088# 0.448579f
C202 source.n32 a_n1850_n1088# 0.591072f
C203 plus.n0 a_n1850_n1088# 0.03111f
C204 plus.t14 a_n1850_n1088# 0.02877f
C205 plus.t10 a_n1850_n1088# 0.02877f
C206 plus.n1 a_n1850_n1088# 0.029642f
C207 plus.n2 a_n1850_n1088# 0.03111f
C208 plus.t7 a_n1850_n1088# 0.02877f
C209 plus.t15 a_n1850_n1088# 0.02877f
C210 plus.t12 a_n1850_n1088# 0.02877f
C211 plus.n3 a_n1850_n1088# 0.029642f
C212 plus.n4 a_n1850_n1088# 0.066206f
C213 plus.t8 a_n1850_n1088# 0.02877f
C214 plus.t4 a_n1850_n1088# 0.032918f
C215 plus.n5 a_n1850_n1088# 0.038446f
C216 plus.n6 a_n1850_n1088# 0.029642f
C217 plus.n7 a_n1850_n1088# 0.011759f
C218 plus.n8 a_n1850_n1088# 0.011375f
C219 plus.n9 a_n1850_n1088# 0.03111f
C220 plus.n10 a_n1850_n1088# 0.03111f
C221 plus.n11 a_n1850_n1088# 0.012814f
C222 plus.n12 a_n1850_n1088# 0.029642f
C223 plus.n13 a_n1850_n1088# 0.012814f
C224 plus.n14 a_n1850_n1088# 0.029642f
C225 plus.n15 a_n1850_n1088# 0.012814f
C226 plus.n16 a_n1850_n1088# 0.03111f
C227 plus.n17 a_n1850_n1088# 0.03111f
C228 plus.n18 a_n1850_n1088# 0.011375f
C229 plus.n19 a_n1850_n1088# 0.011759f
C230 plus.n20 a_n1850_n1088# 0.029642f
C231 plus.t1 a_n1850_n1088# 0.032918f
C232 plus.n21 a_n1850_n1088# 0.038405f
C233 plus.n22 a_n1850_n1088# 0.210688f
C234 plus.n23 a_n1850_n1088# 0.03111f
C235 plus.t6 a_n1850_n1088# 0.032918f
C236 plus.t13 a_n1850_n1088# 0.02877f
C237 plus.t3 a_n1850_n1088# 0.02877f
C238 plus.n24 a_n1850_n1088# 0.029642f
C239 plus.n25 a_n1850_n1088# 0.03111f
C240 plus.t5 a_n1850_n1088# 0.02877f
C241 plus.t11 a_n1850_n1088# 0.02877f
C242 plus.t0 a_n1850_n1088# 0.02877f
C243 plus.n26 a_n1850_n1088# 0.029642f
C244 plus.n27 a_n1850_n1088# 0.066206f
C245 plus.t2 a_n1850_n1088# 0.02877f
C246 plus.t9 a_n1850_n1088# 0.032918f
C247 plus.n28 a_n1850_n1088# 0.038446f
C248 plus.n29 a_n1850_n1088# 0.029642f
C249 plus.n30 a_n1850_n1088# 0.011759f
C250 plus.n31 a_n1850_n1088# 0.011375f
C251 plus.n32 a_n1850_n1088# 0.03111f
C252 plus.n33 a_n1850_n1088# 0.03111f
C253 plus.n34 a_n1850_n1088# 0.012814f
C254 plus.n35 a_n1850_n1088# 0.029642f
C255 plus.n36 a_n1850_n1088# 0.012814f
C256 plus.n37 a_n1850_n1088# 0.029642f
C257 plus.n38 a_n1850_n1088# 0.012814f
C258 plus.n39 a_n1850_n1088# 0.03111f
C259 plus.n40 a_n1850_n1088# 0.03111f
C260 plus.n41 a_n1850_n1088# 0.011375f
C261 plus.n42 a_n1850_n1088# 0.011759f
C262 plus.n43 a_n1850_n1088# 0.029642f
C263 plus.n44 a_n1850_n1088# 0.038405f
C264 plus.n45 a_n1850_n1088# 0.684579f
.ends

