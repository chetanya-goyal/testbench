* NGSPICE file created from diffpair484.ext - technology: sky130A

.subckt diffpair484 minus drain_right drain_left source plus
X0 a_n1496_n3888# a_n1496_n3888# a_n1496_n3888# a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=57 ps=247.6 w=15 l=0.15
X1 source.t19 minus.t0 drain_right.t4 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X2 drain_right.t8 minus.t1 source.t18 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X3 a_n1496_n3888# a_n1496_n3888# a_n1496_n3888# a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X4 a_n1496_n3888# a_n1496_n3888# a_n1496_n3888# a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X5 drain_left.t9 plus.t0 source.t2 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X6 source.t17 minus.t2 drain_right.t7 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X7 drain_right.t2 minus.t3 source.t16 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X8 drain_right.t3 minus.t4 source.t15 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X9 source.t6 plus.t1 drain_left.t8 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X10 source.t14 minus.t5 drain_right.t1 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X11 drain_right.t0 minus.t6 source.t13 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X12 drain_left.t7 plus.t2 source.t1 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X13 drain_right.t6 minus.t7 source.t12 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X14 drain_left.t6 plus.t3 source.t4 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X15 a_n1496_n3888# a_n1496_n3888# a_n1496_n3888# a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X16 source.t5 plus.t4 drain_left.t5 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X17 source.t11 minus.t8 drain_right.t5 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X18 drain_left.t4 plus.t5 source.t8 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=3.75 ps=15.5 w=15 l=0.15
X19 drain_left.t3 plus.t6 source.t7 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X20 source.t0 plus.t7 drain_left.t2 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X21 source.t9 plus.t8 drain_left.t1 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
X22 drain_left.t0 plus.t9 source.t3 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=7.125 ps=30.95 w=15 l=0.15
X23 drain_right.t9 minus.t9 source.t10 a_n1496_n3888# sky130_fd_pr__nfet_01v8 ad=3.75 pd=15.5 as=3.75 ps=15.5 w=15 l=0.15
R0 minus.n9 minus.t4 2662.68
R1 minus.n3 minus.t3 2662.68
R2 minus.n20 minus.t6 2662.68
R3 minus.n14 minus.t1 2662.68
R4 minus.n6 minus.t7 2618.87
R5 minus.n8 minus.t5 2618.87
R6 minus.n2 minus.t2 2618.87
R7 minus.n17 minus.t9 2618.87
R8 minus.n19 minus.t0 2618.87
R9 minus.n13 minus.t8 2618.87
R10 minus.n4 minus.n3 161.489
R11 minus.n15 minus.n14 161.489
R12 minus.n10 minus.n9 161.3
R13 minus.n7 minus.n0 161.3
R14 minus.n6 minus.n5 161.3
R15 minus.n4 minus.n1 161.3
R16 minus.n21 minus.n20 161.3
R17 minus.n18 minus.n11 161.3
R18 minus.n17 minus.n16 161.3
R19 minus.n15 minus.n12 161.3
R20 minus.n7 minus.n6 73.0308
R21 minus.n6 minus.n1 73.0308
R22 minus.n17 minus.n12 73.0308
R23 minus.n18 minus.n17 73.0308
R24 minus.n9 minus.n8 51.1217
R25 minus.n3 minus.n2 51.1217
R26 minus.n14 minus.n13 51.1217
R27 minus.n20 minus.n19 51.1217
R28 minus.n22 minus.n10 37.0744
R29 minus.n8 minus.n7 21.9096
R30 minus.n2 minus.n1 21.9096
R31 minus.n13 minus.n12 21.9096
R32 minus.n19 minus.n18 21.9096
R33 minus.n22 minus.n21 6.51376
R34 minus.n10 minus.n0 0.189894
R35 minus.n5 minus.n0 0.189894
R36 minus.n5 minus.n4 0.189894
R37 minus.n16 minus.n15 0.189894
R38 minus.n16 minus.n11 0.189894
R39 minus.n21 minus.n11 0.189894
R40 minus minus.n22 0.188
R41 drain_right.n1 drain_right.t8 63.4399
R42 drain_right.n7 drain_right.t3 62.8798
R43 drain_right.n6 drain_right.n4 61.44
R44 drain_right.n3 drain_right.n2 61.2445
R45 drain_right.n6 drain_right.n5 60.8798
R46 drain_right.n1 drain_right.n0 60.8796
R47 drain_right drain_right.n3 31.468
R48 drain_right drain_right.n7 5.93339
R49 drain_right.n2 drain_right.t4 2.0005
R50 drain_right.n2 drain_right.t0 2.0005
R51 drain_right.n0 drain_right.t5 2.0005
R52 drain_right.n0 drain_right.t9 2.0005
R53 drain_right.n4 drain_right.t7 2.0005
R54 drain_right.n4 drain_right.t2 2.0005
R55 drain_right.n5 drain_right.t1 2.0005
R56 drain_right.n5 drain_right.t6 2.0005
R57 drain_right.n7 drain_right.n6 0.560845
R58 drain_right.n3 drain_right.n1 0.0852402
R59 source.n5 source.t16 46.201
R60 source.n19 source.t13 46.2008
R61 source.n14 source.t4 46.2008
R62 source.n0 source.t3 46.2008
R63 source.n2 source.n1 44.201
R64 source.n4 source.n3 44.201
R65 source.n7 source.n6 44.201
R66 source.n9 source.n8 44.201
R67 source.n18 source.n17 44.2008
R68 source.n16 source.n15 44.2008
R69 source.n13 source.n12 44.2008
R70 source.n11 source.n10 44.2008
R71 source.n11 source.n9 24.6811
R72 source.n20 source.n0 18.5777
R73 source.n20 source.n19 5.5436
R74 source.n17 source.t10 2.0005
R75 source.n17 source.t19 2.0005
R76 source.n15 source.t18 2.0005
R77 source.n15 source.t11 2.0005
R78 source.n12 source.t2 2.0005
R79 source.n12 source.t9 2.0005
R80 source.n10 source.t8 2.0005
R81 source.n10 source.t6 2.0005
R82 source.n1 source.t7 2.0005
R83 source.n1 source.t5 2.0005
R84 source.n3 source.t1 2.0005
R85 source.n3 source.t0 2.0005
R86 source.n6 source.t12 2.0005
R87 source.n6 source.t17 2.0005
R88 source.n8 source.t15 2.0005
R89 source.n8 source.t14 2.0005
R90 source.n5 source.n4 0.7505
R91 source.n16 source.n14 0.7505
R92 source.n9 source.n7 0.560845
R93 source.n7 source.n5 0.560845
R94 source.n4 source.n2 0.560845
R95 source.n2 source.n0 0.560845
R96 source.n13 source.n11 0.560845
R97 source.n14 source.n13 0.560845
R98 source.n18 source.n16 0.560845
R99 source.n19 source.n18 0.560845
R100 source source.n20 0.188
R101 plus.n3 plus.t2 2662.68
R102 plus.n9 plus.t9 2662.68
R103 plus.n14 plus.t3 2662.68
R104 plus.n20 plus.t5 2662.68
R105 plus.n6 plus.t6 2618.87
R106 plus.n2 plus.t7 2618.87
R107 plus.n8 plus.t4 2618.87
R108 plus.n17 plus.t0 2618.87
R109 plus.n13 plus.t8 2618.87
R110 plus.n19 plus.t1 2618.87
R111 plus.n4 plus.n3 161.489
R112 plus.n15 plus.n14 161.489
R113 plus.n4 plus.n1 161.3
R114 plus.n6 plus.n5 161.3
R115 plus.n7 plus.n0 161.3
R116 plus.n10 plus.n9 161.3
R117 plus.n15 plus.n12 161.3
R118 plus.n17 plus.n16 161.3
R119 plus.n18 plus.n11 161.3
R120 plus.n21 plus.n20 161.3
R121 plus.n6 plus.n1 73.0308
R122 plus.n7 plus.n6 73.0308
R123 plus.n18 plus.n17 73.0308
R124 plus.n17 plus.n12 73.0308
R125 plus.n3 plus.n2 51.1217
R126 plus.n9 plus.n8 51.1217
R127 plus.n20 plus.n19 51.1217
R128 plus.n14 plus.n13 51.1217
R129 plus plus.n21 29.8191
R130 plus.n2 plus.n1 21.9096
R131 plus.n8 plus.n7 21.9096
R132 plus.n19 plus.n18 21.9096
R133 plus.n13 plus.n12 21.9096
R134 plus plus.n10 13.2941
R135 plus.n5 plus.n4 0.189894
R136 plus.n5 plus.n0 0.189894
R137 plus.n10 plus.n0 0.189894
R138 plus.n21 plus.n11 0.189894
R139 plus.n16 plus.n11 0.189894
R140 plus.n16 plus.n15 0.189894
R141 drain_left.n5 drain_left.t7 63.4402
R142 drain_left.n1 drain_left.t4 63.4399
R143 drain_left.n3 drain_left.n2 61.2445
R144 drain_left.n5 drain_left.n4 60.8798
R145 drain_left.n7 drain_left.n6 60.8796
R146 drain_left.n1 drain_left.n0 60.8796
R147 drain_left drain_left.n3 32.0213
R148 drain_left drain_left.n7 6.21356
R149 drain_left.n2 drain_left.t1 2.0005
R150 drain_left.n2 drain_left.t6 2.0005
R151 drain_left.n0 drain_left.t8 2.0005
R152 drain_left.n0 drain_left.t9 2.0005
R153 drain_left.n6 drain_left.t5 2.0005
R154 drain_left.n6 drain_left.t0 2.0005
R155 drain_left.n4 drain_left.t2 2.0005
R156 drain_left.n4 drain_left.t3 2.0005
R157 drain_left.n7 drain_left.n5 0.560845
R158 drain_left.n3 drain_left.n1 0.0852402
C0 source plus 2.38837f
C1 plus minus 5.55903f
C2 drain_right plus 0.299168f
C3 source drain_left 26.284302f
C4 minus drain_left 0.170828f
C5 drain_right drain_left 0.737656f
C6 source minus 2.37352f
C7 drain_right source 26.2711f
C8 plus drain_left 3.18817f
C9 drain_right minus 3.0487f
C10 drain_right a_n1496_n3888# 7.3842f
C11 drain_left a_n1496_n3888# 7.62695f
C12 source a_n1496_n3888# 7.20079f
C13 minus a_n1496_n3888# 5.702885f
C14 plus a_n1496_n3888# 8.122731f
C15 drain_left.t4 a_n1496_n3888# 3.75723f
C16 drain_left.t8 a_n1496_n3888# 0.457306f
C17 drain_left.t9 a_n1496_n3888# 0.457306f
C18 drain_left.n0 a_n1496_n3888# 3.03908f
C19 drain_left.n1 a_n1496_n3888# 0.63824f
C20 drain_left.t1 a_n1496_n3888# 0.457306f
C21 drain_left.t6 a_n1496_n3888# 0.457306f
C22 drain_left.n2 a_n1496_n3888# 3.04085f
C23 drain_left.n3 a_n1496_n3888# 1.62826f
C24 drain_left.t7 a_n1496_n3888# 3.75723f
C25 drain_left.t2 a_n1496_n3888# 0.457306f
C26 drain_left.t3 a_n1496_n3888# 0.457306f
C27 drain_left.n4 a_n1496_n3888# 3.03908f
C28 drain_left.n5 a_n1496_n3888# 0.670291f
C29 drain_left.t5 a_n1496_n3888# 0.457306f
C30 drain_left.t0 a_n1496_n3888# 0.457306f
C31 drain_left.n6 a_n1496_n3888# 3.03907f
C32 drain_left.n7 a_n1496_n3888# 0.513153f
C33 plus.n0 a_n1496_n3888# 0.059576f
C34 plus.t4 a_n1496_n3888# 0.378165f
C35 plus.t6 a_n1496_n3888# 0.378165f
C36 plus.n1 a_n1496_n3888# 0.025273f
C37 plus.t2 a_n1496_n3888# 0.380676f
C38 plus.t7 a_n1496_n3888# 0.378165f
C39 plus.n2 a_n1496_n3888# 0.154438f
C40 plus.n3 a_n1496_n3888# 0.175444f
C41 plus.n4 a_n1496_n3888# 0.128254f
C42 plus.n5 a_n1496_n3888# 0.059576f
C43 plus.n6 a_n1496_n3888# 0.174202f
C44 plus.n7 a_n1496_n3888# 0.025273f
C45 plus.n8 a_n1496_n3888# 0.154438f
C46 plus.t9 a_n1496_n3888# 0.380676f
C47 plus.n9 a_n1496_n3888# 0.175363f
C48 plus.n10 a_n1496_n3888# 0.754784f
C49 plus.n11 a_n1496_n3888# 0.059576f
C50 plus.t5 a_n1496_n3888# 0.380676f
C51 plus.t1 a_n1496_n3888# 0.378165f
C52 plus.t0 a_n1496_n3888# 0.378165f
C53 plus.n12 a_n1496_n3888# 0.025273f
C54 plus.t8 a_n1496_n3888# 0.378165f
C55 plus.n13 a_n1496_n3888# 0.154438f
C56 plus.t3 a_n1496_n3888# 0.380676f
C57 plus.n14 a_n1496_n3888# 0.175444f
C58 plus.n15 a_n1496_n3888# 0.128254f
C59 plus.n16 a_n1496_n3888# 0.059576f
C60 plus.n17 a_n1496_n3888# 0.174202f
C61 plus.n18 a_n1496_n3888# 0.025273f
C62 plus.n19 a_n1496_n3888# 0.154438f
C63 plus.n20 a_n1496_n3888# 0.175363f
C64 plus.n21 a_n1496_n3888# 1.79248f
C65 source.t3 a_n1496_n3888# 3.68516f
C66 source.n0 a_n1496_n3888# 1.64054f
C67 source.t7 a_n1496_n3888# 0.462815f
C68 source.t5 a_n1496_n3888# 0.462815f
C69 source.n1 a_n1496_n3888# 2.99791f
C70 source.n2 a_n1496_n3888# 0.34689f
C71 source.t1 a_n1496_n3888# 0.462815f
C72 source.t0 a_n1496_n3888# 0.462815f
C73 source.n3 a_n1496_n3888# 2.99791f
C74 source.n4 a_n1496_n3888# 0.362638f
C75 source.t16 a_n1496_n3888# 3.68517f
C76 source.n5 a_n1496_n3888# 0.508444f
C77 source.t12 a_n1496_n3888# 0.462815f
C78 source.t17 a_n1496_n3888# 0.462815f
C79 source.n6 a_n1496_n3888# 2.99791f
C80 source.n7 a_n1496_n3888# 0.34689f
C81 source.t15 a_n1496_n3888# 0.462815f
C82 source.t14 a_n1496_n3888# 0.462815f
C83 source.n8 a_n1496_n3888# 2.99791f
C84 source.n9 a_n1496_n3888# 1.97026f
C85 source.t8 a_n1496_n3888# 0.462815f
C86 source.t6 a_n1496_n3888# 0.462815f
C87 source.n10 a_n1496_n3888# 2.9979f
C88 source.n11 a_n1496_n3888# 1.97026f
C89 source.t2 a_n1496_n3888# 0.462815f
C90 source.t9 a_n1496_n3888# 0.462815f
C91 source.n12 a_n1496_n3888# 2.9979f
C92 source.n13 a_n1496_n3888# 0.346893f
C93 source.t4 a_n1496_n3888# 3.68516f
C94 source.n14 a_n1496_n3888# 0.508448f
C95 source.t18 a_n1496_n3888# 0.462815f
C96 source.t11 a_n1496_n3888# 0.462815f
C97 source.n15 a_n1496_n3888# 2.9979f
C98 source.n16 a_n1496_n3888# 0.362641f
C99 source.t10 a_n1496_n3888# 0.462815f
C100 source.t19 a_n1496_n3888# 0.462815f
C101 source.n17 a_n1496_n3888# 2.9979f
C102 source.n18 a_n1496_n3888# 0.346893f
C103 source.t13 a_n1496_n3888# 3.68516f
C104 source.n19 a_n1496_n3888# 0.631796f
C105 source.n20 a_n1496_n3888# 1.88507f
C106 drain_right.t8 a_n1496_n3888# 3.7444f
C107 drain_right.t5 a_n1496_n3888# 0.455744f
C108 drain_right.t9 a_n1496_n3888# 0.455744f
C109 drain_right.n0 a_n1496_n3888# 3.0287f
C110 drain_right.n1 a_n1496_n3888# 0.63606f
C111 drain_right.t4 a_n1496_n3888# 0.455744f
C112 drain_right.t0 a_n1496_n3888# 0.455744f
C113 drain_right.n2 a_n1496_n3888# 3.03046f
C114 drain_right.n3 a_n1496_n3888# 1.56956f
C115 drain_right.t7 a_n1496_n3888# 0.455744f
C116 drain_right.t2 a_n1496_n3888# 0.455744f
C117 drain_right.n4 a_n1496_n3888# 3.03152f
C118 drain_right.t1 a_n1496_n3888# 0.455744f
C119 drain_right.t6 a_n1496_n3888# 0.455744f
C120 drain_right.n5 a_n1496_n3888# 3.02871f
C121 drain_right.n6 a_n1496_n3888# 0.606358f
C122 drain_right.t3 a_n1496_n3888# 3.74111f
C123 drain_right.n7 a_n1496_n3888# 0.584593f
C124 minus.n0 a_n1496_n3888# 0.05789f
C125 minus.t4 a_n1496_n3888# 0.369899f
C126 minus.t5 a_n1496_n3888# 0.367459f
C127 minus.t7 a_n1496_n3888# 0.367459f
C128 minus.n1 a_n1496_n3888# 0.024558f
C129 minus.t2 a_n1496_n3888# 0.367459f
C130 minus.n2 a_n1496_n3888# 0.150066f
C131 minus.t3 a_n1496_n3888# 0.369899f
C132 minus.n3 a_n1496_n3888# 0.170477f
C133 minus.n4 a_n1496_n3888# 0.124624f
C134 minus.n5 a_n1496_n3888# 0.05789f
C135 minus.n6 a_n1496_n3888# 0.16927f
C136 minus.n7 a_n1496_n3888# 0.024558f
C137 minus.n8 a_n1496_n3888# 0.150066f
C138 minus.n9 a_n1496_n3888# 0.170399f
C139 minus.n10 a_n1496_n3888# 2.12443f
C140 minus.n11 a_n1496_n3888# 0.05789f
C141 minus.t0 a_n1496_n3888# 0.367459f
C142 minus.t9 a_n1496_n3888# 0.367459f
C143 minus.n12 a_n1496_n3888# 0.024558f
C144 minus.t1 a_n1496_n3888# 0.369899f
C145 minus.t8 a_n1496_n3888# 0.367459f
C146 minus.n13 a_n1496_n3888# 0.150066f
C147 minus.n14 a_n1496_n3888# 0.170477f
C148 minus.n15 a_n1496_n3888# 0.124624f
C149 minus.n16 a_n1496_n3888# 0.05789f
C150 minus.n17 a_n1496_n3888# 0.16927f
C151 minus.n18 a_n1496_n3888# 0.024558f
C152 minus.n19 a_n1496_n3888# 0.150066f
C153 minus.t6 a_n1496_n3888# 0.369899f
C154 minus.n20 a_n1496_n3888# 0.170399f
C155 minus.n21 a_n1496_n3888# 0.380342f
C156 minus.n22 a_n1496_n3888# 2.57327f
.ends

