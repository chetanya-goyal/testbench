* NGSPICE file created from diffpair303.ext - technology: sky130A

.subckt diffpair303 minus drain_right drain_left source plus
X0 a_n1746_n2088# a_n1746_n2088# a_n1746_n2088# a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.7
X1 source.t15 plus.t0 drain_left.t6 a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X2 source.t14 plus.t1 drain_left.t5 a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X3 source.t7 minus.t0 drain_right.t7 a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X4 source.t13 plus.t2 drain_left.t4 a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X5 drain_left.t3 plus.t3 source.t12 a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X6 drain_left.t1 plus.t4 source.t11 a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X7 drain_right.t6 minus.t1 source.t3 a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X8 source.t6 minus.t2 drain_right.t5 a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X9 source.t10 plus.t5 drain_left.t2 a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X10 drain_left.t7 plus.t6 source.t9 a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X11 a_n1746_n2088# a_n1746_n2088# a_n1746_n2088# a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X12 drain_right.t4 minus.t3 source.t5 a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X13 drain_right.t3 minus.t4 source.t4 a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.7
X14 drain_left.t0 plus.t7 source.t8 a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X15 a_n1746_n2088# a_n1746_n2088# a_n1746_n2088# a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X16 source.t0 minus.t5 drain_right.t2 a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
X17 drain_right.t1 minus.t6 source.t2 a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.7
X18 a_n1746_n2088# a_n1746_n2088# a_n1746_n2088# a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.7
X19 source.t1 minus.t7 drain_right.t0 a_n1746_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.7
R0 plus.n3 plus.t2 284.868
R1 plus.n13 plus.t4 284.868
R2 plus.n8 plus.t6 262.69
R3 plus.n6 plus.t1 262.69
R4 plus.n2 plus.t7 262.69
R5 plus.n18 plus.t0 262.69
R6 plus.n16 plus.t3 262.69
R7 plus.n12 plus.t5 262.69
R8 plus.n5 plus.n4 161.3
R9 plus.n6 plus.n1 161.3
R10 plus.n7 plus.n0 161.3
R11 plus.n9 plus.n8 161.3
R12 plus.n15 plus.n14 161.3
R13 plus.n16 plus.n11 161.3
R14 plus.n17 plus.n10 161.3
R15 plus.n19 plus.n18 161.3
R16 plus.n4 plus.n3 44.862
R17 plus.n14 plus.n13 44.862
R18 plus.n8 plus.n7 28.4823
R19 plus.n18 plus.n17 28.4823
R20 plus plus.n19 27.4763
R21 plus.n5 plus.n2 24.1005
R22 plus.n6 plus.n5 24.1005
R23 plus.n16 plus.n15 24.1005
R24 plus.n15 plus.n12 24.1005
R25 plus.n7 plus.n6 19.7187
R26 plus.n17 plus.n16 19.7187
R27 plus.n3 plus.n2 19.7081
R28 plus.n13 plus.n12 19.7081
R29 plus plus.n9 10.0043
R30 plus.n4 plus.n1 0.189894
R31 plus.n1 plus.n0 0.189894
R32 plus.n9 plus.n0 0.189894
R33 plus.n19 plus.n10 0.189894
R34 plus.n11 plus.n10 0.189894
R35 plus.n14 plus.n11 0.189894
R36 drain_left.n5 drain_left.n3 68.0787
R37 drain_left.n2 drain_left.n1 67.5793
R38 drain_left.n2 drain_left.n0 67.5793
R39 drain_left.n5 drain_left.n4 67.1907
R40 drain_left drain_left.n2 25.9294
R41 drain_left drain_left.n5 6.54115
R42 drain_left.n1 drain_left.t2 3.3005
R43 drain_left.n1 drain_left.t1 3.3005
R44 drain_left.n0 drain_left.t6 3.3005
R45 drain_left.n0 drain_left.t3 3.3005
R46 drain_left.n4 drain_left.t5 3.3005
R47 drain_left.n4 drain_left.t7 3.3005
R48 drain_left.n3 drain_left.t4 3.3005
R49 drain_left.n3 drain_left.t0 3.3005
R50 source.n258 source.n232 289.615
R51 source.n224 source.n198 289.615
R52 source.n192 source.n166 289.615
R53 source.n158 source.n132 289.615
R54 source.n26 source.n0 289.615
R55 source.n60 source.n34 289.615
R56 source.n92 source.n66 289.615
R57 source.n126 source.n100 289.615
R58 source.n243 source.n242 185
R59 source.n240 source.n239 185
R60 source.n249 source.n248 185
R61 source.n251 source.n250 185
R62 source.n236 source.n235 185
R63 source.n257 source.n256 185
R64 source.n259 source.n258 185
R65 source.n209 source.n208 185
R66 source.n206 source.n205 185
R67 source.n215 source.n214 185
R68 source.n217 source.n216 185
R69 source.n202 source.n201 185
R70 source.n223 source.n222 185
R71 source.n225 source.n224 185
R72 source.n177 source.n176 185
R73 source.n174 source.n173 185
R74 source.n183 source.n182 185
R75 source.n185 source.n184 185
R76 source.n170 source.n169 185
R77 source.n191 source.n190 185
R78 source.n193 source.n192 185
R79 source.n143 source.n142 185
R80 source.n140 source.n139 185
R81 source.n149 source.n148 185
R82 source.n151 source.n150 185
R83 source.n136 source.n135 185
R84 source.n157 source.n156 185
R85 source.n159 source.n158 185
R86 source.n27 source.n26 185
R87 source.n25 source.n24 185
R88 source.n4 source.n3 185
R89 source.n19 source.n18 185
R90 source.n17 source.n16 185
R91 source.n8 source.n7 185
R92 source.n11 source.n10 185
R93 source.n61 source.n60 185
R94 source.n59 source.n58 185
R95 source.n38 source.n37 185
R96 source.n53 source.n52 185
R97 source.n51 source.n50 185
R98 source.n42 source.n41 185
R99 source.n45 source.n44 185
R100 source.n93 source.n92 185
R101 source.n91 source.n90 185
R102 source.n70 source.n69 185
R103 source.n85 source.n84 185
R104 source.n83 source.n82 185
R105 source.n74 source.n73 185
R106 source.n77 source.n76 185
R107 source.n127 source.n126 185
R108 source.n125 source.n124 185
R109 source.n104 source.n103 185
R110 source.n119 source.n118 185
R111 source.n117 source.n116 185
R112 source.n108 source.n107 185
R113 source.n111 source.n110 185
R114 source.t5 source.n241 147.661
R115 source.t0 source.n207 147.661
R116 source.t11 source.n175 147.661
R117 source.t15 source.n141 147.661
R118 source.t9 source.n9 147.661
R119 source.t13 source.n43 147.661
R120 source.t4 source.n75 147.661
R121 source.t1 source.n109 147.661
R122 source.n242 source.n239 104.615
R123 source.n249 source.n239 104.615
R124 source.n250 source.n249 104.615
R125 source.n250 source.n235 104.615
R126 source.n257 source.n235 104.615
R127 source.n258 source.n257 104.615
R128 source.n208 source.n205 104.615
R129 source.n215 source.n205 104.615
R130 source.n216 source.n215 104.615
R131 source.n216 source.n201 104.615
R132 source.n223 source.n201 104.615
R133 source.n224 source.n223 104.615
R134 source.n176 source.n173 104.615
R135 source.n183 source.n173 104.615
R136 source.n184 source.n183 104.615
R137 source.n184 source.n169 104.615
R138 source.n191 source.n169 104.615
R139 source.n192 source.n191 104.615
R140 source.n142 source.n139 104.615
R141 source.n149 source.n139 104.615
R142 source.n150 source.n149 104.615
R143 source.n150 source.n135 104.615
R144 source.n157 source.n135 104.615
R145 source.n158 source.n157 104.615
R146 source.n26 source.n25 104.615
R147 source.n25 source.n3 104.615
R148 source.n18 source.n3 104.615
R149 source.n18 source.n17 104.615
R150 source.n17 source.n7 104.615
R151 source.n10 source.n7 104.615
R152 source.n60 source.n59 104.615
R153 source.n59 source.n37 104.615
R154 source.n52 source.n37 104.615
R155 source.n52 source.n51 104.615
R156 source.n51 source.n41 104.615
R157 source.n44 source.n41 104.615
R158 source.n92 source.n91 104.615
R159 source.n91 source.n69 104.615
R160 source.n84 source.n69 104.615
R161 source.n84 source.n83 104.615
R162 source.n83 source.n73 104.615
R163 source.n76 source.n73 104.615
R164 source.n126 source.n125 104.615
R165 source.n125 source.n103 104.615
R166 source.n118 source.n103 104.615
R167 source.n118 source.n117 104.615
R168 source.n117 source.n107 104.615
R169 source.n110 source.n107 104.615
R170 source.n242 source.t5 52.3082
R171 source.n208 source.t0 52.3082
R172 source.n176 source.t11 52.3082
R173 source.n142 source.t15 52.3082
R174 source.n10 source.t9 52.3082
R175 source.n44 source.t13 52.3082
R176 source.n76 source.t4 52.3082
R177 source.n110 source.t1 52.3082
R178 source.n33 source.n32 50.512
R179 source.n99 source.n98 50.512
R180 source.n231 source.n230 50.5119
R181 source.n165 source.n164 50.5119
R182 source.n263 source.n262 32.1853
R183 source.n229 source.n228 32.1853
R184 source.n197 source.n196 32.1853
R185 source.n163 source.n162 32.1853
R186 source.n31 source.n30 32.1853
R187 source.n65 source.n64 32.1853
R188 source.n97 source.n96 32.1853
R189 source.n131 source.n130 32.1853
R190 source.n163 source.n131 17.6302
R191 source.n243 source.n241 15.6674
R192 source.n209 source.n207 15.6674
R193 source.n177 source.n175 15.6674
R194 source.n143 source.n141 15.6674
R195 source.n11 source.n9 15.6674
R196 source.n45 source.n43 15.6674
R197 source.n77 source.n75 15.6674
R198 source.n111 source.n109 15.6674
R199 source.n244 source.n240 12.8005
R200 source.n210 source.n206 12.8005
R201 source.n178 source.n174 12.8005
R202 source.n144 source.n140 12.8005
R203 source.n12 source.n8 12.8005
R204 source.n46 source.n42 12.8005
R205 source.n78 source.n74 12.8005
R206 source.n112 source.n108 12.8005
R207 source.n248 source.n247 12.0247
R208 source.n214 source.n213 12.0247
R209 source.n182 source.n181 12.0247
R210 source.n148 source.n147 12.0247
R211 source.n16 source.n15 12.0247
R212 source.n50 source.n49 12.0247
R213 source.n82 source.n81 12.0247
R214 source.n116 source.n115 12.0247
R215 source.n264 source.n31 11.9233
R216 source.n251 source.n238 11.249
R217 source.n217 source.n204 11.249
R218 source.n185 source.n172 11.249
R219 source.n151 source.n138 11.249
R220 source.n19 source.n6 11.249
R221 source.n53 source.n40 11.249
R222 source.n85 source.n72 11.249
R223 source.n119 source.n106 11.249
R224 source.n252 source.n236 10.4732
R225 source.n218 source.n202 10.4732
R226 source.n186 source.n170 10.4732
R227 source.n152 source.n136 10.4732
R228 source.n20 source.n4 10.4732
R229 source.n54 source.n38 10.4732
R230 source.n86 source.n70 10.4732
R231 source.n120 source.n104 10.4732
R232 source.n256 source.n255 9.69747
R233 source.n222 source.n221 9.69747
R234 source.n190 source.n189 9.69747
R235 source.n156 source.n155 9.69747
R236 source.n24 source.n23 9.69747
R237 source.n58 source.n57 9.69747
R238 source.n90 source.n89 9.69747
R239 source.n124 source.n123 9.69747
R240 source.n262 source.n261 9.45567
R241 source.n228 source.n227 9.45567
R242 source.n196 source.n195 9.45567
R243 source.n162 source.n161 9.45567
R244 source.n30 source.n29 9.45567
R245 source.n64 source.n63 9.45567
R246 source.n96 source.n95 9.45567
R247 source.n130 source.n129 9.45567
R248 source.n261 source.n260 9.3005
R249 source.n234 source.n233 9.3005
R250 source.n255 source.n254 9.3005
R251 source.n253 source.n252 9.3005
R252 source.n238 source.n237 9.3005
R253 source.n247 source.n246 9.3005
R254 source.n245 source.n244 9.3005
R255 source.n227 source.n226 9.3005
R256 source.n200 source.n199 9.3005
R257 source.n221 source.n220 9.3005
R258 source.n219 source.n218 9.3005
R259 source.n204 source.n203 9.3005
R260 source.n213 source.n212 9.3005
R261 source.n211 source.n210 9.3005
R262 source.n195 source.n194 9.3005
R263 source.n168 source.n167 9.3005
R264 source.n189 source.n188 9.3005
R265 source.n187 source.n186 9.3005
R266 source.n172 source.n171 9.3005
R267 source.n181 source.n180 9.3005
R268 source.n179 source.n178 9.3005
R269 source.n161 source.n160 9.3005
R270 source.n134 source.n133 9.3005
R271 source.n155 source.n154 9.3005
R272 source.n153 source.n152 9.3005
R273 source.n138 source.n137 9.3005
R274 source.n147 source.n146 9.3005
R275 source.n145 source.n144 9.3005
R276 source.n29 source.n28 9.3005
R277 source.n2 source.n1 9.3005
R278 source.n23 source.n22 9.3005
R279 source.n21 source.n20 9.3005
R280 source.n6 source.n5 9.3005
R281 source.n15 source.n14 9.3005
R282 source.n13 source.n12 9.3005
R283 source.n63 source.n62 9.3005
R284 source.n36 source.n35 9.3005
R285 source.n57 source.n56 9.3005
R286 source.n55 source.n54 9.3005
R287 source.n40 source.n39 9.3005
R288 source.n49 source.n48 9.3005
R289 source.n47 source.n46 9.3005
R290 source.n95 source.n94 9.3005
R291 source.n68 source.n67 9.3005
R292 source.n89 source.n88 9.3005
R293 source.n87 source.n86 9.3005
R294 source.n72 source.n71 9.3005
R295 source.n81 source.n80 9.3005
R296 source.n79 source.n78 9.3005
R297 source.n129 source.n128 9.3005
R298 source.n102 source.n101 9.3005
R299 source.n123 source.n122 9.3005
R300 source.n121 source.n120 9.3005
R301 source.n106 source.n105 9.3005
R302 source.n115 source.n114 9.3005
R303 source.n113 source.n112 9.3005
R304 source.n259 source.n234 8.92171
R305 source.n225 source.n200 8.92171
R306 source.n193 source.n168 8.92171
R307 source.n159 source.n134 8.92171
R308 source.n27 source.n2 8.92171
R309 source.n61 source.n36 8.92171
R310 source.n93 source.n68 8.92171
R311 source.n127 source.n102 8.92171
R312 source.n260 source.n232 8.14595
R313 source.n226 source.n198 8.14595
R314 source.n194 source.n166 8.14595
R315 source.n160 source.n132 8.14595
R316 source.n28 source.n0 8.14595
R317 source.n62 source.n34 8.14595
R318 source.n94 source.n66 8.14595
R319 source.n128 source.n100 8.14595
R320 source.n262 source.n232 5.81868
R321 source.n228 source.n198 5.81868
R322 source.n196 source.n166 5.81868
R323 source.n162 source.n132 5.81868
R324 source.n30 source.n0 5.81868
R325 source.n64 source.n34 5.81868
R326 source.n96 source.n66 5.81868
R327 source.n130 source.n100 5.81868
R328 source.n264 source.n263 5.7074
R329 source.n260 source.n259 5.04292
R330 source.n226 source.n225 5.04292
R331 source.n194 source.n193 5.04292
R332 source.n160 source.n159 5.04292
R333 source.n28 source.n27 5.04292
R334 source.n62 source.n61 5.04292
R335 source.n94 source.n93 5.04292
R336 source.n128 source.n127 5.04292
R337 source.n245 source.n241 4.38594
R338 source.n211 source.n207 4.38594
R339 source.n179 source.n175 4.38594
R340 source.n145 source.n141 4.38594
R341 source.n13 source.n9 4.38594
R342 source.n47 source.n43 4.38594
R343 source.n79 source.n75 4.38594
R344 source.n113 source.n109 4.38594
R345 source.n256 source.n234 4.26717
R346 source.n222 source.n200 4.26717
R347 source.n190 source.n168 4.26717
R348 source.n156 source.n134 4.26717
R349 source.n24 source.n2 4.26717
R350 source.n58 source.n36 4.26717
R351 source.n90 source.n68 4.26717
R352 source.n124 source.n102 4.26717
R353 source.n255 source.n236 3.49141
R354 source.n221 source.n202 3.49141
R355 source.n189 source.n170 3.49141
R356 source.n155 source.n136 3.49141
R357 source.n23 source.n4 3.49141
R358 source.n57 source.n38 3.49141
R359 source.n89 source.n70 3.49141
R360 source.n123 source.n104 3.49141
R361 source.n230 source.t2 3.3005
R362 source.n230 source.t6 3.3005
R363 source.n164 source.t12 3.3005
R364 source.n164 source.t10 3.3005
R365 source.n32 source.t8 3.3005
R366 source.n32 source.t14 3.3005
R367 source.n98 source.t3 3.3005
R368 source.n98 source.t7 3.3005
R369 source.n252 source.n251 2.71565
R370 source.n218 source.n217 2.71565
R371 source.n186 source.n185 2.71565
R372 source.n152 source.n151 2.71565
R373 source.n20 source.n19 2.71565
R374 source.n54 source.n53 2.71565
R375 source.n86 source.n85 2.71565
R376 source.n120 source.n119 2.71565
R377 source.n248 source.n238 1.93989
R378 source.n214 source.n204 1.93989
R379 source.n182 source.n172 1.93989
R380 source.n148 source.n138 1.93989
R381 source.n16 source.n6 1.93989
R382 source.n50 source.n40 1.93989
R383 source.n82 source.n72 1.93989
R384 source.n116 source.n106 1.93989
R385 source.n247 source.n240 1.16414
R386 source.n213 source.n206 1.16414
R387 source.n181 source.n174 1.16414
R388 source.n147 source.n140 1.16414
R389 source.n15 source.n8 1.16414
R390 source.n49 source.n42 1.16414
R391 source.n81 source.n74 1.16414
R392 source.n115 source.n108 1.16414
R393 source.n131 source.n99 0.888431
R394 source.n99 source.n97 0.888431
R395 source.n65 source.n33 0.888431
R396 source.n33 source.n31 0.888431
R397 source.n165 source.n163 0.888431
R398 source.n197 source.n165 0.888431
R399 source.n231 source.n229 0.888431
R400 source.n263 source.n231 0.888431
R401 source.n97 source.n65 0.470328
R402 source.n229 source.n197 0.470328
R403 source.n244 source.n243 0.388379
R404 source.n210 source.n209 0.388379
R405 source.n178 source.n177 0.388379
R406 source.n144 source.n143 0.388379
R407 source.n12 source.n11 0.388379
R408 source.n46 source.n45 0.388379
R409 source.n78 source.n77 0.388379
R410 source.n112 source.n111 0.388379
R411 source source.n264 0.188
R412 source.n246 source.n245 0.155672
R413 source.n246 source.n237 0.155672
R414 source.n253 source.n237 0.155672
R415 source.n254 source.n253 0.155672
R416 source.n254 source.n233 0.155672
R417 source.n261 source.n233 0.155672
R418 source.n212 source.n211 0.155672
R419 source.n212 source.n203 0.155672
R420 source.n219 source.n203 0.155672
R421 source.n220 source.n219 0.155672
R422 source.n220 source.n199 0.155672
R423 source.n227 source.n199 0.155672
R424 source.n180 source.n179 0.155672
R425 source.n180 source.n171 0.155672
R426 source.n187 source.n171 0.155672
R427 source.n188 source.n187 0.155672
R428 source.n188 source.n167 0.155672
R429 source.n195 source.n167 0.155672
R430 source.n146 source.n145 0.155672
R431 source.n146 source.n137 0.155672
R432 source.n153 source.n137 0.155672
R433 source.n154 source.n153 0.155672
R434 source.n154 source.n133 0.155672
R435 source.n161 source.n133 0.155672
R436 source.n29 source.n1 0.155672
R437 source.n22 source.n1 0.155672
R438 source.n22 source.n21 0.155672
R439 source.n21 source.n5 0.155672
R440 source.n14 source.n5 0.155672
R441 source.n14 source.n13 0.155672
R442 source.n63 source.n35 0.155672
R443 source.n56 source.n35 0.155672
R444 source.n56 source.n55 0.155672
R445 source.n55 source.n39 0.155672
R446 source.n48 source.n39 0.155672
R447 source.n48 source.n47 0.155672
R448 source.n95 source.n67 0.155672
R449 source.n88 source.n67 0.155672
R450 source.n88 source.n87 0.155672
R451 source.n87 source.n71 0.155672
R452 source.n80 source.n71 0.155672
R453 source.n80 source.n79 0.155672
R454 source.n129 source.n101 0.155672
R455 source.n122 source.n101 0.155672
R456 source.n122 source.n121 0.155672
R457 source.n121 source.n105 0.155672
R458 source.n114 source.n105 0.155672
R459 source.n114 source.n113 0.155672
R460 minus.n3 minus.t4 284.868
R461 minus.n13 minus.t5 284.868
R462 minus.n2 minus.t0 262.69
R463 minus.n6 minus.t1 262.69
R464 minus.n8 minus.t7 262.69
R465 minus.n12 minus.t6 262.69
R466 minus.n16 minus.t2 262.69
R467 minus.n18 minus.t3 262.69
R468 minus.n9 minus.n8 161.3
R469 minus.n7 minus.n0 161.3
R470 minus.n6 minus.n5 161.3
R471 minus.n4 minus.n1 161.3
R472 minus.n19 minus.n18 161.3
R473 minus.n17 minus.n10 161.3
R474 minus.n16 minus.n15 161.3
R475 minus.n14 minus.n11 161.3
R476 minus.n4 minus.n3 44.862
R477 minus.n14 minus.n13 44.862
R478 minus.n20 minus.n9 31.3225
R479 minus.n8 minus.n7 28.4823
R480 minus.n18 minus.n17 28.4823
R481 minus.n6 minus.n1 24.1005
R482 minus.n2 minus.n1 24.1005
R483 minus.n12 minus.n11 24.1005
R484 minus.n16 minus.n11 24.1005
R485 minus.n7 minus.n6 19.7187
R486 minus.n17 minus.n16 19.7187
R487 minus.n3 minus.n2 19.7081
R488 minus.n13 minus.n12 19.7081
R489 minus.n20 minus.n19 6.63308
R490 minus.n9 minus.n0 0.189894
R491 minus.n5 minus.n0 0.189894
R492 minus.n5 minus.n4 0.189894
R493 minus.n15 minus.n14 0.189894
R494 minus.n15 minus.n10 0.189894
R495 minus.n19 minus.n10 0.189894
R496 minus minus.n20 0.188
R497 drain_right.n5 drain_right.n3 68.0786
R498 drain_right.n2 drain_right.n1 67.5793
R499 drain_right.n2 drain_right.n0 67.5793
R500 drain_right.n5 drain_right.n4 67.1908
R501 drain_right drain_right.n2 25.3761
R502 drain_right drain_right.n5 6.54115
R503 drain_right.n1 drain_right.t5 3.3005
R504 drain_right.n1 drain_right.t4 3.3005
R505 drain_right.n0 drain_right.t2 3.3005
R506 drain_right.n0 drain_right.t1 3.3005
R507 drain_right.n3 drain_right.t7 3.3005
R508 drain_right.n3 drain_right.t3 3.3005
R509 drain_right.n4 drain_right.t0 3.3005
R510 drain_right.n4 drain_right.t6 3.3005
C0 drain_left minus 0.171089f
C1 drain_left drain_right 0.821811f
C2 plus minus 4.2083f
C3 plus drain_right 0.322995f
C4 drain_left source 6.70116f
C5 plus source 3.03068f
C6 minus drain_right 2.96476f
C7 plus drain_left 3.1336f
C8 source minus 3.01666f
C9 source drain_right 6.70294f
C10 drain_right a_n1746_n2088# 4.49773f
C11 drain_left a_n1746_n2088# 4.74508f
C12 source a_n1746_n2088# 5.407554f
C13 minus a_n1746_n2088# 6.279799f
C14 plus a_n1746_n2088# 7.653199f
C15 drain_right.t2 a_n1746_n2088# 0.126599f
C16 drain_right.t1 a_n1746_n2088# 0.126599f
C17 drain_right.n0 a_n1746_n2088# 1.05779f
C18 drain_right.t5 a_n1746_n2088# 0.126599f
C19 drain_right.t4 a_n1746_n2088# 0.126599f
C20 drain_right.n1 a_n1746_n2088# 1.05779f
C21 drain_right.n2 a_n1746_n2088# 1.57692f
C22 drain_right.t7 a_n1746_n2088# 0.126599f
C23 drain_right.t3 a_n1746_n2088# 0.126599f
C24 drain_right.n3 a_n1746_n2088# 1.0608f
C25 drain_right.t0 a_n1746_n2088# 0.126599f
C26 drain_right.t6 a_n1746_n2088# 0.126599f
C27 drain_right.n4 a_n1746_n2088# 1.05584f
C28 drain_right.n5 a_n1746_n2088# 0.980966f
C29 minus.n0 a_n1746_n2088# 0.045134f
C30 minus.n1 a_n1746_n2088# 0.010242f
C31 minus.t1 a_n1746_n2088# 0.549837f
C32 minus.t4 a_n1746_n2088# 0.5696f
C33 minus.t0 a_n1746_n2088# 0.549837f
C34 minus.n2 a_n1746_n2088# 0.258159f
C35 minus.n3 a_n1746_n2088# 0.238465f
C36 minus.n4 a_n1746_n2088# 0.187689f
C37 minus.n5 a_n1746_n2088# 0.045134f
C38 minus.n6 a_n1746_n2088# 0.254074f
C39 minus.n7 a_n1746_n2088# 0.010242f
C40 minus.t7 a_n1746_n2088# 0.549837f
C41 minus.n8 a_n1746_n2088# 0.251152f
C42 minus.n9 a_n1746_n2088# 1.26823f
C43 minus.n10 a_n1746_n2088# 0.045134f
C44 minus.n11 a_n1746_n2088# 0.010242f
C45 minus.t5 a_n1746_n2088# 0.5696f
C46 minus.t6 a_n1746_n2088# 0.549837f
C47 minus.n12 a_n1746_n2088# 0.258159f
C48 minus.n13 a_n1746_n2088# 0.238465f
C49 minus.n14 a_n1746_n2088# 0.187689f
C50 minus.n15 a_n1746_n2088# 0.045134f
C51 minus.t2 a_n1746_n2088# 0.549837f
C52 minus.n16 a_n1746_n2088# 0.254074f
C53 minus.n17 a_n1746_n2088# 0.010242f
C54 minus.t3 a_n1746_n2088# 0.549837f
C55 minus.n18 a_n1746_n2088# 0.251152f
C56 minus.n19 a_n1746_n2088# 0.309137f
C57 minus.n20 a_n1746_n2088# 1.55419f
C58 source.n0 a_n1746_n2088# 0.030515f
C59 source.n1 a_n1746_n2088# 0.021709f
C60 source.n2 a_n1746_n2088# 0.011666f
C61 source.n3 a_n1746_n2088# 0.027573f
C62 source.n4 a_n1746_n2088# 0.012352f
C63 source.n5 a_n1746_n2088# 0.021709f
C64 source.n6 a_n1746_n2088# 0.011666f
C65 source.n7 a_n1746_n2088# 0.027573f
C66 source.n8 a_n1746_n2088# 0.012352f
C67 source.n9 a_n1746_n2088# 0.092901f
C68 source.t9 a_n1746_n2088# 0.044941f
C69 source.n10 a_n1746_n2088# 0.02068f
C70 source.n11 a_n1746_n2088# 0.016287f
C71 source.n12 a_n1746_n2088# 0.011666f
C72 source.n13 a_n1746_n2088# 0.516554f
C73 source.n14 a_n1746_n2088# 0.021709f
C74 source.n15 a_n1746_n2088# 0.011666f
C75 source.n16 a_n1746_n2088# 0.012352f
C76 source.n17 a_n1746_n2088# 0.027573f
C77 source.n18 a_n1746_n2088# 0.027573f
C78 source.n19 a_n1746_n2088# 0.012352f
C79 source.n20 a_n1746_n2088# 0.011666f
C80 source.n21 a_n1746_n2088# 0.021709f
C81 source.n22 a_n1746_n2088# 0.021709f
C82 source.n23 a_n1746_n2088# 0.011666f
C83 source.n24 a_n1746_n2088# 0.012352f
C84 source.n25 a_n1746_n2088# 0.027573f
C85 source.n26 a_n1746_n2088# 0.059692f
C86 source.n27 a_n1746_n2088# 0.012352f
C87 source.n28 a_n1746_n2088# 0.011666f
C88 source.n29 a_n1746_n2088# 0.05018f
C89 source.n30 a_n1746_n2088# 0.0334f
C90 source.n31 a_n1746_n2088# 0.567127f
C91 source.t8 a_n1746_n2088# 0.102932f
C92 source.t14 a_n1746_n2088# 0.102932f
C93 source.n32 a_n1746_n2088# 0.801647f
C94 source.n33 a_n1746_n2088# 0.327731f
C95 source.n34 a_n1746_n2088# 0.030515f
C96 source.n35 a_n1746_n2088# 0.021709f
C97 source.n36 a_n1746_n2088# 0.011666f
C98 source.n37 a_n1746_n2088# 0.027573f
C99 source.n38 a_n1746_n2088# 0.012352f
C100 source.n39 a_n1746_n2088# 0.021709f
C101 source.n40 a_n1746_n2088# 0.011666f
C102 source.n41 a_n1746_n2088# 0.027573f
C103 source.n42 a_n1746_n2088# 0.012352f
C104 source.n43 a_n1746_n2088# 0.092901f
C105 source.t13 a_n1746_n2088# 0.044941f
C106 source.n44 a_n1746_n2088# 0.02068f
C107 source.n45 a_n1746_n2088# 0.016287f
C108 source.n46 a_n1746_n2088# 0.011666f
C109 source.n47 a_n1746_n2088# 0.516554f
C110 source.n48 a_n1746_n2088# 0.021709f
C111 source.n49 a_n1746_n2088# 0.011666f
C112 source.n50 a_n1746_n2088# 0.012352f
C113 source.n51 a_n1746_n2088# 0.027573f
C114 source.n52 a_n1746_n2088# 0.027573f
C115 source.n53 a_n1746_n2088# 0.012352f
C116 source.n54 a_n1746_n2088# 0.011666f
C117 source.n55 a_n1746_n2088# 0.021709f
C118 source.n56 a_n1746_n2088# 0.021709f
C119 source.n57 a_n1746_n2088# 0.011666f
C120 source.n58 a_n1746_n2088# 0.012352f
C121 source.n59 a_n1746_n2088# 0.027573f
C122 source.n60 a_n1746_n2088# 0.059692f
C123 source.n61 a_n1746_n2088# 0.012352f
C124 source.n62 a_n1746_n2088# 0.011666f
C125 source.n63 a_n1746_n2088# 0.05018f
C126 source.n64 a_n1746_n2088# 0.0334f
C127 source.n65 a_n1746_n2088# 0.11352f
C128 source.n66 a_n1746_n2088# 0.030515f
C129 source.n67 a_n1746_n2088# 0.021709f
C130 source.n68 a_n1746_n2088# 0.011666f
C131 source.n69 a_n1746_n2088# 0.027573f
C132 source.n70 a_n1746_n2088# 0.012352f
C133 source.n71 a_n1746_n2088# 0.021709f
C134 source.n72 a_n1746_n2088# 0.011666f
C135 source.n73 a_n1746_n2088# 0.027573f
C136 source.n74 a_n1746_n2088# 0.012352f
C137 source.n75 a_n1746_n2088# 0.092901f
C138 source.t4 a_n1746_n2088# 0.044941f
C139 source.n76 a_n1746_n2088# 0.02068f
C140 source.n77 a_n1746_n2088# 0.016287f
C141 source.n78 a_n1746_n2088# 0.011666f
C142 source.n79 a_n1746_n2088# 0.516554f
C143 source.n80 a_n1746_n2088# 0.021709f
C144 source.n81 a_n1746_n2088# 0.011666f
C145 source.n82 a_n1746_n2088# 0.012352f
C146 source.n83 a_n1746_n2088# 0.027573f
C147 source.n84 a_n1746_n2088# 0.027573f
C148 source.n85 a_n1746_n2088# 0.012352f
C149 source.n86 a_n1746_n2088# 0.011666f
C150 source.n87 a_n1746_n2088# 0.021709f
C151 source.n88 a_n1746_n2088# 0.021709f
C152 source.n89 a_n1746_n2088# 0.011666f
C153 source.n90 a_n1746_n2088# 0.012352f
C154 source.n91 a_n1746_n2088# 0.027573f
C155 source.n92 a_n1746_n2088# 0.059692f
C156 source.n93 a_n1746_n2088# 0.012352f
C157 source.n94 a_n1746_n2088# 0.011666f
C158 source.n95 a_n1746_n2088# 0.05018f
C159 source.n96 a_n1746_n2088# 0.0334f
C160 source.n97 a_n1746_n2088# 0.11352f
C161 source.t3 a_n1746_n2088# 0.102932f
C162 source.t7 a_n1746_n2088# 0.102932f
C163 source.n98 a_n1746_n2088# 0.801647f
C164 source.n99 a_n1746_n2088# 0.327731f
C165 source.n100 a_n1746_n2088# 0.030515f
C166 source.n101 a_n1746_n2088# 0.021709f
C167 source.n102 a_n1746_n2088# 0.011666f
C168 source.n103 a_n1746_n2088# 0.027573f
C169 source.n104 a_n1746_n2088# 0.012352f
C170 source.n105 a_n1746_n2088# 0.021709f
C171 source.n106 a_n1746_n2088# 0.011666f
C172 source.n107 a_n1746_n2088# 0.027573f
C173 source.n108 a_n1746_n2088# 0.012352f
C174 source.n109 a_n1746_n2088# 0.092901f
C175 source.t1 a_n1746_n2088# 0.044941f
C176 source.n110 a_n1746_n2088# 0.02068f
C177 source.n111 a_n1746_n2088# 0.016287f
C178 source.n112 a_n1746_n2088# 0.011666f
C179 source.n113 a_n1746_n2088# 0.516554f
C180 source.n114 a_n1746_n2088# 0.021709f
C181 source.n115 a_n1746_n2088# 0.011666f
C182 source.n116 a_n1746_n2088# 0.012352f
C183 source.n117 a_n1746_n2088# 0.027573f
C184 source.n118 a_n1746_n2088# 0.027573f
C185 source.n119 a_n1746_n2088# 0.012352f
C186 source.n120 a_n1746_n2088# 0.011666f
C187 source.n121 a_n1746_n2088# 0.021709f
C188 source.n122 a_n1746_n2088# 0.021709f
C189 source.n123 a_n1746_n2088# 0.011666f
C190 source.n124 a_n1746_n2088# 0.012352f
C191 source.n125 a_n1746_n2088# 0.027573f
C192 source.n126 a_n1746_n2088# 0.059692f
C193 source.n127 a_n1746_n2088# 0.012352f
C194 source.n128 a_n1746_n2088# 0.011666f
C195 source.n129 a_n1746_n2088# 0.05018f
C196 source.n130 a_n1746_n2088# 0.0334f
C197 source.n131 a_n1746_n2088# 0.853573f
C198 source.n132 a_n1746_n2088# 0.030515f
C199 source.n133 a_n1746_n2088# 0.021709f
C200 source.n134 a_n1746_n2088# 0.011666f
C201 source.n135 a_n1746_n2088# 0.027573f
C202 source.n136 a_n1746_n2088# 0.012352f
C203 source.n137 a_n1746_n2088# 0.021709f
C204 source.n138 a_n1746_n2088# 0.011666f
C205 source.n139 a_n1746_n2088# 0.027573f
C206 source.n140 a_n1746_n2088# 0.012352f
C207 source.n141 a_n1746_n2088# 0.092901f
C208 source.t15 a_n1746_n2088# 0.044941f
C209 source.n142 a_n1746_n2088# 0.02068f
C210 source.n143 a_n1746_n2088# 0.016287f
C211 source.n144 a_n1746_n2088# 0.011666f
C212 source.n145 a_n1746_n2088# 0.516554f
C213 source.n146 a_n1746_n2088# 0.021709f
C214 source.n147 a_n1746_n2088# 0.011666f
C215 source.n148 a_n1746_n2088# 0.012352f
C216 source.n149 a_n1746_n2088# 0.027573f
C217 source.n150 a_n1746_n2088# 0.027573f
C218 source.n151 a_n1746_n2088# 0.012352f
C219 source.n152 a_n1746_n2088# 0.011666f
C220 source.n153 a_n1746_n2088# 0.021709f
C221 source.n154 a_n1746_n2088# 0.021709f
C222 source.n155 a_n1746_n2088# 0.011666f
C223 source.n156 a_n1746_n2088# 0.012352f
C224 source.n157 a_n1746_n2088# 0.027573f
C225 source.n158 a_n1746_n2088# 0.059692f
C226 source.n159 a_n1746_n2088# 0.012352f
C227 source.n160 a_n1746_n2088# 0.011666f
C228 source.n161 a_n1746_n2088# 0.05018f
C229 source.n162 a_n1746_n2088# 0.0334f
C230 source.n163 a_n1746_n2088# 0.853573f
C231 source.t12 a_n1746_n2088# 0.102932f
C232 source.t10 a_n1746_n2088# 0.102932f
C233 source.n164 a_n1746_n2088# 0.801641f
C234 source.n165 a_n1746_n2088# 0.327736f
C235 source.n166 a_n1746_n2088# 0.030515f
C236 source.n167 a_n1746_n2088# 0.021709f
C237 source.n168 a_n1746_n2088# 0.011666f
C238 source.n169 a_n1746_n2088# 0.027573f
C239 source.n170 a_n1746_n2088# 0.012352f
C240 source.n171 a_n1746_n2088# 0.021709f
C241 source.n172 a_n1746_n2088# 0.011666f
C242 source.n173 a_n1746_n2088# 0.027573f
C243 source.n174 a_n1746_n2088# 0.012352f
C244 source.n175 a_n1746_n2088# 0.092901f
C245 source.t11 a_n1746_n2088# 0.044941f
C246 source.n176 a_n1746_n2088# 0.02068f
C247 source.n177 a_n1746_n2088# 0.016287f
C248 source.n178 a_n1746_n2088# 0.011666f
C249 source.n179 a_n1746_n2088# 0.516554f
C250 source.n180 a_n1746_n2088# 0.021709f
C251 source.n181 a_n1746_n2088# 0.011666f
C252 source.n182 a_n1746_n2088# 0.012352f
C253 source.n183 a_n1746_n2088# 0.027573f
C254 source.n184 a_n1746_n2088# 0.027573f
C255 source.n185 a_n1746_n2088# 0.012352f
C256 source.n186 a_n1746_n2088# 0.011666f
C257 source.n187 a_n1746_n2088# 0.021709f
C258 source.n188 a_n1746_n2088# 0.021709f
C259 source.n189 a_n1746_n2088# 0.011666f
C260 source.n190 a_n1746_n2088# 0.012352f
C261 source.n191 a_n1746_n2088# 0.027573f
C262 source.n192 a_n1746_n2088# 0.059692f
C263 source.n193 a_n1746_n2088# 0.012352f
C264 source.n194 a_n1746_n2088# 0.011666f
C265 source.n195 a_n1746_n2088# 0.05018f
C266 source.n196 a_n1746_n2088# 0.0334f
C267 source.n197 a_n1746_n2088# 0.11352f
C268 source.n198 a_n1746_n2088# 0.030515f
C269 source.n199 a_n1746_n2088# 0.021709f
C270 source.n200 a_n1746_n2088# 0.011666f
C271 source.n201 a_n1746_n2088# 0.027573f
C272 source.n202 a_n1746_n2088# 0.012352f
C273 source.n203 a_n1746_n2088# 0.021709f
C274 source.n204 a_n1746_n2088# 0.011666f
C275 source.n205 a_n1746_n2088# 0.027573f
C276 source.n206 a_n1746_n2088# 0.012352f
C277 source.n207 a_n1746_n2088# 0.092901f
C278 source.t0 a_n1746_n2088# 0.044941f
C279 source.n208 a_n1746_n2088# 0.02068f
C280 source.n209 a_n1746_n2088# 0.016287f
C281 source.n210 a_n1746_n2088# 0.011666f
C282 source.n211 a_n1746_n2088# 0.516554f
C283 source.n212 a_n1746_n2088# 0.021709f
C284 source.n213 a_n1746_n2088# 0.011666f
C285 source.n214 a_n1746_n2088# 0.012352f
C286 source.n215 a_n1746_n2088# 0.027573f
C287 source.n216 a_n1746_n2088# 0.027573f
C288 source.n217 a_n1746_n2088# 0.012352f
C289 source.n218 a_n1746_n2088# 0.011666f
C290 source.n219 a_n1746_n2088# 0.021709f
C291 source.n220 a_n1746_n2088# 0.021709f
C292 source.n221 a_n1746_n2088# 0.011666f
C293 source.n222 a_n1746_n2088# 0.012352f
C294 source.n223 a_n1746_n2088# 0.027573f
C295 source.n224 a_n1746_n2088# 0.059692f
C296 source.n225 a_n1746_n2088# 0.012352f
C297 source.n226 a_n1746_n2088# 0.011666f
C298 source.n227 a_n1746_n2088# 0.05018f
C299 source.n228 a_n1746_n2088# 0.0334f
C300 source.n229 a_n1746_n2088# 0.11352f
C301 source.t2 a_n1746_n2088# 0.102932f
C302 source.t6 a_n1746_n2088# 0.102932f
C303 source.n230 a_n1746_n2088# 0.801641f
C304 source.n231 a_n1746_n2088# 0.327736f
C305 source.n232 a_n1746_n2088# 0.030515f
C306 source.n233 a_n1746_n2088# 0.021709f
C307 source.n234 a_n1746_n2088# 0.011666f
C308 source.n235 a_n1746_n2088# 0.027573f
C309 source.n236 a_n1746_n2088# 0.012352f
C310 source.n237 a_n1746_n2088# 0.021709f
C311 source.n238 a_n1746_n2088# 0.011666f
C312 source.n239 a_n1746_n2088# 0.027573f
C313 source.n240 a_n1746_n2088# 0.012352f
C314 source.n241 a_n1746_n2088# 0.092901f
C315 source.t5 a_n1746_n2088# 0.044941f
C316 source.n242 a_n1746_n2088# 0.02068f
C317 source.n243 a_n1746_n2088# 0.016287f
C318 source.n244 a_n1746_n2088# 0.011666f
C319 source.n245 a_n1746_n2088# 0.516554f
C320 source.n246 a_n1746_n2088# 0.021709f
C321 source.n247 a_n1746_n2088# 0.011666f
C322 source.n248 a_n1746_n2088# 0.012352f
C323 source.n249 a_n1746_n2088# 0.027573f
C324 source.n250 a_n1746_n2088# 0.027573f
C325 source.n251 a_n1746_n2088# 0.012352f
C326 source.n252 a_n1746_n2088# 0.011666f
C327 source.n253 a_n1746_n2088# 0.021709f
C328 source.n254 a_n1746_n2088# 0.021709f
C329 source.n255 a_n1746_n2088# 0.011666f
C330 source.n256 a_n1746_n2088# 0.012352f
C331 source.n257 a_n1746_n2088# 0.027573f
C332 source.n258 a_n1746_n2088# 0.059692f
C333 source.n259 a_n1746_n2088# 0.012352f
C334 source.n260 a_n1746_n2088# 0.011666f
C335 source.n261 a_n1746_n2088# 0.05018f
C336 source.n262 a_n1746_n2088# 0.0334f
C337 source.n263 a_n1746_n2088# 0.255131f
C338 source.n264 a_n1746_n2088# 0.90033f
C339 drain_left.t6 a_n1746_n2088# 0.126542f
C340 drain_left.t3 a_n1746_n2088# 0.126542f
C341 drain_left.n0 a_n1746_n2088# 1.05731f
C342 drain_left.t2 a_n1746_n2088# 0.126542f
C343 drain_left.t1 a_n1746_n2088# 0.126542f
C344 drain_left.n1 a_n1746_n2088# 1.05731f
C345 drain_left.n2 a_n1746_n2088# 1.63048f
C346 drain_left.t4 a_n1746_n2088# 0.126542f
C347 drain_left.t0 a_n1746_n2088# 0.126542f
C348 drain_left.n3 a_n1746_n2088# 1.06032f
C349 drain_left.t5 a_n1746_n2088# 0.126542f
C350 drain_left.t7 a_n1746_n2088# 0.126542f
C351 drain_left.n4 a_n1746_n2088# 1.05536f
C352 drain_left.n5 a_n1746_n2088# 0.98052f
C353 plus.n0 a_n1746_n2088# 0.045988f
C354 plus.t6 a_n1746_n2088# 0.560241f
C355 plus.t1 a_n1746_n2088# 0.560241f
C356 plus.n1 a_n1746_n2088# 0.045988f
C357 plus.t7 a_n1746_n2088# 0.560241f
C358 plus.n2 a_n1746_n2088# 0.263043f
C359 plus.t2 a_n1746_n2088# 0.580377f
C360 plus.n3 a_n1746_n2088# 0.242977f
C361 plus.n4 a_n1746_n2088# 0.19124f
C362 plus.n5 a_n1746_n2088# 0.010436f
C363 plus.n6 a_n1746_n2088# 0.258882f
C364 plus.n7 a_n1746_n2088# 0.010436f
C365 plus.n8 a_n1746_n2088# 0.255905f
C366 plus.n9 a_n1746_n2088# 0.40904f
C367 plus.n10 a_n1746_n2088# 0.045988f
C368 plus.t0 a_n1746_n2088# 0.560241f
C369 plus.n11 a_n1746_n2088# 0.045988f
C370 plus.t3 a_n1746_n2088# 0.560241f
C371 plus.t5 a_n1746_n2088# 0.560241f
C372 plus.n12 a_n1746_n2088# 0.263043f
C373 plus.t4 a_n1746_n2088# 0.580377f
C374 plus.n13 a_n1746_n2088# 0.242977f
C375 plus.n14 a_n1746_n2088# 0.19124f
C376 plus.n15 a_n1746_n2088# 0.010436f
C377 plus.n16 a_n1746_n2088# 0.258882f
C378 plus.n17 a_n1746_n2088# 0.010436f
C379 plus.n18 a_n1746_n2088# 0.255905f
C380 plus.n19 a_n1746_n2088# 1.16863f
.ends

