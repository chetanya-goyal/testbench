* NGSPICE file created from diffpair357.ext - technology: sky130A

.subckt diffpair357 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t19 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X1 source.t1 minus.t0 drain_right.t15 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X2 drain_left.t14 plus.t1 source.t22 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X3 drain_left.t13 plus.t2 source.t21 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X4 drain_right.t14 minus.t1 source.t8 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X5 a_n1850_n2688# a_n1850_n2688# a_n1850_n2688# a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.3
X6 a_n1850_n2688# a_n1850_n2688# a_n1850_n2688# a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X7 source.t31 plus.t3 drain_left.t12 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X8 source.t11 minus.t2 drain_right.t13 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X9 source.t6 minus.t3 drain_right.t12 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X10 drain_right.t11 minus.t4 source.t7 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X11 source.t18 plus.t4 drain_left.t11 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X12 source.t29 plus.t5 drain_left.t10 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X13 source.t28 plus.t6 drain_left.t9 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X14 source.t27 plus.t7 drain_left.t8 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X15 a_n1850_n2688# a_n1850_n2688# a_n1850_n2688# a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X16 drain_left.t7 plus.t8 source.t26 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X17 drain_right.t10 minus.t5 source.t12 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X18 drain_right.t9 minus.t6 source.t10 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X19 source.t13 minus.t7 drain_right.t8 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X20 drain_right.t7 minus.t8 source.t3 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X21 drain_right.t6 minus.t9 source.t0 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X22 source.t16 plus.t9 drain_left.t6 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X23 drain_right.t5 minus.t10 source.t2 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X24 drain_left.t5 plus.t10 source.t20 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X25 a_n1850_n2688# a_n1850_n2688# a_n1850_n2688# a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.3
X26 drain_left.t4 plus.t11 source.t23 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.3
X27 source.t24 plus.t12 drain_left.t3 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X28 drain_left.t2 plus.t13 source.t17 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X29 drain_right.t4 minus.t11 source.t4 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X30 source.t9 minus.t12 drain_right.t3 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X31 source.t5 minus.t13 drain_right.t2 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X32 source.t14 minus.t14 drain_right.t1 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X33 source.t15 minus.t15 drain_right.t0 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.3
X34 source.t25 plus.t14 drain_left.t1 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
X35 drain_left.t0 plus.t15 source.t30 a_n1850_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.3
R0 plus.n5 plus.t3 857.376
R1 plus.n21 plus.t0 857.376
R2 plus.n28 plus.t11 857.376
R3 plus.n44 plus.t9 857.376
R4 plus.n6 plus.t8 827.433
R5 plus.n3 plus.t12 827.433
R6 plus.n12 plus.t15 827.433
R7 plus.n14 plus.t5 827.433
R8 plus.n1 plus.t10 827.433
R9 plus.n20 plus.t14 827.433
R10 plus.n29 plus.t4 827.433
R11 plus.n26 plus.t13 827.433
R12 plus.n35 plus.t6 827.433
R13 plus.n37 plus.t1 827.433
R14 plus.n24 plus.t7 827.433
R15 plus.n43 plus.t2 827.433
R16 plus.n5 plus.n4 161.489
R17 plus.n28 plus.n27 161.489
R18 plus.n7 plus.n4 161.3
R19 plus.n9 plus.n8 161.3
R20 plus.n11 plus.n10 161.3
R21 plus.n13 plus.n2 161.3
R22 plus.n16 plus.n15 161.3
R23 plus.n18 plus.n17 161.3
R24 plus.n19 plus.n0 161.3
R25 plus.n22 plus.n21 161.3
R26 plus.n30 plus.n27 161.3
R27 plus.n32 plus.n31 161.3
R28 plus.n34 plus.n33 161.3
R29 plus.n36 plus.n25 161.3
R30 plus.n39 plus.n38 161.3
R31 plus.n41 plus.n40 161.3
R32 plus.n42 plus.n23 161.3
R33 plus.n45 plus.n44 161.3
R34 plus.n8 plus.n7 73.0308
R35 plus.n19 plus.n18 73.0308
R36 plus.n42 plus.n41 73.0308
R37 plus.n31 plus.n30 73.0308
R38 plus.n11 plus.n3 64.9975
R39 plus.n15 plus.n1 64.9975
R40 plus.n38 plus.n24 64.9975
R41 plus.n34 plus.n26 64.9975
R42 plus.n6 plus.n5 62.0763
R43 plus.n21 plus.n20 62.0763
R44 plus.n44 plus.n43 62.0763
R45 plus.n29 plus.n28 62.0763
R46 plus.n13 plus.n12 46.0096
R47 plus.n14 plus.n13 46.0096
R48 plus.n37 plus.n36 46.0096
R49 plus.n36 plus.n35 46.0096
R50 plus plus.n45 28.8399
R51 plus.n12 plus.n11 27.0217
R52 plus.n15 plus.n14 27.0217
R53 plus.n38 plus.n37 27.0217
R54 plus.n35 plus.n34 27.0217
R55 plus plus.n22 10.974
R56 plus.n7 plus.n6 10.955
R57 plus.n20 plus.n19 10.955
R58 plus.n43 plus.n42 10.955
R59 plus.n30 plus.n29 10.955
R60 plus.n8 plus.n3 8.03383
R61 plus.n18 plus.n1 8.03383
R62 plus.n41 plus.n24 8.03383
R63 plus.n31 plus.n26 8.03383
R64 plus.n9 plus.n4 0.189894
R65 plus.n10 plus.n9 0.189894
R66 plus.n10 plus.n2 0.189894
R67 plus.n16 plus.n2 0.189894
R68 plus.n17 plus.n16 0.189894
R69 plus.n17 plus.n0 0.189894
R70 plus.n22 plus.n0 0.189894
R71 plus.n45 plus.n23 0.189894
R72 plus.n40 plus.n23 0.189894
R73 plus.n40 plus.n39 0.189894
R74 plus.n39 plus.n25 0.189894
R75 plus.n33 plus.n25 0.189894
R76 plus.n33 plus.n32 0.189894
R77 plus.n32 plus.n27 0.189894
R78 source.n7 source.t31 51.0588
R79 source.n8 source.t2 51.0588
R80 source.n15 source.t5 51.0588
R81 source.n31 source.t3 51.0586
R82 source.n24 source.t15 51.0586
R83 source.n23 source.t23 51.0586
R84 source.n16 source.t16 51.0586
R85 source.n0 source.t19 51.0586
R86 source.n2 source.n1 48.8588
R87 source.n4 source.n3 48.8588
R88 source.n6 source.n5 48.8588
R89 source.n10 source.n9 48.8588
R90 source.n12 source.n11 48.8588
R91 source.n14 source.n13 48.8588
R92 source.n30 source.n29 48.8586
R93 source.n28 source.n27 48.8586
R94 source.n26 source.n25 48.8586
R95 source.n22 source.n21 48.8586
R96 source.n20 source.n19 48.8586
R97 source.n18 source.n17 48.8586
R98 source.n16 source.n15 19.5581
R99 source.n32 source.n0 14.0236
R100 source.n32 source.n31 5.53498
R101 source.n29 source.t0 2.2005
R102 source.n29 source.t11 2.2005
R103 source.n27 source.t12 2.2005
R104 source.n27 source.t6 2.2005
R105 source.n25 source.t10 2.2005
R106 source.n25 source.t14 2.2005
R107 source.n21 source.t17 2.2005
R108 source.n21 source.t18 2.2005
R109 source.n19 source.t22 2.2005
R110 source.n19 source.t28 2.2005
R111 source.n17 source.t21 2.2005
R112 source.n17 source.t27 2.2005
R113 source.n1 source.t20 2.2005
R114 source.n1 source.t25 2.2005
R115 source.n3 source.t30 2.2005
R116 source.n3 source.t29 2.2005
R117 source.n5 source.t26 2.2005
R118 source.n5 source.t24 2.2005
R119 source.n9 source.t8 2.2005
R120 source.n9 source.t9 2.2005
R121 source.n11 source.t4 2.2005
R122 source.n11 source.t13 2.2005
R123 source.n13 source.t7 2.2005
R124 source.n13 source.t1 2.2005
R125 source.n15 source.n14 0.543603
R126 source.n14 source.n12 0.543603
R127 source.n12 source.n10 0.543603
R128 source.n10 source.n8 0.543603
R129 source.n7 source.n6 0.543603
R130 source.n6 source.n4 0.543603
R131 source.n4 source.n2 0.543603
R132 source.n2 source.n0 0.543603
R133 source.n18 source.n16 0.543603
R134 source.n20 source.n18 0.543603
R135 source.n22 source.n20 0.543603
R136 source.n23 source.n22 0.543603
R137 source.n26 source.n24 0.543603
R138 source.n28 source.n26 0.543603
R139 source.n30 source.n28 0.543603
R140 source.n31 source.n30 0.543603
R141 source.n8 source.n7 0.470328
R142 source.n24 source.n23 0.470328
R143 source source.n32 0.188
R144 drain_left.n9 drain_left.n7 66.0807
R145 drain_left.n5 drain_left.n3 66.0804
R146 drain_left.n2 drain_left.n0 66.0804
R147 drain_left.n11 drain_left.n10 65.5376
R148 drain_left.n9 drain_left.n8 65.5376
R149 drain_left.n13 drain_left.n12 65.5374
R150 drain_left.n5 drain_left.n4 65.5373
R151 drain_left.n2 drain_left.n1 65.5373
R152 drain_left drain_left.n6 28.6245
R153 drain_left drain_left.n13 6.19632
R154 drain_left.n3 drain_left.t11 2.2005
R155 drain_left.n3 drain_left.t4 2.2005
R156 drain_left.n4 drain_left.t9 2.2005
R157 drain_left.n4 drain_left.t2 2.2005
R158 drain_left.n1 drain_left.t8 2.2005
R159 drain_left.n1 drain_left.t14 2.2005
R160 drain_left.n0 drain_left.t6 2.2005
R161 drain_left.n0 drain_left.t13 2.2005
R162 drain_left.n12 drain_left.t1 2.2005
R163 drain_left.n12 drain_left.t15 2.2005
R164 drain_left.n10 drain_left.t10 2.2005
R165 drain_left.n10 drain_left.t5 2.2005
R166 drain_left.n8 drain_left.t3 2.2005
R167 drain_left.n8 drain_left.t0 2.2005
R168 drain_left.n7 drain_left.t12 2.2005
R169 drain_left.n7 drain_left.t7 2.2005
R170 drain_left.n11 drain_left.n9 0.543603
R171 drain_left.n13 drain_left.n11 0.543603
R172 drain_left.n6 drain_left.n5 0.216706
R173 drain_left.n6 drain_left.n2 0.216706
R174 minus.n21 minus.t13 857.376
R175 minus.n5 minus.t10 857.376
R176 minus.n44 minus.t8 857.376
R177 minus.n28 minus.t15 857.376
R178 minus.n20 minus.t4 827.433
R179 minus.n1 minus.t0 827.433
R180 minus.n14 minus.t11 827.433
R181 minus.n12 minus.t7 827.433
R182 minus.n3 minus.t1 827.433
R183 minus.n6 minus.t12 827.433
R184 minus.n43 minus.t2 827.433
R185 minus.n24 minus.t9 827.433
R186 minus.n37 minus.t3 827.433
R187 minus.n35 minus.t5 827.433
R188 minus.n26 minus.t14 827.433
R189 minus.n29 minus.t6 827.433
R190 minus.n5 minus.n4 161.489
R191 minus.n28 minus.n27 161.489
R192 minus.n22 minus.n21 161.3
R193 minus.n19 minus.n0 161.3
R194 minus.n18 minus.n17 161.3
R195 minus.n16 minus.n15 161.3
R196 minus.n13 minus.n2 161.3
R197 minus.n11 minus.n10 161.3
R198 minus.n9 minus.n8 161.3
R199 minus.n7 minus.n4 161.3
R200 minus.n45 minus.n44 161.3
R201 minus.n42 minus.n23 161.3
R202 minus.n41 minus.n40 161.3
R203 minus.n39 minus.n38 161.3
R204 minus.n36 minus.n25 161.3
R205 minus.n34 minus.n33 161.3
R206 minus.n32 minus.n31 161.3
R207 minus.n30 minus.n27 161.3
R208 minus.n19 minus.n18 73.0308
R209 minus.n8 minus.n7 73.0308
R210 minus.n31 minus.n30 73.0308
R211 minus.n42 minus.n41 73.0308
R212 minus.n15 minus.n1 64.9975
R213 minus.n11 minus.n3 64.9975
R214 minus.n34 minus.n26 64.9975
R215 minus.n38 minus.n24 64.9975
R216 minus.n21 minus.n20 62.0763
R217 minus.n6 minus.n5 62.0763
R218 minus.n29 minus.n28 62.0763
R219 minus.n44 minus.n43 62.0763
R220 minus.n14 minus.n13 46.0096
R221 minus.n13 minus.n12 46.0096
R222 minus.n36 minus.n35 46.0096
R223 minus.n37 minus.n36 46.0096
R224 minus.n46 minus.n22 33.8225
R225 minus.n15 minus.n14 27.0217
R226 minus.n12 minus.n11 27.0217
R227 minus.n35 minus.n34 27.0217
R228 minus.n38 minus.n37 27.0217
R229 minus.n20 minus.n19 10.955
R230 minus.n7 minus.n6 10.955
R231 minus.n30 minus.n29 10.955
R232 minus.n43 minus.n42 10.955
R233 minus.n18 minus.n1 8.03383
R234 minus.n8 minus.n3 8.03383
R235 minus.n31 minus.n26 8.03383
R236 minus.n41 minus.n24 8.03383
R237 minus.n46 minus.n45 6.46641
R238 minus.n22 minus.n0 0.189894
R239 minus.n17 minus.n0 0.189894
R240 minus.n17 minus.n16 0.189894
R241 minus.n16 minus.n2 0.189894
R242 minus.n10 minus.n2 0.189894
R243 minus.n10 minus.n9 0.189894
R244 minus.n9 minus.n4 0.189894
R245 minus.n32 minus.n27 0.189894
R246 minus.n33 minus.n32 0.189894
R247 minus.n33 minus.n25 0.189894
R248 minus.n39 minus.n25 0.189894
R249 minus.n40 minus.n39 0.189894
R250 minus.n40 minus.n23 0.189894
R251 minus.n45 minus.n23 0.189894
R252 minus minus.n46 0.188
R253 drain_right.n9 drain_right.n7 66.0805
R254 drain_right.n5 drain_right.n3 66.0804
R255 drain_right.n2 drain_right.n0 66.0804
R256 drain_right.n9 drain_right.n8 65.5376
R257 drain_right.n11 drain_right.n10 65.5376
R258 drain_right.n13 drain_right.n12 65.5376
R259 drain_right.n5 drain_right.n4 65.5373
R260 drain_right.n2 drain_right.n1 65.5373
R261 drain_right drain_right.n6 28.0713
R262 drain_right drain_right.n13 6.19632
R263 drain_right.n3 drain_right.t13 2.2005
R264 drain_right.n3 drain_right.t7 2.2005
R265 drain_right.n4 drain_right.t12 2.2005
R266 drain_right.n4 drain_right.t6 2.2005
R267 drain_right.n1 drain_right.t1 2.2005
R268 drain_right.n1 drain_right.t10 2.2005
R269 drain_right.n0 drain_right.t0 2.2005
R270 drain_right.n0 drain_right.t9 2.2005
R271 drain_right.n7 drain_right.t3 2.2005
R272 drain_right.n7 drain_right.t5 2.2005
R273 drain_right.n8 drain_right.t8 2.2005
R274 drain_right.n8 drain_right.t14 2.2005
R275 drain_right.n10 drain_right.t15 2.2005
R276 drain_right.n10 drain_right.t4 2.2005
R277 drain_right.n12 drain_right.t2 2.2005
R278 drain_right.n12 drain_right.t11 2.2005
R279 drain_right.n13 drain_right.n11 0.543603
R280 drain_right.n11 drain_right.n9 0.543603
R281 drain_right.n6 drain_right.n5 0.216706
R282 drain_right.n6 drain_right.n2 0.216706
C0 drain_right minus 4.55062f
C1 drain_right drain_left 0.948737f
C2 plus minus 4.90753f
C3 plus drain_left 4.73032f
C4 drain_left minus 0.171647f
C5 drain_right source 23.5792f
C6 plus source 4.38549f
C7 minus source 4.37145f
C8 drain_right plus 0.334364f
C9 drain_left source 23.5789f
C10 drain_right a_n1850_n2688# 5.91935f
C11 drain_left a_n1850_n2688# 6.1986f
C12 source a_n1850_n2688# 7.096548f
C13 minus a_n1850_n2688# 7.029669f
C14 plus a_n1850_n2688# 8.80956f
C15 drain_right.t0 a_n1850_n2688# 0.239925f
C16 drain_right.t9 a_n1850_n2688# 0.239925f
C17 drain_right.n0 a_n1850_n2688# 2.10184f
C18 drain_right.t1 a_n1850_n2688# 0.239925f
C19 drain_right.t10 a_n1850_n2688# 0.239925f
C20 drain_right.n1 a_n1850_n2688# 2.09854f
C21 drain_right.n2 a_n1850_n2688# 0.754951f
C22 drain_right.t13 a_n1850_n2688# 0.239925f
C23 drain_right.t7 a_n1850_n2688# 0.239925f
C24 drain_right.n3 a_n1850_n2688# 2.10184f
C25 drain_right.t12 a_n1850_n2688# 0.239925f
C26 drain_right.t6 a_n1850_n2688# 0.239925f
C27 drain_right.n4 a_n1850_n2688# 2.09854f
C28 drain_right.n5 a_n1850_n2688# 0.754951f
C29 drain_right.n6 a_n1850_n2688# 1.35627f
C30 drain_right.t3 a_n1850_n2688# 0.239925f
C31 drain_right.t5 a_n1850_n2688# 0.239925f
C32 drain_right.n7 a_n1850_n2688# 2.10184f
C33 drain_right.t8 a_n1850_n2688# 0.239925f
C34 drain_right.t14 a_n1850_n2688# 0.239925f
C35 drain_right.n8 a_n1850_n2688# 2.09854f
C36 drain_right.n9 a_n1850_n2688# 0.786868f
C37 drain_right.t15 a_n1850_n2688# 0.239925f
C38 drain_right.t4 a_n1850_n2688# 0.239925f
C39 drain_right.n10 a_n1850_n2688# 2.09854f
C40 drain_right.n11 a_n1850_n2688# 0.388288f
C41 drain_right.t2 a_n1850_n2688# 0.239925f
C42 drain_right.t11 a_n1850_n2688# 0.239925f
C43 drain_right.n12 a_n1850_n2688# 2.09854f
C44 drain_right.n13 a_n1850_n2688# 0.669083f
C45 minus.n0 a_n1850_n2688# 0.050632f
C46 minus.t13 a_n1850_n2688# 0.393028f
C47 minus.t4 a_n1850_n2688# 0.387373f
C48 minus.t0 a_n1850_n2688# 0.387373f
C49 minus.n1 a_n1850_n2688# 0.16176f
C50 minus.n2 a_n1850_n2688# 0.050632f
C51 minus.t11 a_n1850_n2688# 0.387373f
C52 minus.t7 a_n1850_n2688# 0.387373f
C53 minus.t1 a_n1850_n2688# 0.387373f
C54 minus.n3 a_n1850_n2688# 0.16176f
C55 minus.n4 a_n1850_n2688# 0.107753f
C56 minus.t12 a_n1850_n2688# 0.387373f
C57 minus.t10 a_n1850_n2688# 0.393028f
C58 minus.n5 a_n1850_n2688# 0.177183f
C59 minus.n6 a_n1850_n2688# 0.16176f
C60 minus.n7 a_n1850_n2688# 0.019138f
C61 minus.n8 a_n1850_n2688# 0.018513f
C62 minus.n9 a_n1850_n2688# 0.050632f
C63 minus.n10 a_n1850_n2688# 0.050632f
C64 minus.n11 a_n1850_n2688# 0.020855f
C65 minus.n12 a_n1850_n2688# 0.16176f
C66 minus.n13 a_n1850_n2688# 0.020855f
C67 minus.n14 a_n1850_n2688# 0.16176f
C68 minus.n15 a_n1850_n2688# 0.020855f
C69 minus.n16 a_n1850_n2688# 0.050632f
C70 minus.n17 a_n1850_n2688# 0.050632f
C71 minus.n18 a_n1850_n2688# 0.018513f
C72 minus.n19 a_n1850_n2688# 0.019138f
C73 minus.n20 a_n1850_n2688# 0.16176f
C74 minus.n21 a_n1850_n2688# 0.177116f
C75 minus.n22 a_n1850_n2688# 1.60554f
C76 minus.n23 a_n1850_n2688# 0.050632f
C77 minus.t2 a_n1850_n2688# 0.387373f
C78 minus.t9 a_n1850_n2688# 0.387373f
C79 minus.n24 a_n1850_n2688# 0.16176f
C80 minus.n25 a_n1850_n2688# 0.050632f
C81 minus.t3 a_n1850_n2688# 0.387373f
C82 minus.t5 a_n1850_n2688# 0.387373f
C83 minus.t14 a_n1850_n2688# 0.387373f
C84 minus.n26 a_n1850_n2688# 0.16176f
C85 minus.n27 a_n1850_n2688# 0.107753f
C86 minus.t6 a_n1850_n2688# 0.387373f
C87 minus.t15 a_n1850_n2688# 0.393028f
C88 minus.n28 a_n1850_n2688# 0.177183f
C89 minus.n29 a_n1850_n2688# 0.16176f
C90 minus.n30 a_n1850_n2688# 0.019138f
C91 minus.n31 a_n1850_n2688# 0.018513f
C92 minus.n32 a_n1850_n2688# 0.050632f
C93 minus.n33 a_n1850_n2688# 0.050632f
C94 minus.n34 a_n1850_n2688# 0.020855f
C95 minus.n35 a_n1850_n2688# 0.16176f
C96 minus.n36 a_n1850_n2688# 0.020855f
C97 minus.n37 a_n1850_n2688# 0.16176f
C98 minus.n38 a_n1850_n2688# 0.020855f
C99 minus.n39 a_n1850_n2688# 0.050632f
C100 minus.n40 a_n1850_n2688# 0.050632f
C101 minus.n41 a_n1850_n2688# 0.018513f
C102 minus.n42 a_n1850_n2688# 0.019138f
C103 minus.n43 a_n1850_n2688# 0.16176f
C104 minus.t8 a_n1850_n2688# 0.393028f
C105 minus.n44 a_n1850_n2688# 0.177116f
C106 minus.n45 a_n1850_n2688# 0.327006f
C107 minus.n46 a_n1850_n2688# 1.96508f
C108 drain_left.t6 a_n1850_n2688# 0.239654f
C109 drain_left.t13 a_n1850_n2688# 0.239654f
C110 drain_left.n0 a_n1850_n2688# 2.09947f
C111 drain_left.t8 a_n1850_n2688# 0.239654f
C112 drain_left.t14 a_n1850_n2688# 0.239654f
C113 drain_left.n1 a_n1850_n2688# 2.09617f
C114 drain_left.n2 a_n1850_n2688# 0.754099f
C115 drain_left.t11 a_n1850_n2688# 0.239654f
C116 drain_left.t4 a_n1850_n2688# 0.239654f
C117 drain_left.n3 a_n1850_n2688# 2.09947f
C118 drain_left.t9 a_n1850_n2688# 0.239654f
C119 drain_left.t2 a_n1850_n2688# 0.239654f
C120 drain_left.n4 a_n1850_n2688# 2.09617f
C121 drain_left.n5 a_n1850_n2688# 0.754099f
C122 drain_left.n6 a_n1850_n2688# 1.42409f
C123 drain_left.t12 a_n1850_n2688# 0.239654f
C124 drain_left.t7 a_n1850_n2688# 0.239654f
C125 drain_left.n7 a_n1850_n2688# 2.09947f
C126 drain_left.t3 a_n1850_n2688# 0.239654f
C127 drain_left.t0 a_n1850_n2688# 0.239654f
C128 drain_left.n8 a_n1850_n2688# 2.09617f
C129 drain_left.n9 a_n1850_n2688# 0.785972f
C130 drain_left.t10 a_n1850_n2688# 0.239654f
C131 drain_left.t5 a_n1850_n2688# 0.239654f
C132 drain_left.n10 a_n1850_n2688# 2.09617f
C133 drain_left.n11 a_n1850_n2688# 0.387849f
C134 drain_left.t1 a_n1850_n2688# 0.239654f
C135 drain_left.t15 a_n1850_n2688# 0.239654f
C136 drain_left.n12 a_n1850_n2688# 2.09617f
C137 drain_left.n13 a_n1850_n2688# 0.668337f
C138 source.t19 a_n1850_n2688# 2.18538f
C139 source.n0 a_n1850_n2688# 1.25665f
C140 source.t20 a_n1850_n2688# 0.204941f
C141 source.t25 a_n1850_n2688# 0.204941f
C142 source.n1 a_n1850_n2688# 1.71563f
C143 source.n2 a_n1850_n2688# 0.369426f
C144 source.t30 a_n1850_n2688# 0.204941f
C145 source.t29 a_n1850_n2688# 0.204941f
C146 source.n3 a_n1850_n2688# 1.71563f
C147 source.n4 a_n1850_n2688# 0.369426f
C148 source.t26 a_n1850_n2688# 0.204941f
C149 source.t24 a_n1850_n2688# 0.204941f
C150 source.n5 a_n1850_n2688# 1.71563f
C151 source.n6 a_n1850_n2688# 0.369426f
C152 source.t31 a_n1850_n2688# 2.18539f
C153 source.n7 a_n1850_n2688# 0.451798f
C154 source.t2 a_n1850_n2688# 2.18539f
C155 source.n8 a_n1850_n2688# 0.451798f
C156 source.t8 a_n1850_n2688# 0.204941f
C157 source.t9 a_n1850_n2688# 0.204941f
C158 source.n9 a_n1850_n2688# 1.71563f
C159 source.n10 a_n1850_n2688# 0.369426f
C160 source.t4 a_n1850_n2688# 0.204941f
C161 source.t13 a_n1850_n2688# 0.204941f
C162 source.n11 a_n1850_n2688# 1.71563f
C163 source.n12 a_n1850_n2688# 0.369426f
C164 source.t7 a_n1850_n2688# 0.204941f
C165 source.t1 a_n1850_n2688# 0.204941f
C166 source.n13 a_n1850_n2688# 1.71563f
C167 source.n14 a_n1850_n2688# 0.369426f
C168 source.t5 a_n1850_n2688# 2.18539f
C169 source.n15 a_n1850_n2688# 1.67535f
C170 source.t16 a_n1850_n2688# 2.18538f
C171 source.n16 a_n1850_n2688# 1.67535f
C172 source.t21 a_n1850_n2688# 0.204941f
C173 source.t27 a_n1850_n2688# 0.204941f
C174 source.n17 a_n1850_n2688# 1.71563f
C175 source.n18 a_n1850_n2688# 0.369431f
C176 source.t22 a_n1850_n2688# 0.204941f
C177 source.t28 a_n1850_n2688# 0.204941f
C178 source.n19 a_n1850_n2688# 1.71563f
C179 source.n20 a_n1850_n2688# 0.369431f
C180 source.t17 a_n1850_n2688# 0.204941f
C181 source.t18 a_n1850_n2688# 0.204941f
C182 source.n21 a_n1850_n2688# 1.71563f
C183 source.n22 a_n1850_n2688# 0.369431f
C184 source.t23 a_n1850_n2688# 2.18538f
C185 source.n23 a_n1850_n2688# 0.451803f
C186 source.t15 a_n1850_n2688# 2.18538f
C187 source.n24 a_n1850_n2688# 0.451803f
C188 source.t10 a_n1850_n2688# 0.204941f
C189 source.t14 a_n1850_n2688# 0.204941f
C190 source.n25 a_n1850_n2688# 1.71563f
C191 source.n26 a_n1850_n2688# 0.369431f
C192 source.t12 a_n1850_n2688# 0.204941f
C193 source.t6 a_n1850_n2688# 0.204941f
C194 source.n27 a_n1850_n2688# 1.71563f
C195 source.n28 a_n1850_n2688# 0.369431f
C196 source.t0 a_n1850_n2688# 0.204941f
C197 source.t11 a_n1850_n2688# 0.204941f
C198 source.n29 a_n1850_n2688# 1.71563f
C199 source.n30 a_n1850_n2688# 0.369431f
C200 source.t3 a_n1850_n2688# 2.18538f
C201 source.n31 a_n1850_n2688# 0.614469f
C202 source.n32 a_n1850_n2688# 1.50007f
C203 plus.n0 a_n1850_n2688# 0.051375f
C204 plus.t14 a_n1850_n2688# 0.393055f
C205 plus.t10 a_n1850_n2688# 0.393055f
C206 plus.n1 a_n1850_n2688# 0.164133f
C207 plus.n2 a_n1850_n2688# 0.051375f
C208 plus.t5 a_n1850_n2688# 0.393055f
C209 plus.t15 a_n1850_n2688# 0.393055f
C210 plus.t12 a_n1850_n2688# 0.393055f
C211 plus.n3 a_n1850_n2688# 0.164133f
C212 plus.n4 a_n1850_n2688# 0.109333f
C213 plus.t8 a_n1850_n2688# 0.393055f
C214 plus.t3 a_n1850_n2688# 0.398793f
C215 plus.n5 a_n1850_n2688# 0.179782f
C216 plus.n6 a_n1850_n2688# 0.164133f
C217 plus.n7 a_n1850_n2688# 0.019418f
C218 plus.n8 a_n1850_n2688# 0.018785f
C219 plus.n9 a_n1850_n2688# 0.051375f
C220 plus.n10 a_n1850_n2688# 0.051375f
C221 plus.n11 a_n1850_n2688# 0.02116f
C222 plus.n12 a_n1850_n2688# 0.164133f
C223 plus.n13 a_n1850_n2688# 0.02116f
C224 plus.n14 a_n1850_n2688# 0.164133f
C225 plus.n15 a_n1850_n2688# 0.02116f
C226 plus.n16 a_n1850_n2688# 0.051375f
C227 plus.n17 a_n1850_n2688# 0.051375f
C228 plus.n18 a_n1850_n2688# 0.018785f
C229 plus.n19 a_n1850_n2688# 0.019418f
C230 plus.n20 a_n1850_n2688# 0.164133f
C231 plus.t0 a_n1850_n2688# 0.398793f
C232 plus.n21 a_n1850_n2688# 0.179714f
C233 plus.n22 a_n1850_n2688# 0.500463f
C234 plus.n23 a_n1850_n2688# 0.051375f
C235 plus.t9 a_n1850_n2688# 0.398793f
C236 plus.t2 a_n1850_n2688# 0.393055f
C237 plus.t7 a_n1850_n2688# 0.393055f
C238 plus.n24 a_n1850_n2688# 0.164133f
C239 plus.n25 a_n1850_n2688# 0.051375f
C240 plus.t1 a_n1850_n2688# 0.393055f
C241 plus.t6 a_n1850_n2688# 0.393055f
C242 plus.t13 a_n1850_n2688# 0.393055f
C243 plus.n26 a_n1850_n2688# 0.164133f
C244 plus.n27 a_n1850_n2688# 0.109333f
C245 plus.t4 a_n1850_n2688# 0.393055f
C246 plus.t11 a_n1850_n2688# 0.398793f
C247 plus.n28 a_n1850_n2688# 0.179782f
C248 plus.n29 a_n1850_n2688# 0.164133f
C249 plus.n30 a_n1850_n2688# 0.019418f
C250 plus.n31 a_n1850_n2688# 0.018785f
C251 plus.n32 a_n1850_n2688# 0.051375f
C252 plus.n33 a_n1850_n2688# 0.051375f
C253 plus.n34 a_n1850_n2688# 0.02116f
C254 plus.n35 a_n1850_n2688# 0.164133f
C255 plus.n36 a_n1850_n2688# 0.02116f
C256 plus.n37 a_n1850_n2688# 0.164133f
C257 plus.n38 a_n1850_n2688# 0.02116f
C258 plus.n39 a_n1850_n2688# 0.051375f
C259 plus.n40 a_n1850_n2688# 0.051375f
C260 plus.n41 a_n1850_n2688# 0.018785f
C261 plus.n42 a_n1850_n2688# 0.019418f
C262 plus.n43 a_n1850_n2688# 0.164133f
C263 plus.n44 a_n1850_n2688# 0.179714f
C264 plus.n45 a_n1850_n2688# 1.42029f
.ends

