* NGSPICE file created from diffpair447.ext - technology: sky130A

.subckt diffpair447 minus drain_right drain_left source plus
X0 source.t31 plus.t0 drain_left.t10 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X1 drain_left.t15 plus.t1 source.t30 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X2 drain_right.t15 minus.t0 source.t2 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X3 drain_right.t14 minus.t1 source.t9 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X4 source.t6 minus.t2 drain_right.t13 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.5
X5 source.t7 minus.t3 drain_right.t12 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X6 source.t29 plus.t2 drain_left.t12 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.5
X7 source.t10 minus.t4 drain_right.t11 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X8 drain_left.t4 plus.t3 source.t28 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X9 drain_right.t10 minus.t5 source.t5 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X10 a_n2210_n3288# a_n2210_n3288# a_n2210_n3288# a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.5
X11 drain_left.t13 plus.t4 source.t27 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X12 drain_right.t9 minus.t6 source.t14 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X13 drain_right.t8 minus.t7 source.t15 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.5
X14 drain_left.t14 plus.t5 source.t26 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X15 source.t25 plus.t6 drain_left.t11 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X16 drain_right.t7 minus.t8 source.t3 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X17 source.t11 minus.t9 drain_right.t6 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X18 source.t24 plus.t7 drain_left.t5 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X19 source.t4 minus.t10 drain_right.t5 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X20 source.t8 minus.t11 drain_right.t4 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.5
X21 a_n2210_n3288# a_n2210_n3288# a_n2210_n3288# a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.5
X22 source.t12 minus.t12 drain_right.t3 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X23 drain_right.t2 minus.t13 source.t0 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X24 drain_right.t1 minus.t14 source.t13 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.5
X25 a_n2210_n3288# a_n2210_n3288# a_n2210_n3288# a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.5
X26 drain_left.t9 plus.t8 source.t23 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X27 source.t1 minus.t15 drain_right.t0 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X28 source.t22 plus.t9 drain_left.t8 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X29 drain_left.t0 plus.t10 source.t21 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.5
X30 source.t20 plus.t11 drain_left.t1 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X31 drain_left.t6 plus.t12 source.t19 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.5
X32 source.t18 plus.t13 drain_left.t2 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
X33 a_n2210_n3288# a_n2210_n3288# a_n2210_n3288# a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.5
X34 source.t17 plus.t14 drain_left.t7 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.5
X35 drain_left.t3 plus.t15 source.t16 a_n2210_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.5
R0 plus.n5 plus.t2 677.948
R1 plus.n27 plus.t10 677.948
R2 plus.n20 plus.t12 656.966
R3 plus.n19 plus.t7 656.966
R4 plus.n1 plus.t15 656.966
R5 plus.n13 plus.t9 656.966
R6 plus.n12 plus.t5 656.966
R7 plus.n4 plus.t13 656.966
R8 plus.n6 plus.t8 656.966
R9 plus.n42 plus.t14 656.966
R10 plus.n41 plus.t3 656.966
R11 plus.n23 plus.t6 656.966
R12 plus.n35 plus.t1 656.966
R13 plus.n34 plus.t0 656.966
R14 plus.n26 plus.t4 656.966
R15 plus.n28 plus.t11 656.966
R16 plus.n8 plus.n7 161.3
R17 plus.n9 plus.n4 161.3
R18 plus.n11 plus.n10 161.3
R19 plus.n12 plus.n3 161.3
R20 plus.n13 plus.n2 161.3
R21 plus.n15 plus.n14 161.3
R22 plus.n16 plus.n1 161.3
R23 plus.n18 plus.n17 161.3
R24 plus.n19 plus.n0 161.3
R25 plus.n21 plus.n20 161.3
R26 plus.n30 plus.n29 161.3
R27 plus.n31 plus.n26 161.3
R28 plus.n33 plus.n32 161.3
R29 plus.n34 plus.n25 161.3
R30 plus.n35 plus.n24 161.3
R31 plus.n37 plus.n36 161.3
R32 plus.n38 plus.n23 161.3
R33 plus.n40 plus.n39 161.3
R34 plus.n41 plus.n22 161.3
R35 plus.n43 plus.n42 161.3
R36 plus.n8 plus.n5 70.4033
R37 plus.n30 plus.n27 70.4033
R38 plus.n20 plus.n19 48.2005
R39 plus.n13 plus.n12 48.2005
R40 plus.n42 plus.n41 48.2005
R41 plus.n35 plus.n34 48.2005
R42 plus.n18 plus.n1 37.246
R43 plus.n7 plus.n4 37.246
R44 plus.n40 plus.n23 37.246
R45 plus.n29 plus.n26 37.246
R46 plus.n14 plus.n1 35.7853
R47 plus.n11 plus.n4 35.7853
R48 plus.n36 plus.n23 35.7853
R49 plus.n33 plus.n26 35.7853
R50 plus plus.n43 31.4346
R51 plus.n6 plus.n5 20.9576
R52 plus.n28 plus.n27 20.9576
R53 plus.n14 plus.n13 12.4157
R54 plus.n12 plus.n11 12.4157
R55 plus.n36 plus.n35 12.4157
R56 plus.n34 plus.n33 12.4157
R57 plus plus.n21 12.205
R58 plus.n19 plus.n18 10.955
R59 plus.n7 plus.n6 10.955
R60 plus.n41 plus.n40 10.955
R61 plus.n29 plus.n28 10.955
R62 plus.n9 plus.n8 0.189894
R63 plus.n10 plus.n9 0.189894
R64 plus.n10 plus.n3 0.189894
R65 plus.n3 plus.n2 0.189894
R66 plus.n15 plus.n2 0.189894
R67 plus.n16 plus.n15 0.189894
R68 plus.n17 plus.n16 0.189894
R69 plus.n17 plus.n0 0.189894
R70 plus.n21 plus.n0 0.189894
R71 plus.n43 plus.n22 0.189894
R72 plus.n39 plus.n22 0.189894
R73 plus.n39 plus.n38 0.189894
R74 plus.n38 plus.n37 0.189894
R75 plus.n37 plus.n24 0.189894
R76 plus.n25 plus.n24 0.189894
R77 plus.n32 plus.n25 0.189894
R78 plus.n32 plus.n31 0.189894
R79 plus.n31 plus.n30 0.189894
R80 drain_left.n9 drain_left.n7 60.2682
R81 drain_left.n5 drain_left.n3 60.268
R82 drain_left.n2 drain_left.n0 60.268
R83 drain_left.n11 drain_left.n10 59.5527
R84 drain_left.n9 drain_left.n8 59.5527
R85 drain_left.n5 drain_left.n4 59.5525
R86 drain_left.n2 drain_left.n1 59.5525
R87 drain_left.n13 drain_left.n12 59.5525
R88 drain_left drain_left.n6 32.0179
R89 drain_left drain_left.n13 6.36873
R90 drain_left.n3 drain_left.t1 1.6505
R91 drain_left.n3 drain_left.t0 1.6505
R92 drain_left.n4 drain_left.t10 1.6505
R93 drain_left.n4 drain_left.t13 1.6505
R94 drain_left.n1 drain_left.t11 1.6505
R95 drain_left.n1 drain_left.t15 1.6505
R96 drain_left.n0 drain_left.t7 1.6505
R97 drain_left.n0 drain_left.t4 1.6505
R98 drain_left.n12 drain_left.t5 1.6505
R99 drain_left.n12 drain_left.t6 1.6505
R100 drain_left.n10 drain_left.t8 1.6505
R101 drain_left.n10 drain_left.t3 1.6505
R102 drain_left.n8 drain_left.t2 1.6505
R103 drain_left.n8 drain_left.t14 1.6505
R104 drain_left.n7 drain_left.t12 1.6505
R105 drain_left.n7 drain_left.t9 1.6505
R106 drain_left.n11 drain_left.n9 0.716017
R107 drain_left.n13 drain_left.n11 0.716017
R108 drain_left.n6 drain_left.n5 0.302913
R109 drain_left.n6 drain_left.n2 0.302913
R110 source.n546 source.n486 289.615
R111 source.n474 source.n414 289.615
R112 source.n408 source.n348 289.615
R113 source.n336 source.n276 289.615
R114 source.n60 source.n0 289.615
R115 source.n132 source.n72 289.615
R116 source.n198 source.n138 289.615
R117 source.n270 source.n210 289.615
R118 source.n506 source.n505 185
R119 source.n511 source.n510 185
R120 source.n513 source.n512 185
R121 source.n502 source.n501 185
R122 source.n519 source.n518 185
R123 source.n521 source.n520 185
R124 source.n498 source.n497 185
R125 source.n528 source.n527 185
R126 source.n529 source.n496 185
R127 source.n531 source.n530 185
R128 source.n494 source.n493 185
R129 source.n537 source.n536 185
R130 source.n539 source.n538 185
R131 source.n490 source.n489 185
R132 source.n545 source.n544 185
R133 source.n547 source.n546 185
R134 source.n434 source.n433 185
R135 source.n439 source.n438 185
R136 source.n441 source.n440 185
R137 source.n430 source.n429 185
R138 source.n447 source.n446 185
R139 source.n449 source.n448 185
R140 source.n426 source.n425 185
R141 source.n456 source.n455 185
R142 source.n457 source.n424 185
R143 source.n459 source.n458 185
R144 source.n422 source.n421 185
R145 source.n465 source.n464 185
R146 source.n467 source.n466 185
R147 source.n418 source.n417 185
R148 source.n473 source.n472 185
R149 source.n475 source.n474 185
R150 source.n368 source.n367 185
R151 source.n373 source.n372 185
R152 source.n375 source.n374 185
R153 source.n364 source.n363 185
R154 source.n381 source.n380 185
R155 source.n383 source.n382 185
R156 source.n360 source.n359 185
R157 source.n390 source.n389 185
R158 source.n391 source.n358 185
R159 source.n393 source.n392 185
R160 source.n356 source.n355 185
R161 source.n399 source.n398 185
R162 source.n401 source.n400 185
R163 source.n352 source.n351 185
R164 source.n407 source.n406 185
R165 source.n409 source.n408 185
R166 source.n296 source.n295 185
R167 source.n301 source.n300 185
R168 source.n303 source.n302 185
R169 source.n292 source.n291 185
R170 source.n309 source.n308 185
R171 source.n311 source.n310 185
R172 source.n288 source.n287 185
R173 source.n318 source.n317 185
R174 source.n319 source.n286 185
R175 source.n321 source.n320 185
R176 source.n284 source.n283 185
R177 source.n327 source.n326 185
R178 source.n329 source.n328 185
R179 source.n280 source.n279 185
R180 source.n335 source.n334 185
R181 source.n337 source.n336 185
R182 source.n61 source.n60 185
R183 source.n59 source.n58 185
R184 source.n4 source.n3 185
R185 source.n53 source.n52 185
R186 source.n51 source.n50 185
R187 source.n8 source.n7 185
R188 source.n45 source.n44 185
R189 source.n43 source.n10 185
R190 source.n42 source.n41 185
R191 source.n13 source.n11 185
R192 source.n36 source.n35 185
R193 source.n34 source.n33 185
R194 source.n17 source.n16 185
R195 source.n28 source.n27 185
R196 source.n26 source.n25 185
R197 source.n21 source.n20 185
R198 source.n133 source.n132 185
R199 source.n131 source.n130 185
R200 source.n76 source.n75 185
R201 source.n125 source.n124 185
R202 source.n123 source.n122 185
R203 source.n80 source.n79 185
R204 source.n117 source.n116 185
R205 source.n115 source.n82 185
R206 source.n114 source.n113 185
R207 source.n85 source.n83 185
R208 source.n108 source.n107 185
R209 source.n106 source.n105 185
R210 source.n89 source.n88 185
R211 source.n100 source.n99 185
R212 source.n98 source.n97 185
R213 source.n93 source.n92 185
R214 source.n199 source.n198 185
R215 source.n197 source.n196 185
R216 source.n142 source.n141 185
R217 source.n191 source.n190 185
R218 source.n189 source.n188 185
R219 source.n146 source.n145 185
R220 source.n183 source.n182 185
R221 source.n181 source.n148 185
R222 source.n180 source.n179 185
R223 source.n151 source.n149 185
R224 source.n174 source.n173 185
R225 source.n172 source.n171 185
R226 source.n155 source.n154 185
R227 source.n166 source.n165 185
R228 source.n164 source.n163 185
R229 source.n159 source.n158 185
R230 source.n271 source.n270 185
R231 source.n269 source.n268 185
R232 source.n214 source.n213 185
R233 source.n263 source.n262 185
R234 source.n261 source.n260 185
R235 source.n218 source.n217 185
R236 source.n255 source.n254 185
R237 source.n253 source.n220 185
R238 source.n252 source.n251 185
R239 source.n223 source.n221 185
R240 source.n246 source.n245 185
R241 source.n244 source.n243 185
R242 source.n227 source.n226 185
R243 source.n238 source.n237 185
R244 source.n236 source.n235 185
R245 source.n231 source.n230 185
R246 source.n507 source.t15 149.524
R247 source.n435 source.t6 149.524
R248 source.n369 source.t21 149.524
R249 source.n297 source.t17 149.524
R250 source.n22 source.t19 149.524
R251 source.n94 source.t29 149.524
R252 source.n160 source.t13 149.524
R253 source.n232 source.t8 149.524
R254 source.n511 source.n505 104.615
R255 source.n512 source.n511 104.615
R256 source.n512 source.n501 104.615
R257 source.n519 source.n501 104.615
R258 source.n520 source.n519 104.615
R259 source.n520 source.n497 104.615
R260 source.n528 source.n497 104.615
R261 source.n529 source.n528 104.615
R262 source.n530 source.n529 104.615
R263 source.n530 source.n493 104.615
R264 source.n537 source.n493 104.615
R265 source.n538 source.n537 104.615
R266 source.n538 source.n489 104.615
R267 source.n545 source.n489 104.615
R268 source.n546 source.n545 104.615
R269 source.n439 source.n433 104.615
R270 source.n440 source.n439 104.615
R271 source.n440 source.n429 104.615
R272 source.n447 source.n429 104.615
R273 source.n448 source.n447 104.615
R274 source.n448 source.n425 104.615
R275 source.n456 source.n425 104.615
R276 source.n457 source.n456 104.615
R277 source.n458 source.n457 104.615
R278 source.n458 source.n421 104.615
R279 source.n465 source.n421 104.615
R280 source.n466 source.n465 104.615
R281 source.n466 source.n417 104.615
R282 source.n473 source.n417 104.615
R283 source.n474 source.n473 104.615
R284 source.n373 source.n367 104.615
R285 source.n374 source.n373 104.615
R286 source.n374 source.n363 104.615
R287 source.n381 source.n363 104.615
R288 source.n382 source.n381 104.615
R289 source.n382 source.n359 104.615
R290 source.n390 source.n359 104.615
R291 source.n391 source.n390 104.615
R292 source.n392 source.n391 104.615
R293 source.n392 source.n355 104.615
R294 source.n399 source.n355 104.615
R295 source.n400 source.n399 104.615
R296 source.n400 source.n351 104.615
R297 source.n407 source.n351 104.615
R298 source.n408 source.n407 104.615
R299 source.n301 source.n295 104.615
R300 source.n302 source.n301 104.615
R301 source.n302 source.n291 104.615
R302 source.n309 source.n291 104.615
R303 source.n310 source.n309 104.615
R304 source.n310 source.n287 104.615
R305 source.n318 source.n287 104.615
R306 source.n319 source.n318 104.615
R307 source.n320 source.n319 104.615
R308 source.n320 source.n283 104.615
R309 source.n327 source.n283 104.615
R310 source.n328 source.n327 104.615
R311 source.n328 source.n279 104.615
R312 source.n335 source.n279 104.615
R313 source.n336 source.n335 104.615
R314 source.n60 source.n59 104.615
R315 source.n59 source.n3 104.615
R316 source.n52 source.n3 104.615
R317 source.n52 source.n51 104.615
R318 source.n51 source.n7 104.615
R319 source.n44 source.n7 104.615
R320 source.n44 source.n43 104.615
R321 source.n43 source.n42 104.615
R322 source.n42 source.n11 104.615
R323 source.n35 source.n11 104.615
R324 source.n35 source.n34 104.615
R325 source.n34 source.n16 104.615
R326 source.n27 source.n16 104.615
R327 source.n27 source.n26 104.615
R328 source.n26 source.n20 104.615
R329 source.n132 source.n131 104.615
R330 source.n131 source.n75 104.615
R331 source.n124 source.n75 104.615
R332 source.n124 source.n123 104.615
R333 source.n123 source.n79 104.615
R334 source.n116 source.n79 104.615
R335 source.n116 source.n115 104.615
R336 source.n115 source.n114 104.615
R337 source.n114 source.n83 104.615
R338 source.n107 source.n83 104.615
R339 source.n107 source.n106 104.615
R340 source.n106 source.n88 104.615
R341 source.n99 source.n88 104.615
R342 source.n99 source.n98 104.615
R343 source.n98 source.n92 104.615
R344 source.n198 source.n197 104.615
R345 source.n197 source.n141 104.615
R346 source.n190 source.n141 104.615
R347 source.n190 source.n189 104.615
R348 source.n189 source.n145 104.615
R349 source.n182 source.n145 104.615
R350 source.n182 source.n181 104.615
R351 source.n181 source.n180 104.615
R352 source.n180 source.n149 104.615
R353 source.n173 source.n149 104.615
R354 source.n173 source.n172 104.615
R355 source.n172 source.n154 104.615
R356 source.n165 source.n154 104.615
R357 source.n165 source.n164 104.615
R358 source.n164 source.n158 104.615
R359 source.n270 source.n269 104.615
R360 source.n269 source.n213 104.615
R361 source.n262 source.n213 104.615
R362 source.n262 source.n261 104.615
R363 source.n261 source.n217 104.615
R364 source.n254 source.n217 104.615
R365 source.n254 source.n253 104.615
R366 source.n253 source.n252 104.615
R367 source.n252 source.n221 104.615
R368 source.n245 source.n221 104.615
R369 source.n245 source.n244 104.615
R370 source.n244 source.n226 104.615
R371 source.n237 source.n226 104.615
R372 source.n237 source.n236 104.615
R373 source.n236 source.n230 104.615
R374 source.t15 source.n505 52.3082
R375 source.t6 source.n433 52.3082
R376 source.t21 source.n367 52.3082
R377 source.t17 source.n295 52.3082
R378 source.t19 source.n20 52.3082
R379 source.t29 source.n92 52.3082
R380 source.t13 source.n158 52.3082
R381 source.t8 source.n230 52.3082
R382 source.n67 source.n66 42.8739
R383 source.n69 source.n68 42.8739
R384 source.n71 source.n70 42.8739
R385 source.n205 source.n204 42.8739
R386 source.n207 source.n206 42.8739
R387 source.n209 source.n208 42.8739
R388 source.n485 source.n484 42.8737
R389 source.n483 source.n482 42.8737
R390 source.n481 source.n480 42.8737
R391 source.n347 source.n346 42.8737
R392 source.n345 source.n344 42.8737
R393 source.n343 source.n342 42.8737
R394 source.n551 source.n550 29.8581
R395 source.n479 source.n478 29.8581
R396 source.n413 source.n412 29.8581
R397 source.n341 source.n340 29.8581
R398 source.n65 source.n64 29.8581
R399 source.n137 source.n136 29.8581
R400 source.n203 source.n202 29.8581
R401 source.n275 source.n274 29.8581
R402 source.n341 source.n275 22.0032
R403 source.n552 source.n65 16.3826
R404 source.n531 source.n496 13.1884
R405 source.n459 source.n424 13.1884
R406 source.n393 source.n358 13.1884
R407 source.n321 source.n286 13.1884
R408 source.n45 source.n10 13.1884
R409 source.n117 source.n82 13.1884
R410 source.n183 source.n148 13.1884
R411 source.n255 source.n220 13.1884
R412 source.n527 source.n526 12.8005
R413 source.n532 source.n494 12.8005
R414 source.n455 source.n454 12.8005
R415 source.n460 source.n422 12.8005
R416 source.n389 source.n388 12.8005
R417 source.n394 source.n356 12.8005
R418 source.n317 source.n316 12.8005
R419 source.n322 source.n284 12.8005
R420 source.n46 source.n8 12.8005
R421 source.n41 source.n12 12.8005
R422 source.n118 source.n80 12.8005
R423 source.n113 source.n84 12.8005
R424 source.n184 source.n146 12.8005
R425 source.n179 source.n150 12.8005
R426 source.n256 source.n218 12.8005
R427 source.n251 source.n222 12.8005
R428 source.n525 source.n498 12.0247
R429 source.n536 source.n535 12.0247
R430 source.n453 source.n426 12.0247
R431 source.n464 source.n463 12.0247
R432 source.n387 source.n360 12.0247
R433 source.n398 source.n397 12.0247
R434 source.n315 source.n288 12.0247
R435 source.n326 source.n325 12.0247
R436 source.n50 source.n49 12.0247
R437 source.n40 source.n13 12.0247
R438 source.n122 source.n121 12.0247
R439 source.n112 source.n85 12.0247
R440 source.n188 source.n187 12.0247
R441 source.n178 source.n151 12.0247
R442 source.n260 source.n259 12.0247
R443 source.n250 source.n223 12.0247
R444 source.n522 source.n521 11.249
R445 source.n539 source.n492 11.249
R446 source.n450 source.n449 11.249
R447 source.n467 source.n420 11.249
R448 source.n384 source.n383 11.249
R449 source.n401 source.n354 11.249
R450 source.n312 source.n311 11.249
R451 source.n329 source.n282 11.249
R452 source.n53 source.n6 11.249
R453 source.n37 source.n36 11.249
R454 source.n125 source.n78 11.249
R455 source.n109 source.n108 11.249
R456 source.n191 source.n144 11.249
R457 source.n175 source.n174 11.249
R458 source.n263 source.n216 11.249
R459 source.n247 source.n246 11.249
R460 source.n518 source.n500 10.4732
R461 source.n540 source.n490 10.4732
R462 source.n446 source.n428 10.4732
R463 source.n468 source.n418 10.4732
R464 source.n380 source.n362 10.4732
R465 source.n402 source.n352 10.4732
R466 source.n308 source.n290 10.4732
R467 source.n330 source.n280 10.4732
R468 source.n54 source.n4 10.4732
R469 source.n33 source.n15 10.4732
R470 source.n126 source.n76 10.4732
R471 source.n105 source.n87 10.4732
R472 source.n192 source.n142 10.4732
R473 source.n171 source.n153 10.4732
R474 source.n264 source.n214 10.4732
R475 source.n243 source.n225 10.4732
R476 source.n507 source.n506 10.2747
R477 source.n435 source.n434 10.2747
R478 source.n369 source.n368 10.2747
R479 source.n297 source.n296 10.2747
R480 source.n22 source.n21 10.2747
R481 source.n94 source.n93 10.2747
R482 source.n160 source.n159 10.2747
R483 source.n232 source.n231 10.2747
R484 source.n517 source.n502 9.69747
R485 source.n544 source.n543 9.69747
R486 source.n445 source.n430 9.69747
R487 source.n472 source.n471 9.69747
R488 source.n379 source.n364 9.69747
R489 source.n406 source.n405 9.69747
R490 source.n307 source.n292 9.69747
R491 source.n334 source.n333 9.69747
R492 source.n58 source.n57 9.69747
R493 source.n32 source.n17 9.69747
R494 source.n130 source.n129 9.69747
R495 source.n104 source.n89 9.69747
R496 source.n196 source.n195 9.69747
R497 source.n170 source.n155 9.69747
R498 source.n268 source.n267 9.69747
R499 source.n242 source.n227 9.69747
R500 source.n550 source.n549 9.45567
R501 source.n478 source.n477 9.45567
R502 source.n412 source.n411 9.45567
R503 source.n340 source.n339 9.45567
R504 source.n64 source.n63 9.45567
R505 source.n136 source.n135 9.45567
R506 source.n202 source.n201 9.45567
R507 source.n274 source.n273 9.45567
R508 source.n549 source.n548 9.3005
R509 source.n488 source.n487 9.3005
R510 source.n543 source.n542 9.3005
R511 source.n541 source.n540 9.3005
R512 source.n492 source.n491 9.3005
R513 source.n535 source.n534 9.3005
R514 source.n533 source.n532 9.3005
R515 source.n509 source.n508 9.3005
R516 source.n504 source.n503 9.3005
R517 source.n515 source.n514 9.3005
R518 source.n517 source.n516 9.3005
R519 source.n500 source.n499 9.3005
R520 source.n523 source.n522 9.3005
R521 source.n525 source.n524 9.3005
R522 source.n526 source.n495 9.3005
R523 source.n477 source.n476 9.3005
R524 source.n416 source.n415 9.3005
R525 source.n471 source.n470 9.3005
R526 source.n469 source.n468 9.3005
R527 source.n420 source.n419 9.3005
R528 source.n463 source.n462 9.3005
R529 source.n461 source.n460 9.3005
R530 source.n437 source.n436 9.3005
R531 source.n432 source.n431 9.3005
R532 source.n443 source.n442 9.3005
R533 source.n445 source.n444 9.3005
R534 source.n428 source.n427 9.3005
R535 source.n451 source.n450 9.3005
R536 source.n453 source.n452 9.3005
R537 source.n454 source.n423 9.3005
R538 source.n411 source.n410 9.3005
R539 source.n350 source.n349 9.3005
R540 source.n405 source.n404 9.3005
R541 source.n403 source.n402 9.3005
R542 source.n354 source.n353 9.3005
R543 source.n397 source.n396 9.3005
R544 source.n395 source.n394 9.3005
R545 source.n371 source.n370 9.3005
R546 source.n366 source.n365 9.3005
R547 source.n377 source.n376 9.3005
R548 source.n379 source.n378 9.3005
R549 source.n362 source.n361 9.3005
R550 source.n385 source.n384 9.3005
R551 source.n387 source.n386 9.3005
R552 source.n388 source.n357 9.3005
R553 source.n339 source.n338 9.3005
R554 source.n278 source.n277 9.3005
R555 source.n333 source.n332 9.3005
R556 source.n331 source.n330 9.3005
R557 source.n282 source.n281 9.3005
R558 source.n325 source.n324 9.3005
R559 source.n323 source.n322 9.3005
R560 source.n299 source.n298 9.3005
R561 source.n294 source.n293 9.3005
R562 source.n305 source.n304 9.3005
R563 source.n307 source.n306 9.3005
R564 source.n290 source.n289 9.3005
R565 source.n313 source.n312 9.3005
R566 source.n315 source.n314 9.3005
R567 source.n316 source.n285 9.3005
R568 source.n24 source.n23 9.3005
R569 source.n19 source.n18 9.3005
R570 source.n30 source.n29 9.3005
R571 source.n32 source.n31 9.3005
R572 source.n15 source.n14 9.3005
R573 source.n38 source.n37 9.3005
R574 source.n40 source.n39 9.3005
R575 source.n12 source.n9 9.3005
R576 source.n63 source.n62 9.3005
R577 source.n2 source.n1 9.3005
R578 source.n57 source.n56 9.3005
R579 source.n55 source.n54 9.3005
R580 source.n6 source.n5 9.3005
R581 source.n49 source.n48 9.3005
R582 source.n47 source.n46 9.3005
R583 source.n96 source.n95 9.3005
R584 source.n91 source.n90 9.3005
R585 source.n102 source.n101 9.3005
R586 source.n104 source.n103 9.3005
R587 source.n87 source.n86 9.3005
R588 source.n110 source.n109 9.3005
R589 source.n112 source.n111 9.3005
R590 source.n84 source.n81 9.3005
R591 source.n135 source.n134 9.3005
R592 source.n74 source.n73 9.3005
R593 source.n129 source.n128 9.3005
R594 source.n127 source.n126 9.3005
R595 source.n78 source.n77 9.3005
R596 source.n121 source.n120 9.3005
R597 source.n119 source.n118 9.3005
R598 source.n162 source.n161 9.3005
R599 source.n157 source.n156 9.3005
R600 source.n168 source.n167 9.3005
R601 source.n170 source.n169 9.3005
R602 source.n153 source.n152 9.3005
R603 source.n176 source.n175 9.3005
R604 source.n178 source.n177 9.3005
R605 source.n150 source.n147 9.3005
R606 source.n201 source.n200 9.3005
R607 source.n140 source.n139 9.3005
R608 source.n195 source.n194 9.3005
R609 source.n193 source.n192 9.3005
R610 source.n144 source.n143 9.3005
R611 source.n187 source.n186 9.3005
R612 source.n185 source.n184 9.3005
R613 source.n234 source.n233 9.3005
R614 source.n229 source.n228 9.3005
R615 source.n240 source.n239 9.3005
R616 source.n242 source.n241 9.3005
R617 source.n225 source.n224 9.3005
R618 source.n248 source.n247 9.3005
R619 source.n250 source.n249 9.3005
R620 source.n222 source.n219 9.3005
R621 source.n273 source.n272 9.3005
R622 source.n212 source.n211 9.3005
R623 source.n267 source.n266 9.3005
R624 source.n265 source.n264 9.3005
R625 source.n216 source.n215 9.3005
R626 source.n259 source.n258 9.3005
R627 source.n257 source.n256 9.3005
R628 source.n514 source.n513 8.92171
R629 source.n547 source.n488 8.92171
R630 source.n442 source.n441 8.92171
R631 source.n475 source.n416 8.92171
R632 source.n376 source.n375 8.92171
R633 source.n409 source.n350 8.92171
R634 source.n304 source.n303 8.92171
R635 source.n337 source.n278 8.92171
R636 source.n61 source.n2 8.92171
R637 source.n29 source.n28 8.92171
R638 source.n133 source.n74 8.92171
R639 source.n101 source.n100 8.92171
R640 source.n199 source.n140 8.92171
R641 source.n167 source.n166 8.92171
R642 source.n271 source.n212 8.92171
R643 source.n239 source.n238 8.92171
R644 source.n510 source.n504 8.14595
R645 source.n548 source.n486 8.14595
R646 source.n438 source.n432 8.14595
R647 source.n476 source.n414 8.14595
R648 source.n372 source.n366 8.14595
R649 source.n410 source.n348 8.14595
R650 source.n300 source.n294 8.14595
R651 source.n338 source.n276 8.14595
R652 source.n62 source.n0 8.14595
R653 source.n25 source.n19 8.14595
R654 source.n134 source.n72 8.14595
R655 source.n97 source.n91 8.14595
R656 source.n200 source.n138 8.14595
R657 source.n163 source.n157 8.14595
R658 source.n272 source.n210 8.14595
R659 source.n235 source.n229 8.14595
R660 source.n509 source.n506 7.3702
R661 source.n437 source.n434 7.3702
R662 source.n371 source.n368 7.3702
R663 source.n299 source.n296 7.3702
R664 source.n24 source.n21 7.3702
R665 source.n96 source.n93 7.3702
R666 source.n162 source.n159 7.3702
R667 source.n234 source.n231 7.3702
R668 source.n510 source.n509 5.81868
R669 source.n550 source.n486 5.81868
R670 source.n438 source.n437 5.81868
R671 source.n478 source.n414 5.81868
R672 source.n372 source.n371 5.81868
R673 source.n412 source.n348 5.81868
R674 source.n300 source.n299 5.81868
R675 source.n340 source.n276 5.81868
R676 source.n64 source.n0 5.81868
R677 source.n25 source.n24 5.81868
R678 source.n136 source.n72 5.81868
R679 source.n97 source.n96 5.81868
R680 source.n202 source.n138 5.81868
R681 source.n163 source.n162 5.81868
R682 source.n274 source.n210 5.81868
R683 source.n235 source.n234 5.81868
R684 source.n552 source.n551 5.62119
R685 source.n513 source.n504 5.04292
R686 source.n548 source.n547 5.04292
R687 source.n441 source.n432 5.04292
R688 source.n476 source.n475 5.04292
R689 source.n375 source.n366 5.04292
R690 source.n410 source.n409 5.04292
R691 source.n303 source.n294 5.04292
R692 source.n338 source.n337 5.04292
R693 source.n62 source.n61 5.04292
R694 source.n28 source.n19 5.04292
R695 source.n134 source.n133 5.04292
R696 source.n100 source.n91 5.04292
R697 source.n200 source.n199 5.04292
R698 source.n166 source.n157 5.04292
R699 source.n272 source.n271 5.04292
R700 source.n238 source.n229 5.04292
R701 source.n514 source.n502 4.26717
R702 source.n544 source.n488 4.26717
R703 source.n442 source.n430 4.26717
R704 source.n472 source.n416 4.26717
R705 source.n376 source.n364 4.26717
R706 source.n406 source.n350 4.26717
R707 source.n304 source.n292 4.26717
R708 source.n334 source.n278 4.26717
R709 source.n58 source.n2 4.26717
R710 source.n29 source.n17 4.26717
R711 source.n130 source.n74 4.26717
R712 source.n101 source.n89 4.26717
R713 source.n196 source.n140 4.26717
R714 source.n167 source.n155 4.26717
R715 source.n268 source.n212 4.26717
R716 source.n239 source.n227 4.26717
R717 source.n518 source.n517 3.49141
R718 source.n543 source.n490 3.49141
R719 source.n446 source.n445 3.49141
R720 source.n471 source.n418 3.49141
R721 source.n380 source.n379 3.49141
R722 source.n405 source.n352 3.49141
R723 source.n308 source.n307 3.49141
R724 source.n333 source.n280 3.49141
R725 source.n57 source.n4 3.49141
R726 source.n33 source.n32 3.49141
R727 source.n129 source.n76 3.49141
R728 source.n105 source.n104 3.49141
R729 source.n195 source.n142 3.49141
R730 source.n171 source.n170 3.49141
R731 source.n267 source.n214 3.49141
R732 source.n243 source.n242 3.49141
R733 source.n508 source.n507 2.84303
R734 source.n436 source.n435 2.84303
R735 source.n370 source.n369 2.84303
R736 source.n298 source.n297 2.84303
R737 source.n23 source.n22 2.84303
R738 source.n95 source.n94 2.84303
R739 source.n161 source.n160 2.84303
R740 source.n233 source.n232 2.84303
R741 source.n521 source.n500 2.71565
R742 source.n540 source.n539 2.71565
R743 source.n449 source.n428 2.71565
R744 source.n468 source.n467 2.71565
R745 source.n383 source.n362 2.71565
R746 source.n402 source.n401 2.71565
R747 source.n311 source.n290 2.71565
R748 source.n330 source.n329 2.71565
R749 source.n54 source.n53 2.71565
R750 source.n36 source.n15 2.71565
R751 source.n126 source.n125 2.71565
R752 source.n108 source.n87 2.71565
R753 source.n192 source.n191 2.71565
R754 source.n174 source.n153 2.71565
R755 source.n264 source.n263 2.71565
R756 source.n246 source.n225 2.71565
R757 source.n522 source.n498 1.93989
R758 source.n536 source.n492 1.93989
R759 source.n450 source.n426 1.93989
R760 source.n464 source.n420 1.93989
R761 source.n384 source.n360 1.93989
R762 source.n398 source.n354 1.93989
R763 source.n312 source.n288 1.93989
R764 source.n326 source.n282 1.93989
R765 source.n50 source.n6 1.93989
R766 source.n37 source.n13 1.93989
R767 source.n122 source.n78 1.93989
R768 source.n109 source.n85 1.93989
R769 source.n188 source.n144 1.93989
R770 source.n175 source.n151 1.93989
R771 source.n260 source.n216 1.93989
R772 source.n247 source.n223 1.93989
R773 source.n484 source.t0 1.6505
R774 source.n484 source.t12 1.6505
R775 source.n482 source.t3 1.6505
R776 source.n482 source.t10 1.6505
R777 source.n480 source.t9 1.6505
R778 source.n480 source.t11 1.6505
R779 source.n346 source.t27 1.6505
R780 source.n346 source.t20 1.6505
R781 source.n344 source.t30 1.6505
R782 source.n344 source.t31 1.6505
R783 source.n342 source.t28 1.6505
R784 source.n342 source.t25 1.6505
R785 source.n66 source.t16 1.6505
R786 source.n66 source.t24 1.6505
R787 source.n68 source.t26 1.6505
R788 source.n68 source.t22 1.6505
R789 source.n70 source.t23 1.6505
R790 source.n70 source.t18 1.6505
R791 source.n204 source.t14 1.6505
R792 source.n204 source.t7 1.6505
R793 source.n206 source.t5 1.6505
R794 source.n206 source.t1 1.6505
R795 source.n208 source.t2 1.6505
R796 source.n208 source.t4 1.6505
R797 source.n527 source.n525 1.16414
R798 source.n535 source.n494 1.16414
R799 source.n455 source.n453 1.16414
R800 source.n463 source.n422 1.16414
R801 source.n389 source.n387 1.16414
R802 source.n397 source.n356 1.16414
R803 source.n317 source.n315 1.16414
R804 source.n325 source.n284 1.16414
R805 source.n49 source.n8 1.16414
R806 source.n41 source.n40 1.16414
R807 source.n121 source.n80 1.16414
R808 source.n113 source.n112 1.16414
R809 source.n187 source.n146 1.16414
R810 source.n179 source.n178 1.16414
R811 source.n259 source.n218 1.16414
R812 source.n251 source.n250 1.16414
R813 source.n275 source.n209 0.716017
R814 source.n209 source.n207 0.716017
R815 source.n207 source.n205 0.716017
R816 source.n205 source.n203 0.716017
R817 source.n137 source.n71 0.716017
R818 source.n71 source.n69 0.716017
R819 source.n69 source.n67 0.716017
R820 source.n67 source.n65 0.716017
R821 source.n343 source.n341 0.716017
R822 source.n345 source.n343 0.716017
R823 source.n347 source.n345 0.716017
R824 source.n413 source.n347 0.716017
R825 source.n481 source.n479 0.716017
R826 source.n483 source.n481 0.716017
R827 source.n485 source.n483 0.716017
R828 source.n551 source.n485 0.716017
R829 source.n203 source.n137 0.470328
R830 source.n479 source.n413 0.470328
R831 source.n526 source.n496 0.388379
R832 source.n532 source.n531 0.388379
R833 source.n454 source.n424 0.388379
R834 source.n460 source.n459 0.388379
R835 source.n388 source.n358 0.388379
R836 source.n394 source.n393 0.388379
R837 source.n316 source.n286 0.388379
R838 source.n322 source.n321 0.388379
R839 source.n46 source.n45 0.388379
R840 source.n12 source.n10 0.388379
R841 source.n118 source.n117 0.388379
R842 source.n84 source.n82 0.388379
R843 source.n184 source.n183 0.388379
R844 source.n150 source.n148 0.388379
R845 source.n256 source.n255 0.388379
R846 source.n222 source.n220 0.388379
R847 source source.n552 0.188
R848 source.n508 source.n503 0.155672
R849 source.n515 source.n503 0.155672
R850 source.n516 source.n515 0.155672
R851 source.n516 source.n499 0.155672
R852 source.n523 source.n499 0.155672
R853 source.n524 source.n523 0.155672
R854 source.n524 source.n495 0.155672
R855 source.n533 source.n495 0.155672
R856 source.n534 source.n533 0.155672
R857 source.n534 source.n491 0.155672
R858 source.n541 source.n491 0.155672
R859 source.n542 source.n541 0.155672
R860 source.n542 source.n487 0.155672
R861 source.n549 source.n487 0.155672
R862 source.n436 source.n431 0.155672
R863 source.n443 source.n431 0.155672
R864 source.n444 source.n443 0.155672
R865 source.n444 source.n427 0.155672
R866 source.n451 source.n427 0.155672
R867 source.n452 source.n451 0.155672
R868 source.n452 source.n423 0.155672
R869 source.n461 source.n423 0.155672
R870 source.n462 source.n461 0.155672
R871 source.n462 source.n419 0.155672
R872 source.n469 source.n419 0.155672
R873 source.n470 source.n469 0.155672
R874 source.n470 source.n415 0.155672
R875 source.n477 source.n415 0.155672
R876 source.n370 source.n365 0.155672
R877 source.n377 source.n365 0.155672
R878 source.n378 source.n377 0.155672
R879 source.n378 source.n361 0.155672
R880 source.n385 source.n361 0.155672
R881 source.n386 source.n385 0.155672
R882 source.n386 source.n357 0.155672
R883 source.n395 source.n357 0.155672
R884 source.n396 source.n395 0.155672
R885 source.n396 source.n353 0.155672
R886 source.n403 source.n353 0.155672
R887 source.n404 source.n403 0.155672
R888 source.n404 source.n349 0.155672
R889 source.n411 source.n349 0.155672
R890 source.n298 source.n293 0.155672
R891 source.n305 source.n293 0.155672
R892 source.n306 source.n305 0.155672
R893 source.n306 source.n289 0.155672
R894 source.n313 source.n289 0.155672
R895 source.n314 source.n313 0.155672
R896 source.n314 source.n285 0.155672
R897 source.n323 source.n285 0.155672
R898 source.n324 source.n323 0.155672
R899 source.n324 source.n281 0.155672
R900 source.n331 source.n281 0.155672
R901 source.n332 source.n331 0.155672
R902 source.n332 source.n277 0.155672
R903 source.n339 source.n277 0.155672
R904 source.n63 source.n1 0.155672
R905 source.n56 source.n1 0.155672
R906 source.n56 source.n55 0.155672
R907 source.n55 source.n5 0.155672
R908 source.n48 source.n5 0.155672
R909 source.n48 source.n47 0.155672
R910 source.n47 source.n9 0.155672
R911 source.n39 source.n9 0.155672
R912 source.n39 source.n38 0.155672
R913 source.n38 source.n14 0.155672
R914 source.n31 source.n14 0.155672
R915 source.n31 source.n30 0.155672
R916 source.n30 source.n18 0.155672
R917 source.n23 source.n18 0.155672
R918 source.n135 source.n73 0.155672
R919 source.n128 source.n73 0.155672
R920 source.n128 source.n127 0.155672
R921 source.n127 source.n77 0.155672
R922 source.n120 source.n77 0.155672
R923 source.n120 source.n119 0.155672
R924 source.n119 source.n81 0.155672
R925 source.n111 source.n81 0.155672
R926 source.n111 source.n110 0.155672
R927 source.n110 source.n86 0.155672
R928 source.n103 source.n86 0.155672
R929 source.n103 source.n102 0.155672
R930 source.n102 source.n90 0.155672
R931 source.n95 source.n90 0.155672
R932 source.n201 source.n139 0.155672
R933 source.n194 source.n139 0.155672
R934 source.n194 source.n193 0.155672
R935 source.n193 source.n143 0.155672
R936 source.n186 source.n143 0.155672
R937 source.n186 source.n185 0.155672
R938 source.n185 source.n147 0.155672
R939 source.n177 source.n147 0.155672
R940 source.n177 source.n176 0.155672
R941 source.n176 source.n152 0.155672
R942 source.n169 source.n152 0.155672
R943 source.n169 source.n168 0.155672
R944 source.n168 source.n156 0.155672
R945 source.n161 source.n156 0.155672
R946 source.n273 source.n211 0.155672
R947 source.n266 source.n211 0.155672
R948 source.n266 source.n265 0.155672
R949 source.n265 source.n215 0.155672
R950 source.n258 source.n215 0.155672
R951 source.n258 source.n257 0.155672
R952 source.n257 source.n219 0.155672
R953 source.n249 source.n219 0.155672
R954 source.n249 source.n248 0.155672
R955 source.n248 source.n224 0.155672
R956 source.n241 source.n224 0.155672
R957 source.n241 source.n240 0.155672
R958 source.n240 source.n228 0.155672
R959 source.n233 source.n228 0.155672
R960 minus.n5 minus.t14 677.948
R961 minus.n27 minus.t2 677.948
R962 minus.n6 minus.t3 656.966
R963 minus.n8 minus.t6 656.966
R964 minus.n12 minus.t15 656.966
R965 minus.n13 minus.t5 656.966
R966 minus.n1 minus.t10 656.966
R967 minus.n19 minus.t0 656.966
R968 minus.n20 minus.t11 656.966
R969 minus.n28 minus.t1 656.966
R970 minus.n30 minus.t9 656.966
R971 minus.n34 minus.t8 656.966
R972 minus.n35 minus.t4 656.966
R973 minus.n23 minus.t13 656.966
R974 minus.n41 minus.t12 656.966
R975 minus.n42 minus.t7 656.966
R976 minus.n21 minus.n20 161.3
R977 minus.n19 minus.n0 161.3
R978 minus.n18 minus.n17 161.3
R979 minus.n16 minus.n1 161.3
R980 minus.n15 minus.n14 161.3
R981 minus.n13 minus.n2 161.3
R982 minus.n12 minus.n11 161.3
R983 minus.n10 minus.n3 161.3
R984 minus.n9 minus.n8 161.3
R985 minus.n7 minus.n4 161.3
R986 minus.n43 minus.n42 161.3
R987 minus.n41 minus.n22 161.3
R988 minus.n40 minus.n39 161.3
R989 minus.n38 minus.n23 161.3
R990 minus.n37 minus.n36 161.3
R991 minus.n35 minus.n24 161.3
R992 minus.n34 minus.n33 161.3
R993 minus.n32 minus.n25 161.3
R994 minus.n31 minus.n30 161.3
R995 minus.n29 minus.n26 161.3
R996 minus.n5 minus.n4 70.4033
R997 minus.n27 minus.n26 70.4033
R998 minus.n13 minus.n12 48.2005
R999 minus.n20 minus.n19 48.2005
R1000 minus.n35 minus.n34 48.2005
R1001 minus.n42 minus.n41 48.2005
R1002 minus.n44 minus.n21 37.5535
R1003 minus.n8 minus.n7 37.246
R1004 minus.n18 minus.n1 37.246
R1005 minus.n30 minus.n29 37.246
R1006 minus.n40 minus.n23 37.246
R1007 minus.n8 minus.n3 35.7853
R1008 minus.n14 minus.n1 35.7853
R1009 minus.n30 minus.n25 35.7853
R1010 minus.n36 minus.n23 35.7853
R1011 minus.n6 minus.n5 20.9576
R1012 minus.n28 minus.n27 20.9576
R1013 minus.n12 minus.n3 12.4157
R1014 minus.n14 minus.n13 12.4157
R1015 minus.n34 minus.n25 12.4157
R1016 minus.n36 minus.n35 12.4157
R1017 minus.n7 minus.n6 10.955
R1018 minus.n19 minus.n18 10.955
R1019 minus.n29 minus.n28 10.955
R1020 minus.n41 minus.n40 10.955
R1021 minus.n44 minus.n43 6.56111
R1022 minus.n21 minus.n0 0.189894
R1023 minus.n17 minus.n0 0.189894
R1024 minus.n17 minus.n16 0.189894
R1025 minus.n16 minus.n15 0.189894
R1026 minus.n15 minus.n2 0.189894
R1027 minus.n11 minus.n2 0.189894
R1028 minus.n11 minus.n10 0.189894
R1029 minus.n10 minus.n9 0.189894
R1030 minus.n9 minus.n4 0.189894
R1031 minus.n31 minus.n26 0.189894
R1032 minus.n32 minus.n31 0.189894
R1033 minus.n33 minus.n32 0.189894
R1034 minus.n33 minus.n24 0.189894
R1035 minus.n37 minus.n24 0.189894
R1036 minus.n38 minus.n37 0.189894
R1037 minus.n39 minus.n38 0.189894
R1038 minus.n39 minus.n22 0.189894
R1039 minus.n43 minus.n22 0.189894
R1040 minus minus.n44 0.188
R1041 drain_right.n5 drain_right.n3 60.268
R1042 drain_right.n2 drain_right.n0 60.268
R1043 drain_right.n9 drain_right.n7 60.268
R1044 drain_right.n9 drain_right.n8 59.5527
R1045 drain_right.n11 drain_right.n10 59.5527
R1046 drain_right.n13 drain_right.n12 59.5527
R1047 drain_right.n5 drain_right.n4 59.5525
R1048 drain_right.n2 drain_right.n1 59.5525
R1049 drain_right drain_right.n6 31.4647
R1050 drain_right drain_right.n13 6.36873
R1051 drain_right.n3 drain_right.t3 1.6505
R1052 drain_right.n3 drain_right.t8 1.6505
R1053 drain_right.n4 drain_right.t11 1.6505
R1054 drain_right.n4 drain_right.t2 1.6505
R1055 drain_right.n1 drain_right.t6 1.6505
R1056 drain_right.n1 drain_right.t7 1.6505
R1057 drain_right.n0 drain_right.t13 1.6505
R1058 drain_right.n0 drain_right.t14 1.6505
R1059 drain_right.n7 drain_right.t12 1.6505
R1060 drain_right.n7 drain_right.t1 1.6505
R1061 drain_right.n8 drain_right.t0 1.6505
R1062 drain_right.n8 drain_right.t9 1.6505
R1063 drain_right.n10 drain_right.t5 1.6505
R1064 drain_right.n10 drain_right.t10 1.6505
R1065 drain_right.n12 drain_right.t4 1.6505
R1066 drain_right.n12 drain_right.t15 1.6505
R1067 drain_right.n13 drain_right.n11 0.716017
R1068 drain_right.n11 drain_right.n9 0.716017
R1069 drain_right.n6 drain_right.n5 0.302913
R1070 drain_right.n6 drain_right.n2 0.302913
C0 minus source 8.23696f
C1 plus drain_right 0.372806f
C2 plus drain_left 8.57739f
C3 plus minus 5.90663f
C4 drain_left drain_right 1.15071f
C5 minus drain_right 8.36021f
C6 drain_left minus 0.172419f
C7 plus source 8.250999f
C8 drain_right source 23.5319f
C9 drain_left source 23.530699f
C10 drain_right a_n2210_n3288# 6.57098f
C11 drain_left a_n2210_n3288# 6.89323f
C12 source a_n2210_n3288# 8.997727f
C13 minus a_n2210_n3288# 8.740124f
C14 plus a_n2210_n3288# 10.608491f
C15 drain_right.t13 a_n2210_n3288# 0.277535f
C16 drain_right.t14 a_n2210_n3288# 0.277535f
C17 drain_right.n0 a_n2210_n3288# 2.47429f
C18 drain_right.t6 a_n2210_n3288# 0.277535f
C19 drain_right.t7 a_n2210_n3288# 0.277535f
C20 drain_right.n1 a_n2210_n3288# 2.46963f
C21 drain_right.n2 a_n2210_n3288# 0.731579f
C22 drain_right.t3 a_n2210_n3288# 0.277535f
C23 drain_right.t8 a_n2210_n3288# 0.277535f
C24 drain_right.n3 a_n2210_n3288# 2.47429f
C25 drain_right.t11 a_n2210_n3288# 0.277535f
C26 drain_right.t2 a_n2210_n3288# 0.277535f
C27 drain_right.n4 a_n2210_n3288# 2.46963f
C28 drain_right.n5 a_n2210_n3288# 0.731579f
C29 drain_right.n6 a_n2210_n3288# 1.4977f
C30 drain_right.t12 a_n2210_n3288# 0.277535f
C31 drain_right.t1 a_n2210_n3288# 0.277535f
C32 drain_right.n7 a_n2210_n3288# 2.47429f
C33 drain_right.t0 a_n2210_n3288# 0.277535f
C34 drain_right.t9 a_n2210_n3288# 0.277535f
C35 drain_right.n8 a_n2210_n3288# 2.46964f
C36 drain_right.n9 a_n2210_n3288# 0.768283f
C37 drain_right.t5 a_n2210_n3288# 0.277535f
C38 drain_right.t10 a_n2210_n3288# 0.277535f
C39 drain_right.n10 a_n2210_n3288# 2.46964f
C40 drain_right.n11 a_n2210_n3288# 0.380572f
C41 drain_right.t4 a_n2210_n3288# 0.277535f
C42 drain_right.t15 a_n2210_n3288# 0.277535f
C43 drain_right.n12 a_n2210_n3288# 2.46964f
C44 drain_right.n13 a_n2210_n3288# 0.632018f
C45 minus.n0 a_n2210_n3288# 0.045066f
C46 minus.t10 a_n2210_n3288# 0.771034f
C47 minus.n1 a_n2210_n3288# 0.315743f
C48 minus.n2 a_n2210_n3288# 0.045066f
C49 minus.n3 a_n2210_n3288# 0.010226f
C50 minus.t15 a_n2210_n3288# 0.771034f
C51 minus.n4 a_n2210_n3288# 0.143482f
C52 minus.t3 a_n2210_n3288# 0.771034f
C53 minus.t14 a_n2210_n3288# 0.780661f
C54 minus.n5 a_n2210_n3288# 0.301721f
C55 minus.n6 a_n2210_n3288# 0.313104f
C56 minus.n7 a_n2210_n3288# 0.010226f
C57 minus.t6 a_n2210_n3288# 0.771034f
C58 minus.n8 a_n2210_n3288# 0.315743f
C59 minus.n9 a_n2210_n3288# 0.045066f
C60 minus.n10 a_n2210_n3288# 0.045066f
C61 minus.n11 a_n2210_n3288# 0.045066f
C62 minus.n12 a_n2210_n3288# 0.313382f
C63 minus.t5 a_n2210_n3288# 0.771034f
C64 minus.n13 a_n2210_n3288# 0.313382f
C65 minus.n14 a_n2210_n3288# 0.010226f
C66 minus.n15 a_n2210_n3288# 0.045066f
C67 minus.n16 a_n2210_n3288# 0.045066f
C68 minus.n17 a_n2210_n3288# 0.045066f
C69 minus.n18 a_n2210_n3288# 0.010226f
C70 minus.t0 a_n2210_n3288# 0.771034f
C71 minus.n19 a_n2210_n3288# 0.313104f
C72 minus.t11 a_n2210_n3288# 0.771034f
C73 minus.n20 a_n2210_n3288# 0.31102f
C74 minus.n21 a_n2210_n3288# 1.6885f
C75 minus.n22 a_n2210_n3288# 0.045066f
C76 minus.t13 a_n2210_n3288# 0.771034f
C77 minus.n23 a_n2210_n3288# 0.315743f
C78 minus.n24 a_n2210_n3288# 0.045066f
C79 minus.n25 a_n2210_n3288# 0.010226f
C80 minus.n26 a_n2210_n3288# 0.143482f
C81 minus.t2 a_n2210_n3288# 0.780661f
C82 minus.n27 a_n2210_n3288# 0.301721f
C83 minus.t1 a_n2210_n3288# 0.771034f
C84 minus.n28 a_n2210_n3288# 0.313104f
C85 minus.n29 a_n2210_n3288# 0.010226f
C86 minus.t9 a_n2210_n3288# 0.771034f
C87 minus.n30 a_n2210_n3288# 0.315743f
C88 minus.n31 a_n2210_n3288# 0.045066f
C89 minus.n32 a_n2210_n3288# 0.045066f
C90 minus.n33 a_n2210_n3288# 0.045066f
C91 minus.t8 a_n2210_n3288# 0.771034f
C92 minus.n34 a_n2210_n3288# 0.313382f
C93 minus.t4 a_n2210_n3288# 0.771034f
C94 minus.n35 a_n2210_n3288# 0.313382f
C95 minus.n36 a_n2210_n3288# 0.010226f
C96 minus.n37 a_n2210_n3288# 0.045066f
C97 minus.n38 a_n2210_n3288# 0.045066f
C98 minus.n39 a_n2210_n3288# 0.045066f
C99 minus.n40 a_n2210_n3288# 0.010226f
C100 minus.t12 a_n2210_n3288# 0.771034f
C101 minus.n41 a_n2210_n3288# 0.313104f
C102 minus.t7 a_n2210_n3288# 0.771034f
C103 minus.n42 a_n2210_n3288# 0.31102f
C104 minus.n43 a_n2210_n3288# 0.301097f
C105 minus.n44 a_n2210_n3288# 2.04079f
C106 source.n0 a_n2210_n3288# 0.032843f
C107 source.n1 a_n2210_n3288# 0.024794f
C108 source.n2 a_n2210_n3288# 0.013323f
C109 source.n3 a_n2210_n3288# 0.031492f
C110 source.n4 a_n2210_n3288# 0.014107f
C111 source.n5 a_n2210_n3288# 0.024794f
C112 source.n6 a_n2210_n3288# 0.013323f
C113 source.n7 a_n2210_n3288# 0.031492f
C114 source.n8 a_n2210_n3288# 0.014107f
C115 source.n9 a_n2210_n3288# 0.024794f
C116 source.n10 a_n2210_n3288# 0.013715f
C117 source.n11 a_n2210_n3288# 0.031492f
C118 source.n12 a_n2210_n3288# 0.013323f
C119 source.n13 a_n2210_n3288# 0.014107f
C120 source.n14 a_n2210_n3288# 0.024794f
C121 source.n15 a_n2210_n3288# 0.013323f
C122 source.n16 a_n2210_n3288# 0.031492f
C123 source.n17 a_n2210_n3288# 0.014107f
C124 source.n18 a_n2210_n3288# 0.024794f
C125 source.n19 a_n2210_n3288# 0.013323f
C126 source.n20 a_n2210_n3288# 0.023619f
C127 source.n21 a_n2210_n3288# 0.022262f
C128 source.t19 a_n2210_n3288# 0.053187f
C129 source.n22 a_n2210_n3288# 0.178764f
C130 source.n23 a_n2210_n3288# 1.25083f
C131 source.n24 a_n2210_n3288# 0.013323f
C132 source.n25 a_n2210_n3288# 0.014107f
C133 source.n26 a_n2210_n3288# 0.031492f
C134 source.n27 a_n2210_n3288# 0.031492f
C135 source.n28 a_n2210_n3288# 0.014107f
C136 source.n29 a_n2210_n3288# 0.013323f
C137 source.n30 a_n2210_n3288# 0.024794f
C138 source.n31 a_n2210_n3288# 0.024794f
C139 source.n32 a_n2210_n3288# 0.013323f
C140 source.n33 a_n2210_n3288# 0.014107f
C141 source.n34 a_n2210_n3288# 0.031492f
C142 source.n35 a_n2210_n3288# 0.031492f
C143 source.n36 a_n2210_n3288# 0.014107f
C144 source.n37 a_n2210_n3288# 0.013323f
C145 source.n38 a_n2210_n3288# 0.024794f
C146 source.n39 a_n2210_n3288# 0.024794f
C147 source.n40 a_n2210_n3288# 0.013323f
C148 source.n41 a_n2210_n3288# 0.014107f
C149 source.n42 a_n2210_n3288# 0.031492f
C150 source.n43 a_n2210_n3288# 0.031492f
C151 source.n44 a_n2210_n3288# 0.031492f
C152 source.n45 a_n2210_n3288# 0.013715f
C153 source.n46 a_n2210_n3288# 0.013323f
C154 source.n47 a_n2210_n3288# 0.024794f
C155 source.n48 a_n2210_n3288# 0.024794f
C156 source.n49 a_n2210_n3288# 0.013323f
C157 source.n50 a_n2210_n3288# 0.014107f
C158 source.n51 a_n2210_n3288# 0.031492f
C159 source.n52 a_n2210_n3288# 0.031492f
C160 source.n53 a_n2210_n3288# 0.014107f
C161 source.n54 a_n2210_n3288# 0.013323f
C162 source.n55 a_n2210_n3288# 0.024794f
C163 source.n56 a_n2210_n3288# 0.024794f
C164 source.n57 a_n2210_n3288# 0.013323f
C165 source.n58 a_n2210_n3288# 0.014107f
C166 source.n59 a_n2210_n3288# 0.031492f
C167 source.n60 a_n2210_n3288# 0.064624f
C168 source.n61 a_n2210_n3288# 0.014107f
C169 source.n62 a_n2210_n3288# 0.013323f
C170 source.n63 a_n2210_n3288# 0.053246f
C171 source.n64 a_n2210_n3288# 0.035666f
C172 source.n65 a_n2210_n3288# 1.02044f
C173 source.t16 a_n2210_n3288# 0.235119f
C174 source.t24 a_n2210_n3288# 0.235119f
C175 source.n66 a_n2210_n3288# 2.01309f
C176 source.n67 a_n2210_n3288# 0.36782f
C177 source.t26 a_n2210_n3288# 0.235119f
C178 source.t22 a_n2210_n3288# 0.235119f
C179 source.n68 a_n2210_n3288# 2.01309f
C180 source.n69 a_n2210_n3288# 0.36782f
C181 source.t23 a_n2210_n3288# 0.235119f
C182 source.t18 a_n2210_n3288# 0.235119f
C183 source.n70 a_n2210_n3288# 2.01309f
C184 source.n71 a_n2210_n3288# 0.36782f
C185 source.n72 a_n2210_n3288# 0.032843f
C186 source.n73 a_n2210_n3288# 0.024794f
C187 source.n74 a_n2210_n3288# 0.013323f
C188 source.n75 a_n2210_n3288# 0.031492f
C189 source.n76 a_n2210_n3288# 0.014107f
C190 source.n77 a_n2210_n3288# 0.024794f
C191 source.n78 a_n2210_n3288# 0.013323f
C192 source.n79 a_n2210_n3288# 0.031492f
C193 source.n80 a_n2210_n3288# 0.014107f
C194 source.n81 a_n2210_n3288# 0.024794f
C195 source.n82 a_n2210_n3288# 0.013715f
C196 source.n83 a_n2210_n3288# 0.031492f
C197 source.n84 a_n2210_n3288# 0.013323f
C198 source.n85 a_n2210_n3288# 0.014107f
C199 source.n86 a_n2210_n3288# 0.024794f
C200 source.n87 a_n2210_n3288# 0.013323f
C201 source.n88 a_n2210_n3288# 0.031492f
C202 source.n89 a_n2210_n3288# 0.014107f
C203 source.n90 a_n2210_n3288# 0.024794f
C204 source.n91 a_n2210_n3288# 0.013323f
C205 source.n92 a_n2210_n3288# 0.023619f
C206 source.n93 a_n2210_n3288# 0.022262f
C207 source.t29 a_n2210_n3288# 0.053187f
C208 source.n94 a_n2210_n3288# 0.178764f
C209 source.n95 a_n2210_n3288# 1.25083f
C210 source.n96 a_n2210_n3288# 0.013323f
C211 source.n97 a_n2210_n3288# 0.014107f
C212 source.n98 a_n2210_n3288# 0.031492f
C213 source.n99 a_n2210_n3288# 0.031492f
C214 source.n100 a_n2210_n3288# 0.014107f
C215 source.n101 a_n2210_n3288# 0.013323f
C216 source.n102 a_n2210_n3288# 0.024794f
C217 source.n103 a_n2210_n3288# 0.024794f
C218 source.n104 a_n2210_n3288# 0.013323f
C219 source.n105 a_n2210_n3288# 0.014107f
C220 source.n106 a_n2210_n3288# 0.031492f
C221 source.n107 a_n2210_n3288# 0.031492f
C222 source.n108 a_n2210_n3288# 0.014107f
C223 source.n109 a_n2210_n3288# 0.013323f
C224 source.n110 a_n2210_n3288# 0.024794f
C225 source.n111 a_n2210_n3288# 0.024794f
C226 source.n112 a_n2210_n3288# 0.013323f
C227 source.n113 a_n2210_n3288# 0.014107f
C228 source.n114 a_n2210_n3288# 0.031492f
C229 source.n115 a_n2210_n3288# 0.031492f
C230 source.n116 a_n2210_n3288# 0.031492f
C231 source.n117 a_n2210_n3288# 0.013715f
C232 source.n118 a_n2210_n3288# 0.013323f
C233 source.n119 a_n2210_n3288# 0.024794f
C234 source.n120 a_n2210_n3288# 0.024794f
C235 source.n121 a_n2210_n3288# 0.013323f
C236 source.n122 a_n2210_n3288# 0.014107f
C237 source.n123 a_n2210_n3288# 0.031492f
C238 source.n124 a_n2210_n3288# 0.031492f
C239 source.n125 a_n2210_n3288# 0.014107f
C240 source.n126 a_n2210_n3288# 0.013323f
C241 source.n127 a_n2210_n3288# 0.024794f
C242 source.n128 a_n2210_n3288# 0.024794f
C243 source.n129 a_n2210_n3288# 0.013323f
C244 source.n130 a_n2210_n3288# 0.014107f
C245 source.n131 a_n2210_n3288# 0.031492f
C246 source.n132 a_n2210_n3288# 0.064624f
C247 source.n133 a_n2210_n3288# 0.014107f
C248 source.n134 a_n2210_n3288# 0.013323f
C249 source.n135 a_n2210_n3288# 0.053246f
C250 source.n136 a_n2210_n3288# 0.035666f
C251 source.n137 a_n2210_n3288# 0.113587f
C252 source.n138 a_n2210_n3288# 0.032843f
C253 source.n139 a_n2210_n3288# 0.024794f
C254 source.n140 a_n2210_n3288# 0.013323f
C255 source.n141 a_n2210_n3288# 0.031492f
C256 source.n142 a_n2210_n3288# 0.014107f
C257 source.n143 a_n2210_n3288# 0.024794f
C258 source.n144 a_n2210_n3288# 0.013323f
C259 source.n145 a_n2210_n3288# 0.031492f
C260 source.n146 a_n2210_n3288# 0.014107f
C261 source.n147 a_n2210_n3288# 0.024794f
C262 source.n148 a_n2210_n3288# 0.013715f
C263 source.n149 a_n2210_n3288# 0.031492f
C264 source.n150 a_n2210_n3288# 0.013323f
C265 source.n151 a_n2210_n3288# 0.014107f
C266 source.n152 a_n2210_n3288# 0.024794f
C267 source.n153 a_n2210_n3288# 0.013323f
C268 source.n154 a_n2210_n3288# 0.031492f
C269 source.n155 a_n2210_n3288# 0.014107f
C270 source.n156 a_n2210_n3288# 0.024794f
C271 source.n157 a_n2210_n3288# 0.013323f
C272 source.n158 a_n2210_n3288# 0.023619f
C273 source.n159 a_n2210_n3288# 0.022262f
C274 source.t13 a_n2210_n3288# 0.053187f
C275 source.n160 a_n2210_n3288# 0.178764f
C276 source.n161 a_n2210_n3288# 1.25083f
C277 source.n162 a_n2210_n3288# 0.013323f
C278 source.n163 a_n2210_n3288# 0.014107f
C279 source.n164 a_n2210_n3288# 0.031492f
C280 source.n165 a_n2210_n3288# 0.031492f
C281 source.n166 a_n2210_n3288# 0.014107f
C282 source.n167 a_n2210_n3288# 0.013323f
C283 source.n168 a_n2210_n3288# 0.024794f
C284 source.n169 a_n2210_n3288# 0.024794f
C285 source.n170 a_n2210_n3288# 0.013323f
C286 source.n171 a_n2210_n3288# 0.014107f
C287 source.n172 a_n2210_n3288# 0.031492f
C288 source.n173 a_n2210_n3288# 0.031492f
C289 source.n174 a_n2210_n3288# 0.014107f
C290 source.n175 a_n2210_n3288# 0.013323f
C291 source.n176 a_n2210_n3288# 0.024794f
C292 source.n177 a_n2210_n3288# 0.024794f
C293 source.n178 a_n2210_n3288# 0.013323f
C294 source.n179 a_n2210_n3288# 0.014107f
C295 source.n180 a_n2210_n3288# 0.031492f
C296 source.n181 a_n2210_n3288# 0.031492f
C297 source.n182 a_n2210_n3288# 0.031492f
C298 source.n183 a_n2210_n3288# 0.013715f
C299 source.n184 a_n2210_n3288# 0.013323f
C300 source.n185 a_n2210_n3288# 0.024794f
C301 source.n186 a_n2210_n3288# 0.024794f
C302 source.n187 a_n2210_n3288# 0.013323f
C303 source.n188 a_n2210_n3288# 0.014107f
C304 source.n189 a_n2210_n3288# 0.031492f
C305 source.n190 a_n2210_n3288# 0.031492f
C306 source.n191 a_n2210_n3288# 0.014107f
C307 source.n192 a_n2210_n3288# 0.013323f
C308 source.n193 a_n2210_n3288# 0.024794f
C309 source.n194 a_n2210_n3288# 0.024794f
C310 source.n195 a_n2210_n3288# 0.013323f
C311 source.n196 a_n2210_n3288# 0.014107f
C312 source.n197 a_n2210_n3288# 0.031492f
C313 source.n198 a_n2210_n3288# 0.064624f
C314 source.n199 a_n2210_n3288# 0.014107f
C315 source.n200 a_n2210_n3288# 0.013323f
C316 source.n201 a_n2210_n3288# 0.053246f
C317 source.n202 a_n2210_n3288# 0.035666f
C318 source.n203 a_n2210_n3288# 0.113587f
C319 source.t14 a_n2210_n3288# 0.235119f
C320 source.t7 a_n2210_n3288# 0.235119f
C321 source.n204 a_n2210_n3288# 2.01309f
C322 source.n205 a_n2210_n3288# 0.36782f
C323 source.t5 a_n2210_n3288# 0.235119f
C324 source.t1 a_n2210_n3288# 0.235119f
C325 source.n206 a_n2210_n3288# 2.01309f
C326 source.n207 a_n2210_n3288# 0.36782f
C327 source.t2 a_n2210_n3288# 0.235119f
C328 source.t4 a_n2210_n3288# 0.235119f
C329 source.n208 a_n2210_n3288# 2.01309f
C330 source.n209 a_n2210_n3288# 0.36782f
C331 source.n210 a_n2210_n3288# 0.032843f
C332 source.n211 a_n2210_n3288# 0.024794f
C333 source.n212 a_n2210_n3288# 0.013323f
C334 source.n213 a_n2210_n3288# 0.031492f
C335 source.n214 a_n2210_n3288# 0.014107f
C336 source.n215 a_n2210_n3288# 0.024794f
C337 source.n216 a_n2210_n3288# 0.013323f
C338 source.n217 a_n2210_n3288# 0.031492f
C339 source.n218 a_n2210_n3288# 0.014107f
C340 source.n219 a_n2210_n3288# 0.024794f
C341 source.n220 a_n2210_n3288# 0.013715f
C342 source.n221 a_n2210_n3288# 0.031492f
C343 source.n222 a_n2210_n3288# 0.013323f
C344 source.n223 a_n2210_n3288# 0.014107f
C345 source.n224 a_n2210_n3288# 0.024794f
C346 source.n225 a_n2210_n3288# 0.013323f
C347 source.n226 a_n2210_n3288# 0.031492f
C348 source.n227 a_n2210_n3288# 0.014107f
C349 source.n228 a_n2210_n3288# 0.024794f
C350 source.n229 a_n2210_n3288# 0.013323f
C351 source.n230 a_n2210_n3288# 0.023619f
C352 source.n231 a_n2210_n3288# 0.022262f
C353 source.t8 a_n2210_n3288# 0.053187f
C354 source.n232 a_n2210_n3288# 0.178764f
C355 source.n233 a_n2210_n3288# 1.25083f
C356 source.n234 a_n2210_n3288# 0.013323f
C357 source.n235 a_n2210_n3288# 0.014107f
C358 source.n236 a_n2210_n3288# 0.031492f
C359 source.n237 a_n2210_n3288# 0.031492f
C360 source.n238 a_n2210_n3288# 0.014107f
C361 source.n239 a_n2210_n3288# 0.013323f
C362 source.n240 a_n2210_n3288# 0.024794f
C363 source.n241 a_n2210_n3288# 0.024794f
C364 source.n242 a_n2210_n3288# 0.013323f
C365 source.n243 a_n2210_n3288# 0.014107f
C366 source.n244 a_n2210_n3288# 0.031492f
C367 source.n245 a_n2210_n3288# 0.031492f
C368 source.n246 a_n2210_n3288# 0.014107f
C369 source.n247 a_n2210_n3288# 0.013323f
C370 source.n248 a_n2210_n3288# 0.024794f
C371 source.n249 a_n2210_n3288# 0.024794f
C372 source.n250 a_n2210_n3288# 0.013323f
C373 source.n251 a_n2210_n3288# 0.014107f
C374 source.n252 a_n2210_n3288# 0.031492f
C375 source.n253 a_n2210_n3288# 0.031492f
C376 source.n254 a_n2210_n3288# 0.031492f
C377 source.n255 a_n2210_n3288# 0.013715f
C378 source.n256 a_n2210_n3288# 0.013323f
C379 source.n257 a_n2210_n3288# 0.024794f
C380 source.n258 a_n2210_n3288# 0.024794f
C381 source.n259 a_n2210_n3288# 0.013323f
C382 source.n260 a_n2210_n3288# 0.014107f
C383 source.n261 a_n2210_n3288# 0.031492f
C384 source.n262 a_n2210_n3288# 0.031492f
C385 source.n263 a_n2210_n3288# 0.014107f
C386 source.n264 a_n2210_n3288# 0.013323f
C387 source.n265 a_n2210_n3288# 0.024794f
C388 source.n266 a_n2210_n3288# 0.024794f
C389 source.n267 a_n2210_n3288# 0.013323f
C390 source.n268 a_n2210_n3288# 0.014107f
C391 source.n269 a_n2210_n3288# 0.031492f
C392 source.n270 a_n2210_n3288# 0.064624f
C393 source.n271 a_n2210_n3288# 0.014107f
C394 source.n272 a_n2210_n3288# 0.013323f
C395 source.n273 a_n2210_n3288# 0.053246f
C396 source.n274 a_n2210_n3288# 0.035666f
C397 source.n275 a_n2210_n3288# 1.41527f
C398 source.n276 a_n2210_n3288# 0.032843f
C399 source.n277 a_n2210_n3288# 0.024794f
C400 source.n278 a_n2210_n3288# 0.013323f
C401 source.n279 a_n2210_n3288# 0.031492f
C402 source.n280 a_n2210_n3288# 0.014107f
C403 source.n281 a_n2210_n3288# 0.024794f
C404 source.n282 a_n2210_n3288# 0.013323f
C405 source.n283 a_n2210_n3288# 0.031492f
C406 source.n284 a_n2210_n3288# 0.014107f
C407 source.n285 a_n2210_n3288# 0.024794f
C408 source.n286 a_n2210_n3288# 0.013715f
C409 source.n287 a_n2210_n3288# 0.031492f
C410 source.n288 a_n2210_n3288# 0.014107f
C411 source.n289 a_n2210_n3288# 0.024794f
C412 source.n290 a_n2210_n3288# 0.013323f
C413 source.n291 a_n2210_n3288# 0.031492f
C414 source.n292 a_n2210_n3288# 0.014107f
C415 source.n293 a_n2210_n3288# 0.024794f
C416 source.n294 a_n2210_n3288# 0.013323f
C417 source.n295 a_n2210_n3288# 0.023619f
C418 source.n296 a_n2210_n3288# 0.022262f
C419 source.t17 a_n2210_n3288# 0.053187f
C420 source.n297 a_n2210_n3288# 0.178764f
C421 source.n298 a_n2210_n3288# 1.25083f
C422 source.n299 a_n2210_n3288# 0.013323f
C423 source.n300 a_n2210_n3288# 0.014107f
C424 source.n301 a_n2210_n3288# 0.031492f
C425 source.n302 a_n2210_n3288# 0.031492f
C426 source.n303 a_n2210_n3288# 0.014107f
C427 source.n304 a_n2210_n3288# 0.013323f
C428 source.n305 a_n2210_n3288# 0.024794f
C429 source.n306 a_n2210_n3288# 0.024794f
C430 source.n307 a_n2210_n3288# 0.013323f
C431 source.n308 a_n2210_n3288# 0.014107f
C432 source.n309 a_n2210_n3288# 0.031492f
C433 source.n310 a_n2210_n3288# 0.031492f
C434 source.n311 a_n2210_n3288# 0.014107f
C435 source.n312 a_n2210_n3288# 0.013323f
C436 source.n313 a_n2210_n3288# 0.024794f
C437 source.n314 a_n2210_n3288# 0.024794f
C438 source.n315 a_n2210_n3288# 0.013323f
C439 source.n316 a_n2210_n3288# 0.013323f
C440 source.n317 a_n2210_n3288# 0.014107f
C441 source.n318 a_n2210_n3288# 0.031492f
C442 source.n319 a_n2210_n3288# 0.031492f
C443 source.n320 a_n2210_n3288# 0.031492f
C444 source.n321 a_n2210_n3288# 0.013715f
C445 source.n322 a_n2210_n3288# 0.013323f
C446 source.n323 a_n2210_n3288# 0.024794f
C447 source.n324 a_n2210_n3288# 0.024794f
C448 source.n325 a_n2210_n3288# 0.013323f
C449 source.n326 a_n2210_n3288# 0.014107f
C450 source.n327 a_n2210_n3288# 0.031492f
C451 source.n328 a_n2210_n3288# 0.031492f
C452 source.n329 a_n2210_n3288# 0.014107f
C453 source.n330 a_n2210_n3288# 0.013323f
C454 source.n331 a_n2210_n3288# 0.024794f
C455 source.n332 a_n2210_n3288# 0.024794f
C456 source.n333 a_n2210_n3288# 0.013323f
C457 source.n334 a_n2210_n3288# 0.014107f
C458 source.n335 a_n2210_n3288# 0.031492f
C459 source.n336 a_n2210_n3288# 0.064624f
C460 source.n337 a_n2210_n3288# 0.014107f
C461 source.n338 a_n2210_n3288# 0.013323f
C462 source.n339 a_n2210_n3288# 0.053246f
C463 source.n340 a_n2210_n3288# 0.035666f
C464 source.n341 a_n2210_n3288# 1.41527f
C465 source.t28 a_n2210_n3288# 0.235119f
C466 source.t25 a_n2210_n3288# 0.235119f
C467 source.n342 a_n2210_n3288# 2.01308f
C468 source.n343 a_n2210_n3288# 0.367832f
C469 source.t30 a_n2210_n3288# 0.235119f
C470 source.t31 a_n2210_n3288# 0.235119f
C471 source.n344 a_n2210_n3288# 2.01308f
C472 source.n345 a_n2210_n3288# 0.367832f
C473 source.t27 a_n2210_n3288# 0.235119f
C474 source.t20 a_n2210_n3288# 0.235119f
C475 source.n346 a_n2210_n3288# 2.01308f
C476 source.n347 a_n2210_n3288# 0.367832f
C477 source.n348 a_n2210_n3288# 0.032843f
C478 source.n349 a_n2210_n3288# 0.024794f
C479 source.n350 a_n2210_n3288# 0.013323f
C480 source.n351 a_n2210_n3288# 0.031492f
C481 source.n352 a_n2210_n3288# 0.014107f
C482 source.n353 a_n2210_n3288# 0.024794f
C483 source.n354 a_n2210_n3288# 0.013323f
C484 source.n355 a_n2210_n3288# 0.031492f
C485 source.n356 a_n2210_n3288# 0.014107f
C486 source.n357 a_n2210_n3288# 0.024794f
C487 source.n358 a_n2210_n3288# 0.013715f
C488 source.n359 a_n2210_n3288# 0.031492f
C489 source.n360 a_n2210_n3288# 0.014107f
C490 source.n361 a_n2210_n3288# 0.024794f
C491 source.n362 a_n2210_n3288# 0.013323f
C492 source.n363 a_n2210_n3288# 0.031492f
C493 source.n364 a_n2210_n3288# 0.014107f
C494 source.n365 a_n2210_n3288# 0.024794f
C495 source.n366 a_n2210_n3288# 0.013323f
C496 source.n367 a_n2210_n3288# 0.023619f
C497 source.n368 a_n2210_n3288# 0.022262f
C498 source.t21 a_n2210_n3288# 0.053187f
C499 source.n369 a_n2210_n3288# 0.178764f
C500 source.n370 a_n2210_n3288# 1.25083f
C501 source.n371 a_n2210_n3288# 0.013323f
C502 source.n372 a_n2210_n3288# 0.014107f
C503 source.n373 a_n2210_n3288# 0.031492f
C504 source.n374 a_n2210_n3288# 0.031492f
C505 source.n375 a_n2210_n3288# 0.014107f
C506 source.n376 a_n2210_n3288# 0.013323f
C507 source.n377 a_n2210_n3288# 0.024794f
C508 source.n378 a_n2210_n3288# 0.024794f
C509 source.n379 a_n2210_n3288# 0.013323f
C510 source.n380 a_n2210_n3288# 0.014107f
C511 source.n381 a_n2210_n3288# 0.031492f
C512 source.n382 a_n2210_n3288# 0.031492f
C513 source.n383 a_n2210_n3288# 0.014107f
C514 source.n384 a_n2210_n3288# 0.013323f
C515 source.n385 a_n2210_n3288# 0.024794f
C516 source.n386 a_n2210_n3288# 0.024794f
C517 source.n387 a_n2210_n3288# 0.013323f
C518 source.n388 a_n2210_n3288# 0.013323f
C519 source.n389 a_n2210_n3288# 0.014107f
C520 source.n390 a_n2210_n3288# 0.031492f
C521 source.n391 a_n2210_n3288# 0.031492f
C522 source.n392 a_n2210_n3288# 0.031492f
C523 source.n393 a_n2210_n3288# 0.013715f
C524 source.n394 a_n2210_n3288# 0.013323f
C525 source.n395 a_n2210_n3288# 0.024794f
C526 source.n396 a_n2210_n3288# 0.024794f
C527 source.n397 a_n2210_n3288# 0.013323f
C528 source.n398 a_n2210_n3288# 0.014107f
C529 source.n399 a_n2210_n3288# 0.031492f
C530 source.n400 a_n2210_n3288# 0.031492f
C531 source.n401 a_n2210_n3288# 0.014107f
C532 source.n402 a_n2210_n3288# 0.013323f
C533 source.n403 a_n2210_n3288# 0.024794f
C534 source.n404 a_n2210_n3288# 0.024794f
C535 source.n405 a_n2210_n3288# 0.013323f
C536 source.n406 a_n2210_n3288# 0.014107f
C537 source.n407 a_n2210_n3288# 0.031492f
C538 source.n408 a_n2210_n3288# 0.064624f
C539 source.n409 a_n2210_n3288# 0.014107f
C540 source.n410 a_n2210_n3288# 0.013323f
C541 source.n411 a_n2210_n3288# 0.053246f
C542 source.n412 a_n2210_n3288# 0.035666f
C543 source.n413 a_n2210_n3288# 0.113587f
C544 source.n414 a_n2210_n3288# 0.032843f
C545 source.n415 a_n2210_n3288# 0.024794f
C546 source.n416 a_n2210_n3288# 0.013323f
C547 source.n417 a_n2210_n3288# 0.031492f
C548 source.n418 a_n2210_n3288# 0.014107f
C549 source.n419 a_n2210_n3288# 0.024794f
C550 source.n420 a_n2210_n3288# 0.013323f
C551 source.n421 a_n2210_n3288# 0.031492f
C552 source.n422 a_n2210_n3288# 0.014107f
C553 source.n423 a_n2210_n3288# 0.024794f
C554 source.n424 a_n2210_n3288# 0.013715f
C555 source.n425 a_n2210_n3288# 0.031492f
C556 source.n426 a_n2210_n3288# 0.014107f
C557 source.n427 a_n2210_n3288# 0.024794f
C558 source.n428 a_n2210_n3288# 0.013323f
C559 source.n429 a_n2210_n3288# 0.031492f
C560 source.n430 a_n2210_n3288# 0.014107f
C561 source.n431 a_n2210_n3288# 0.024794f
C562 source.n432 a_n2210_n3288# 0.013323f
C563 source.n433 a_n2210_n3288# 0.023619f
C564 source.n434 a_n2210_n3288# 0.022262f
C565 source.t6 a_n2210_n3288# 0.053187f
C566 source.n435 a_n2210_n3288# 0.178764f
C567 source.n436 a_n2210_n3288# 1.25083f
C568 source.n437 a_n2210_n3288# 0.013323f
C569 source.n438 a_n2210_n3288# 0.014107f
C570 source.n439 a_n2210_n3288# 0.031492f
C571 source.n440 a_n2210_n3288# 0.031492f
C572 source.n441 a_n2210_n3288# 0.014107f
C573 source.n442 a_n2210_n3288# 0.013323f
C574 source.n443 a_n2210_n3288# 0.024794f
C575 source.n444 a_n2210_n3288# 0.024794f
C576 source.n445 a_n2210_n3288# 0.013323f
C577 source.n446 a_n2210_n3288# 0.014107f
C578 source.n447 a_n2210_n3288# 0.031492f
C579 source.n448 a_n2210_n3288# 0.031492f
C580 source.n449 a_n2210_n3288# 0.014107f
C581 source.n450 a_n2210_n3288# 0.013323f
C582 source.n451 a_n2210_n3288# 0.024794f
C583 source.n452 a_n2210_n3288# 0.024794f
C584 source.n453 a_n2210_n3288# 0.013323f
C585 source.n454 a_n2210_n3288# 0.013323f
C586 source.n455 a_n2210_n3288# 0.014107f
C587 source.n456 a_n2210_n3288# 0.031492f
C588 source.n457 a_n2210_n3288# 0.031492f
C589 source.n458 a_n2210_n3288# 0.031492f
C590 source.n459 a_n2210_n3288# 0.013715f
C591 source.n460 a_n2210_n3288# 0.013323f
C592 source.n461 a_n2210_n3288# 0.024794f
C593 source.n462 a_n2210_n3288# 0.024794f
C594 source.n463 a_n2210_n3288# 0.013323f
C595 source.n464 a_n2210_n3288# 0.014107f
C596 source.n465 a_n2210_n3288# 0.031492f
C597 source.n466 a_n2210_n3288# 0.031492f
C598 source.n467 a_n2210_n3288# 0.014107f
C599 source.n468 a_n2210_n3288# 0.013323f
C600 source.n469 a_n2210_n3288# 0.024794f
C601 source.n470 a_n2210_n3288# 0.024794f
C602 source.n471 a_n2210_n3288# 0.013323f
C603 source.n472 a_n2210_n3288# 0.014107f
C604 source.n473 a_n2210_n3288# 0.031492f
C605 source.n474 a_n2210_n3288# 0.064624f
C606 source.n475 a_n2210_n3288# 0.014107f
C607 source.n476 a_n2210_n3288# 0.013323f
C608 source.n477 a_n2210_n3288# 0.053246f
C609 source.n478 a_n2210_n3288# 0.035666f
C610 source.n479 a_n2210_n3288# 0.113587f
C611 source.t9 a_n2210_n3288# 0.235119f
C612 source.t11 a_n2210_n3288# 0.235119f
C613 source.n480 a_n2210_n3288# 2.01308f
C614 source.n481 a_n2210_n3288# 0.367832f
C615 source.t3 a_n2210_n3288# 0.235119f
C616 source.t10 a_n2210_n3288# 0.235119f
C617 source.n482 a_n2210_n3288# 2.01308f
C618 source.n483 a_n2210_n3288# 0.367832f
C619 source.t0 a_n2210_n3288# 0.235119f
C620 source.t12 a_n2210_n3288# 0.235119f
C621 source.n484 a_n2210_n3288# 2.01308f
C622 source.n485 a_n2210_n3288# 0.367832f
C623 source.n486 a_n2210_n3288# 0.032843f
C624 source.n487 a_n2210_n3288# 0.024794f
C625 source.n488 a_n2210_n3288# 0.013323f
C626 source.n489 a_n2210_n3288# 0.031492f
C627 source.n490 a_n2210_n3288# 0.014107f
C628 source.n491 a_n2210_n3288# 0.024794f
C629 source.n492 a_n2210_n3288# 0.013323f
C630 source.n493 a_n2210_n3288# 0.031492f
C631 source.n494 a_n2210_n3288# 0.014107f
C632 source.n495 a_n2210_n3288# 0.024794f
C633 source.n496 a_n2210_n3288# 0.013715f
C634 source.n497 a_n2210_n3288# 0.031492f
C635 source.n498 a_n2210_n3288# 0.014107f
C636 source.n499 a_n2210_n3288# 0.024794f
C637 source.n500 a_n2210_n3288# 0.013323f
C638 source.n501 a_n2210_n3288# 0.031492f
C639 source.n502 a_n2210_n3288# 0.014107f
C640 source.n503 a_n2210_n3288# 0.024794f
C641 source.n504 a_n2210_n3288# 0.013323f
C642 source.n505 a_n2210_n3288# 0.023619f
C643 source.n506 a_n2210_n3288# 0.022262f
C644 source.t15 a_n2210_n3288# 0.053187f
C645 source.n507 a_n2210_n3288# 0.178764f
C646 source.n508 a_n2210_n3288# 1.25083f
C647 source.n509 a_n2210_n3288# 0.013323f
C648 source.n510 a_n2210_n3288# 0.014107f
C649 source.n511 a_n2210_n3288# 0.031492f
C650 source.n512 a_n2210_n3288# 0.031492f
C651 source.n513 a_n2210_n3288# 0.014107f
C652 source.n514 a_n2210_n3288# 0.013323f
C653 source.n515 a_n2210_n3288# 0.024794f
C654 source.n516 a_n2210_n3288# 0.024794f
C655 source.n517 a_n2210_n3288# 0.013323f
C656 source.n518 a_n2210_n3288# 0.014107f
C657 source.n519 a_n2210_n3288# 0.031492f
C658 source.n520 a_n2210_n3288# 0.031492f
C659 source.n521 a_n2210_n3288# 0.014107f
C660 source.n522 a_n2210_n3288# 0.013323f
C661 source.n523 a_n2210_n3288# 0.024794f
C662 source.n524 a_n2210_n3288# 0.024794f
C663 source.n525 a_n2210_n3288# 0.013323f
C664 source.n526 a_n2210_n3288# 0.013323f
C665 source.n527 a_n2210_n3288# 0.014107f
C666 source.n528 a_n2210_n3288# 0.031492f
C667 source.n529 a_n2210_n3288# 0.031492f
C668 source.n530 a_n2210_n3288# 0.031492f
C669 source.n531 a_n2210_n3288# 0.013715f
C670 source.n532 a_n2210_n3288# 0.013323f
C671 source.n533 a_n2210_n3288# 0.024794f
C672 source.n534 a_n2210_n3288# 0.024794f
C673 source.n535 a_n2210_n3288# 0.013323f
C674 source.n536 a_n2210_n3288# 0.014107f
C675 source.n537 a_n2210_n3288# 0.031492f
C676 source.n538 a_n2210_n3288# 0.031492f
C677 source.n539 a_n2210_n3288# 0.014107f
C678 source.n540 a_n2210_n3288# 0.013323f
C679 source.n541 a_n2210_n3288# 0.024794f
C680 source.n542 a_n2210_n3288# 0.024794f
C681 source.n543 a_n2210_n3288# 0.013323f
C682 source.n544 a_n2210_n3288# 0.014107f
C683 source.n545 a_n2210_n3288# 0.031492f
C684 source.n546 a_n2210_n3288# 0.064624f
C685 source.n547 a_n2210_n3288# 0.014107f
C686 source.n548 a_n2210_n3288# 0.013323f
C687 source.n549 a_n2210_n3288# 0.053246f
C688 source.n550 a_n2210_n3288# 0.035666f
C689 source.n551 a_n2210_n3288# 0.264498f
C690 source.n552 a_n2210_n3288# 1.56323f
C691 drain_left.t7 a_n2210_n3288# 0.278276f
C692 drain_left.t4 a_n2210_n3288# 0.278276f
C693 drain_left.n0 a_n2210_n3288# 2.4809f
C694 drain_left.t11 a_n2210_n3288# 0.278276f
C695 drain_left.t15 a_n2210_n3288# 0.278276f
C696 drain_left.n1 a_n2210_n3288# 2.47622f
C697 drain_left.n2 a_n2210_n3288# 0.733533f
C698 drain_left.t1 a_n2210_n3288# 0.278276f
C699 drain_left.t0 a_n2210_n3288# 0.278276f
C700 drain_left.n3 a_n2210_n3288# 2.4809f
C701 drain_left.t10 a_n2210_n3288# 0.278276f
C702 drain_left.t13 a_n2210_n3288# 0.278276f
C703 drain_left.n4 a_n2210_n3288# 2.47622f
C704 drain_left.n5 a_n2210_n3288# 0.733533f
C705 drain_left.n6 a_n2210_n3288# 1.56219f
C706 drain_left.t12 a_n2210_n3288# 0.278276f
C707 drain_left.t9 a_n2210_n3288# 0.278276f
C708 drain_left.n7 a_n2210_n3288# 2.48091f
C709 drain_left.t2 a_n2210_n3288# 0.278276f
C710 drain_left.t14 a_n2210_n3288# 0.278276f
C711 drain_left.n8 a_n2210_n3288# 2.47623f
C712 drain_left.n9 a_n2210_n3288# 0.770325f
C713 drain_left.t8 a_n2210_n3288# 0.278276f
C714 drain_left.t3 a_n2210_n3288# 0.278276f
C715 drain_left.n10 a_n2210_n3288# 2.47623f
C716 drain_left.n11 a_n2210_n3288# 0.381588f
C717 drain_left.t5 a_n2210_n3288# 0.278276f
C718 drain_left.t6 a_n2210_n3288# 0.278276f
C719 drain_left.n12 a_n2210_n3288# 2.47622f
C720 drain_left.n13 a_n2210_n3288# 0.633717f
C721 plus.n0 a_n2210_n3288# 0.045852f
C722 plus.t12 a_n2210_n3288# 0.784492f
C723 plus.t7 a_n2210_n3288# 0.784492f
C724 plus.t15 a_n2210_n3288# 0.784492f
C725 plus.n1 a_n2210_n3288# 0.321255f
C726 plus.n2 a_n2210_n3288# 0.045852f
C727 plus.t9 a_n2210_n3288# 0.784492f
C728 plus.t5 a_n2210_n3288# 0.784492f
C729 plus.n3 a_n2210_n3288# 0.045852f
C730 plus.t13 a_n2210_n3288# 0.784492f
C731 plus.n4 a_n2210_n3288# 0.321255f
C732 plus.t2 a_n2210_n3288# 0.794287f
C733 plus.n5 a_n2210_n3288# 0.306987f
C734 plus.t8 a_n2210_n3288# 0.784492f
C735 plus.n6 a_n2210_n3288# 0.318569f
C736 plus.n7 a_n2210_n3288# 0.010405f
C737 plus.n8 a_n2210_n3288# 0.145987f
C738 plus.n9 a_n2210_n3288# 0.045852f
C739 plus.n10 a_n2210_n3288# 0.045852f
C740 plus.n11 a_n2210_n3288# 0.010405f
C741 plus.n12 a_n2210_n3288# 0.318852f
C742 plus.n13 a_n2210_n3288# 0.318852f
C743 plus.n14 a_n2210_n3288# 0.010405f
C744 plus.n15 a_n2210_n3288# 0.045852f
C745 plus.n16 a_n2210_n3288# 0.045852f
C746 plus.n17 a_n2210_n3288# 0.045852f
C747 plus.n18 a_n2210_n3288# 0.010405f
C748 plus.n19 a_n2210_n3288# 0.318569f
C749 plus.n20 a_n2210_n3288# 0.316449f
C750 plus.n21 a_n2210_n3288# 0.519707f
C751 plus.n22 a_n2210_n3288# 0.045852f
C752 plus.t14 a_n2210_n3288# 0.784492f
C753 plus.t3 a_n2210_n3288# 0.784492f
C754 plus.t6 a_n2210_n3288# 0.784492f
C755 plus.n23 a_n2210_n3288# 0.321255f
C756 plus.n24 a_n2210_n3288# 0.045852f
C757 plus.t1 a_n2210_n3288# 0.784492f
C758 plus.n25 a_n2210_n3288# 0.045852f
C759 plus.t0 a_n2210_n3288# 0.784492f
C760 plus.t4 a_n2210_n3288# 0.784492f
C761 plus.n26 a_n2210_n3288# 0.321255f
C762 plus.t10 a_n2210_n3288# 0.794287f
C763 plus.n27 a_n2210_n3288# 0.306987f
C764 plus.t11 a_n2210_n3288# 0.784492f
C765 plus.n28 a_n2210_n3288# 0.318569f
C766 plus.n29 a_n2210_n3288# 0.010405f
C767 plus.n30 a_n2210_n3288# 0.145987f
C768 plus.n31 a_n2210_n3288# 0.045852f
C769 plus.n32 a_n2210_n3288# 0.045852f
C770 plus.n33 a_n2210_n3288# 0.010405f
C771 plus.n34 a_n2210_n3288# 0.318852f
C772 plus.n35 a_n2210_n3288# 0.318852f
C773 plus.n36 a_n2210_n3288# 0.010405f
C774 plus.n37 a_n2210_n3288# 0.045852f
C775 plus.n38 a_n2210_n3288# 0.045852f
C776 plus.n39 a_n2210_n3288# 0.045852f
C777 plus.n40 a_n2210_n3288# 0.010405f
C778 plus.n41 a_n2210_n3288# 0.318569f
C779 plus.n42 a_n2210_n3288# 0.316449f
C780 plus.n43 a_n2210_n3288# 1.45825f
.ends

