* NGSPICE file created from diffpair579.ext - technology: sky130A

.subckt diffpair579 minus drain_right drain_left source plus
X0 drain_left.t23 plus.t0 source.t32 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X1 drain_left.t22 plus.t1 source.t28 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X2 source.t31 plus.t2 drain_left.t21 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X3 drain_right.t23 minus.t0 source.t22 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X4 drain_right.t22 minus.t1 source.t21 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X5 source.t30 plus.t3 drain_left.t20 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X6 a_n2094_n4888# a_n2094_n4888# a_n2094_n4888# a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.2
X7 source.t16 minus.t2 drain_right.t21 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X8 a_n2094_n4888# a_n2094_n4888# a_n2094_n4888# a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X9 source.t44 plus.t4 drain_left.t19 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X10 drain_left.t18 plus.t5 source.t46 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X11 source.t15 minus.t3 drain_right.t20 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X12 source.t20 minus.t4 drain_right.t19 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X13 source.t17 minus.t5 drain_right.t18 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X14 source.t8 minus.t6 drain_right.t17 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X15 source.t11 minus.t7 drain_right.t16 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X16 drain_left.t17 plus.t6 source.t45 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X17 drain_right.t15 minus.t8 source.t0 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X18 drain_right.t14 minus.t9 source.t1 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X19 source.t4 minus.t10 drain_right.t13 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X20 drain_right.t12 minus.t11 source.t7 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X21 drain_right.t11 minus.t12 source.t10 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X22 drain_right.t10 minus.t13 source.t5 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X23 drain_left.t16 plus.t7 source.t47 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X24 source.t29 plus.t8 drain_left.t15 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X25 a_n2094_n4888# a_n2094_n4888# a_n2094_n4888# a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X26 drain_right.t9 minus.t14 source.t13 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X27 drain_right.t8 minus.t15 source.t6 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X28 source.t18 minus.t16 drain_right.t7 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X29 drain_right.t6 minus.t17 source.t23 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X30 source.t12 minus.t18 drain_right.t5 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X31 source.t40 plus.t9 drain_left.t14 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X32 drain_right.t4 minus.t19 source.t2 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X33 drain_right.t3 minus.t20 source.t3 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X34 source.t9 minus.t21 drain_right.t2 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X35 drain_left.t13 plus.t10 source.t38 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X36 source.t36 plus.t11 drain_left.t12 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X37 a_n2094_n4888# a_n2094_n4888# a_n2094_n4888# a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X38 source.t34 plus.t12 drain_left.t11 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X39 drain_left.t10 plus.t13 source.t27 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X40 drain_left.t9 plus.t14 source.t43 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X41 source.t24 plus.t15 drain_left.t8 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X42 source.t14 minus.t22 drain_right.t1 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X43 source.t19 minus.t23 drain_right.t0 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X44 source.t26 plus.t16 drain_left.t7 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X45 source.t39 plus.t17 drain_left.t6 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X46 drain_left.t5 plus.t18 source.t37 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X47 source.t35 plus.t19 drain_left.t4 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X48 drain_left.t3 plus.t20 source.t33 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X49 drain_left.t2 plus.t21 source.t42 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X50 source.t25 plus.t22 drain_left.t1 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X51 drain_left.t0 plus.t23 source.t41 a_n2094_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
R0 plus.n6 plus.t8 2627.27
R1 plus.n29 plus.t18 2627.27
R2 plus.n37 plus.t0 2627.27
R3 plus.n60 plus.t19 2627.27
R4 plus.n7 plus.t5 2566.65
R5 plus.n5 plus.t22 2566.65
R6 plus.n12 plus.t13 2566.65
R7 plus.n14 plus.t12 2566.65
R8 plus.n3 plus.t7 2566.65
R9 plus.n19 plus.t4 2566.65
R10 plus.n21 plus.t21 2566.65
R11 plus.n1 plus.t11 2566.65
R12 plus.n26 plus.t6 2566.65
R13 plus.n28 plus.t2 2566.65
R14 plus.n38 plus.t3 2566.65
R15 plus.n36 plus.t1 2566.65
R16 plus.n43 plus.t16 2566.65
R17 plus.n45 plus.t23 2566.65
R18 plus.n34 plus.t17 2566.65
R19 plus.n50 plus.t20 2566.65
R20 plus.n52 plus.t15 2566.65
R21 plus.n32 plus.t10 2566.65
R22 plus.n57 plus.t9 2566.65
R23 plus.n59 plus.t14 2566.65
R24 plus.n9 plus.n6 161.489
R25 plus.n40 plus.n37 161.489
R26 plus.n9 plus.n8 161.3
R27 plus.n11 plus.n10 161.3
R28 plus.n13 plus.n4 161.3
R29 plus.n16 plus.n15 161.3
R30 plus.n18 plus.n17 161.3
R31 plus.n20 plus.n2 161.3
R32 plus.n23 plus.n22 161.3
R33 plus.n25 plus.n24 161.3
R34 plus.n27 plus.n0 161.3
R35 plus.n30 plus.n29 161.3
R36 plus.n40 plus.n39 161.3
R37 plus.n42 plus.n41 161.3
R38 plus.n44 plus.n35 161.3
R39 plus.n47 plus.n46 161.3
R40 plus.n49 plus.n48 161.3
R41 plus.n51 plus.n33 161.3
R42 plus.n54 plus.n53 161.3
R43 plus.n56 plus.n55 161.3
R44 plus.n58 plus.n31 161.3
R45 plus.n61 plus.n60 161.3
R46 plus.n8 plus.n7 56.2338
R47 plus.n28 plus.n27 56.2338
R48 plus.n59 plus.n58 56.2338
R49 plus.n39 plus.n38 56.2338
R50 plus.n11 plus.n5 51.852
R51 plus.n26 plus.n25 51.852
R52 plus.n57 plus.n56 51.852
R53 plus.n42 plus.n36 51.852
R54 plus.n13 plus.n12 47.4702
R55 plus.n22 plus.n1 47.4702
R56 plus.n53 plus.n32 47.4702
R57 plus.n44 plus.n43 47.4702
R58 plus.n15 plus.n14 43.0884
R59 plus.n21 plus.n20 43.0884
R60 plus.n52 plus.n51 43.0884
R61 plus.n46 plus.n45 43.0884
R62 plus.n18 plus.n3 38.7066
R63 plus.n19 plus.n18 38.7066
R64 plus.n50 plus.n49 38.7066
R65 plus.n49 plus.n34 38.7066
R66 plus.n15 plus.n3 34.3247
R67 plus.n20 plus.n19 34.3247
R68 plus.n51 plus.n50 34.3247
R69 plus.n46 plus.n34 34.3247
R70 plus plus.n61 33.9536
R71 plus.n14 plus.n13 29.9429
R72 plus.n22 plus.n21 29.9429
R73 plus.n53 plus.n52 29.9429
R74 plus.n45 plus.n44 29.9429
R75 plus.n12 plus.n11 25.5611
R76 plus.n25 plus.n1 25.5611
R77 plus.n56 plus.n32 25.5611
R78 plus.n43 plus.n42 25.5611
R79 plus.n8 plus.n5 21.1793
R80 plus.n27 plus.n26 21.1793
R81 plus.n58 plus.n57 21.1793
R82 plus.n39 plus.n36 21.1793
R83 plus.n7 plus.n6 16.7975
R84 plus.n29 plus.n28 16.7975
R85 plus.n60 plus.n59 16.7975
R86 plus.n38 plus.n37 16.7975
R87 plus plus.n30 15.1634
R88 plus.n10 plus.n9 0.189894
R89 plus.n10 plus.n4 0.189894
R90 plus.n16 plus.n4 0.189894
R91 plus.n17 plus.n16 0.189894
R92 plus.n17 plus.n2 0.189894
R93 plus.n23 plus.n2 0.189894
R94 plus.n24 plus.n23 0.189894
R95 plus.n24 plus.n0 0.189894
R96 plus.n30 plus.n0 0.189894
R97 plus.n61 plus.n31 0.189894
R98 plus.n55 plus.n31 0.189894
R99 plus.n55 plus.n54 0.189894
R100 plus.n54 plus.n33 0.189894
R101 plus.n48 plus.n33 0.189894
R102 plus.n48 plus.n47 0.189894
R103 plus.n47 plus.n35 0.189894
R104 plus.n41 plus.n35 0.189894
R105 plus.n41 plus.n40 0.189894
R106 source.n0 source.t37 44.1297
R107 source.n11 source.t29 44.1296
R108 source.n12 source.t2 44.1296
R109 source.n23 source.t16 44.1296
R110 source.n47 source.t0 44.1295
R111 source.n36 source.t8 44.1295
R112 source.n35 source.t32 44.1295
R113 source.n24 source.t35 44.1295
R114 source.n2 source.n1 43.1397
R115 source.n4 source.n3 43.1397
R116 source.n6 source.n5 43.1397
R117 source.n8 source.n7 43.1397
R118 source.n10 source.n9 43.1397
R119 source.n14 source.n13 43.1397
R120 source.n16 source.n15 43.1397
R121 source.n18 source.n17 43.1397
R122 source.n20 source.n19 43.1397
R123 source.n22 source.n21 43.1397
R124 source.n46 source.n45 43.1396
R125 source.n44 source.n43 43.1396
R126 source.n42 source.n41 43.1396
R127 source.n40 source.n39 43.1396
R128 source.n38 source.n37 43.1396
R129 source.n34 source.n33 43.1396
R130 source.n32 source.n31 43.1396
R131 source.n30 source.n29 43.1396
R132 source.n28 source.n27 43.1396
R133 source.n26 source.n25 43.1396
R134 source.n24 source.n23 27.8052
R135 source.n48 source.n0 22.3138
R136 source.n48 source.n47 5.49188
R137 source.n45 source.t1 0.9905
R138 source.n45 source.t15 0.9905
R139 source.n43 source.t13 0.9905
R140 source.n43 source.t18 0.9905
R141 source.n41 source.t6 0.9905
R142 source.n41 source.t12 0.9905
R143 source.n39 source.t10 0.9905
R144 source.n39 source.t9 0.9905
R145 source.n37 source.t5 0.9905
R146 source.n37 source.t20 0.9905
R147 source.n33 source.t28 0.9905
R148 source.n33 source.t30 0.9905
R149 source.n31 source.t41 0.9905
R150 source.n31 source.t26 0.9905
R151 source.n29 source.t33 0.9905
R152 source.n29 source.t39 0.9905
R153 source.n27 source.t38 0.9905
R154 source.n27 source.t24 0.9905
R155 source.n25 source.t43 0.9905
R156 source.n25 source.t40 0.9905
R157 source.n1 source.t45 0.9905
R158 source.n1 source.t31 0.9905
R159 source.n3 source.t42 0.9905
R160 source.n3 source.t36 0.9905
R161 source.n5 source.t47 0.9905
R162 source.n5 source.t44 0.9905
R163 source.n7 source.t27 0.9905
R164 source.n7 source.t34 0.9905
R165 source.n9 source.t46 0.9905
R166 source.n9 source.t25 0.9905
R167 source.n13 source.t22 0.9905
R168 source.n13 source.t11 0.9905
R169 source.n15 source.t3 0.9905
R170 source.n15 source.t14 0.9905
R171 source.n17 source.t21 0.9905
R172 source.n17 source.t17 0.9905
R173 source.n19 source.t23 0.9905
R174 source.n19 source.t19 0.9905
R175 source.n21 source.t7 0.9905
R176 source.n21 source.t4 0.9905
R177 source.n12 source.n11 0.470328
R178 source.n36 source.n35 0.470328
R179 source.n23 source.n22 0.457397
R180 source.n22 source.n20 0.457397
R181 source.n20 source.n18 0.457397
R182 source.n18 source.n16 0.457397
R183 source.n16 source.n14 0.457397
R184 source.n14 source.n12 0.457397
R185 source.n11 source.n10 0.457397
R186 source.n10 source.n8 0.457397
R187 source.n8 source.n6 0.457397
R188 source.n6 source.n4 0.457397
R189 source.n4 source.n2 0.457397
R190 source.n2 source.n0 0.457397
R191 source.n26 source.n24 0.457397
R192 source.n28 source.n26 0.457397
R193 source.n30 source.n28 0.457397
R194 source.n32 source.n30 0.457397
R195 source.n34 source.n32 0.457397
R196 source.n35 source.n34 0.457397
R197 source.n38 source.n36 0.457397
R198 source.n40 source.n38 0.457397
R199 source.n42 source.n40 0.457397
R200 source.n44 source.n42 0.457397
R201 source.n46 source.n44 0.457397
R202 source.n47 source.n46 0.457397
R203 source source.n48 0.188
R204 drain_left.n13 drain_left.n11 60.2753
R205 drain_left.n7 drain_left.n5 60.2753
R206 drain_left.n2 drain_left.n0 60.2753
R207 drain_left.n21 drain_left.n20 59.8185
R208 drain_left.n19 drain_left.n18 59.8185
R209 drain_left.n17 drain_left.n16 59.8185
R210 drain_left.n15 drain_left.n14 59.8185
R211 drain_left.n13 drain_left.n12 59.8185
R212 drain_left.n7 drain_left.n6 59.8184
R213 drain_left.n9 drain_left.n8 59.8184
R214 drain_left.n4 drain_left.n3 59.8184
R215 drain_left.n2 drain_left.n1 59.8184
R216 drain_left drain_left.n10 37.7682
R217 drain_left drain_left.n21 6.11011
R218 drain_left.n5 drain_left.t20 0.9905
R219 drain_left.n5 drain_left.t23 0.9905
R220 drain_left.n6 drain_left.t7 0.9905
R221 drain_left.n6 drain_left.t22 0.9905
R222 drain_left.n8 drain_left.t6 0.9905
R223 drain_left.n8 drain_left.t0 0.9905
R224 drain_left.n3 drain_left.t8 0.9905
R225 drain_left.n3 drain_left.t3 0.9905
R226 drain_left.n1 drain_left.t14 0.9905
R227 drain_left.n1 drain_left.t13 0.9905
R228 drain_left.n0 drain_left.t4 0.9905
R229 drain_left.n0 drain_left.t9 0.9905
R230 drain_left.n20 drain_left.t21 0.9905
R231 drain_left.n20 drain_left.t5 0.9905
R232 drain_left.n18 drain_left.t12 0.9905
R233 drain_left.n18 drain_left.t17 0.9905
R234 drain_left.n16 drain_left.t19 0.9905
R235 drain_left.n16 drain_left.t2 0.9905
R236 drain_left.n14 drain_left.t11 0.9905
R237 drain_left.n14 drain_left.t16 0.9905
R238 drain_left.n12 drain_left.t1 0.9905
R239 drain_left.n12 drain_left.t10 0.9905
R240 drain_left.n11 drain_left.t15 0.9905
R241 drain_left.n11 drain_left.t18 0.9905
R242 drain_left.n9 drain_left.n7 0.457397
R243 drain_left.n4 drain_left.n2 0.457397
R244 drain_left.n15 drain_left.n13 0.457397
R245 drain_left.n17 drain_left.n15 0.457397
R246 drain_left.n19 drain_left.n17 0.457397
R247 drain_left.n21 drain_left.n19 0.457397
R248 drain_left.n10 drain_left.n9 0.173602
R249 drain_left.n10 drain_left.n4 0.173602
R250 minus.n29 minus.t2 2627.27
R251 minus.n6 minus.t19 2627.27
R252 minus.n60 minus.t8 2627.27
R253 minus.n37 minus.t6 2627.27
R254 minus.n28 minus.t11 2566.65
R255 minus.n26 minus.t10 2566.65
R256 minus.n1 minus.t17 2566.65
R257 minus.n21 minus.t23 2566.65
R258 minus.n19 minus.t1 2566.65
R259 minus.n3 minus.t5 2566.65
R260 minus.n14 minus.t20 2566.65
R261 minus.n12 minus.t22 2566.65
R262 minus.n5 minus.t0 2566.65
R263 minus.n7 minus.t7 2566.65
R264 minus.n59 minus.t3 2566.65
R265 minus.n57 minus.t9 2566.65
R266 minus.n32 minus.t16 2566.65
R267 minus.n52 minus.t14 2566.65
R268 minus.n50 minus.t18 2566.65
R269 minus.n34 minus.t15 2566.65
R270 minus.n45 minus.t21 2566.65
R271 minus.n43 minus.t12 2566.65
R272 minus.n36 minus.t4 2566.65
R273 minus.n38 minus.t13 2566.65
R274 minus.n9 minus.n6 161.489
R275 minus.n40 minus.n37 161.489
R276 minus.n30 minus.n29 161.3
R277 minus.n27 minus.n0 161.3
R278 minus.n25 minus.n24 161.3
R279 minus.n23 minus.n22 161.3
R280 minus.n20 minus.n2 161.3
R281 minus.n18 minus.n17 161.3
R282 minus.n16 minus.n15 161.3
R283 minus.n13 minus.n4 161.3
R284 minus.n11 minus.n10 161.3
R285 minus.n9 minus.n8 161.3
R286 minus.n61 minus.n60 161.3
R287 minus.n58 minus.n31 161.3
R288 minus.n56 minus.n55 161.3
R289 minus.n54 minus.n53 161.3
R290 minus.n51 minus.n33 161.3
R291 minus.n49 minus.n48 161.3
R292 minus.n47 minus.n46 161.3
R293 minus.n44 minus.n35 161.3
R294 minus.n42 minus.n41 161.3
R295 minus.n40 minus.n39 161.3
R296 minus.n28 minus.n27 56.2338
R297 minus.n8 minus.n7 56.2338
R298 minus.n39 minus.n38 56.2338
R299 minus.n59 minus.n58 56.2338
R300 minus.n26 minus.n25 51.852
R301 minus.n11 minus.n5 51.852
R302 minus.n42 minus.n36 51.852
R303 minus.n57 minus.n56 51.852
R304 minus.n22 minus.n1 47.4702
R305 minus.n13 minus.n12 47.4702
R306 minus.n44 minus.n43 47.4702
R307 minus.n53 minus.n32 47.4702
R308 minus.n62 minus.n30 43.1028
R309 minus.n21 minus.n20 43.0884
R310 minus.n15 minus.n14 43.0884
R311 minus.n46 minus.n45 43.0884
R312 minus.n52 minus.n51 43.0884
R313 minus.n19 minus.n18 38.7066
R314 minus.n18 minus.n3 38.7066
R315 minus.n49 minus.n34 38.7066
R316 minus.n50 minus.n49 38.7066
R317 minus.n20 minus.n19 34.3247
R318 minus.n15 minus.n3 34.3247
R319 minus.n46 minus.n34 34.3247
R320 minus.n51 minus.n50 34.3247
R321 minus.n22 minus.n21 29.9429
R322 minus.n14 minus.n13 29.9429
R323 minus.n45 minus.n44 29.9429
R324 minus.n53 minus.n52 29.9429
R325 minus.n25 minus.n1 25.5611
R326 minus.n12 minus.n11 25.5611
R327 minus.n43 minus.n42 25.5611
R328 minus.n56 minus.n32 25.5611
R329 minus.n27 minus.n26 21.1793
R330 minus.n8 minus.n5 21.1793
R331 minus.n39 minus.n36 21.1793
R332 minus.n58 minus.n57 21.1793
R333 minus.n29 minus.n28 16.7975
R334 minus.n7 minus.n6 16.7975
R335 minus.n38 minus.n37 16.7975
R336 minus.n60 minus.n59 16.7975
R337 minus.n62 minus.n61 6.48914
R338 minus.n30 minus.n0 0.189894
R339 minus.n24 minus.n0 0.189894
R340 minus.n24 minus.n23 0.189894
R341 minus.n23 minus.n2 0.189894
R342 minus.n17 minus.n2 0.189894
R343 minus.n17 minus.n16 0.189894
R344 minus.n16 minus.n4 0.189894
R345 minus.n10 minus.n4 0.189894
R346 minus.n10 minus.n9 0.189894
R347 minus.n41 minus.n40 0.189894
R348 minus.n41 minus.n35 0.189894
R349 minus.n47 minus.n35 0.189894
R350 minus.n48 minus.n47 0.189894
R351 minus.n48 minus.n33 0.189894
R352 minus.n54 minus.n33 0.189894
R353 minus.n55 minus.n54 0.189894
R354 minus.n55 minus.n31 0.189894
R355 minus.n61 minus.n31 0.189894
R356 minus minus.n62 0.188
R357 drain_right.n13 drain_right.n11 60.2753
R358 drain_right.n7 drain_right.n5 60.2753
R359 drain_right.n2 drain_right.n0 60.2753
R360 drain_right.n13 drain_right.n12 59.8185
R361 drain_right.n15 drain_right.n14 59.8185
R362 drain_right.n17 drain_right.n16 59.8185
R363 drain_right.n19 drain_right.n18 59.8185
R364 drain_right.n21 drain_right.n20 59.8185
R365 drain_right.n7 drain_right.n6 59.8184
R366 drain_right.n9 drain_right.n8 59.8184
R367 drain_right.n4 drain_right.n3 59.8184
R368 drain_right.n2 drain_right.n1 59.8184
R369 drain_right drain_right.n10 37.215
R370 drain_right drain_right.n21 6.11011
R371 drain_right.n5 drain_right.t20 0.9905
R372 drain_right.n5 drain_right.t15 0.9905
R373 drain_right.n6 drain_right.t7 0.9905
R374 drain_right.n6 drain_right.t14 0.9905
R375 drain_right.n8 drain_right.t5 0.9905
R376 drain_right.n8 drain_right.t9 0.9905
R377 drain_right.n3 drain_right.t2 0.9905
R378 drain_right.n3 drain_right.t8 0.9905
R379 drain_right.n1 drain_right.t19 0.9905
R380 drain_right.n1 drain_right.t11 0.9905
R381 drain_right.n0 drain_right.t17 0.9905
R382 drain_right.n0 drain_right.t10 0.9905
R383 drain_right.n11 drain_right.t16 0.9905
R384 drain_right.n11 drain_right.t4 0.9905
R385 drain_right.n12 drain_right.t1 0.9905
R386 drain_right.n12 drain_right.t23 0.9905
R387 drain_right.n14 drain_right.t18 0.9905
R388 drain_right.n14 drain_right.t3 0.9905
R389 drain_right.n16 drain_right.t0 0.9905
R390 drain_right.n16 drain_right.t22 0.9905
R391 drain_right.n18 drain_right.t13 0.9905
R392 drain_right.n18 drain_right.t6 0.9905
R393 drain_right.n20 drain_right.t21 0.9905
R394 drain_right.n20 drain_right.t12 0.9905
R395 drain_right.n9 drain_right.n7 0.457397
R396 drain_right.n4 drain_right.n2 0.457397
R397 drain_right.n21 drain_right.n19 0.457397
R398 drain_right.n19 drain_right.n17 0.457397
R399 drain_right.n17 drain_right.n15 0.457397
R400 drain_right.n15 drain_right.n13 0.457397
R401 drain_right.n10 drain_right.n9 0.173602
R402 drain_right.n10 drain_right.n4 0.173602
C0 source minus 9.27291f
C1 plus drain_left 10.1416f
C2 drain_left drain_right 1.11966f
C3 plus minus 7.24759f
C4 minus drain_right 9.936501f
C5 plus source 9.28695f
C6 source drain_right 87.098f
C7 drain_left minus 0.171754f
C8 plus drain_right 0.359911f
C9 source drain_left 87.0977f
C10 drain_right a_n2094_n4888# 9.341461f
C11 drain_left a_n2094_n4888# 9.669019f
C12 source a_n2094_n4888# 12.903711f
C13 minus a_n2094_n4888# 8.689123f
C14 plus a_n2094_n4888# 11.337231f
C15 drain_right.t17 a_n2094_n4888# 0.624036f
C16 drain_right.t10 a_n2094_n4888# 0.624036f
C17 drain_right.n0 a_n2094_n4888# 5.7086f
C18 drain_right.t19 a_n2094_n4888# 0.624036f
C19 drain_right.t11 a_n2094_n4888# 0.624036f
C20 drain_right.n1 a_n2094_n4888# 5.70507f
C21 drain_right.n2 a_n2094_n4888# 0.91128f
C22 drain_right.t2 a_n2094_n4888# 0.624036f
C23 drain_right.t8 a_n2094_n4888# 0.624036f
C24 drain_right.n3 a_n2094_n4888# 5.70507f
C25 drain_right.n4 a_n2094_n4888# 0.418633f
C26 drain_right.t20 a_n2094_n4888# 0.624036f
C27 drain_right.t15 a_n2094_n4888# 0.624036f
C28 drain_right.n5 a_n2094_n4888# 5.7086f
C29 drain_right.t7 a_n2094_n4888# 0.624036f
C30 drain_right.t14 a_n2094_n4888# 0.624036f
C31 drain_right.n6 a_n2094_n4888# 5.70507f
C32 drain_right.n7 a_n2094_n4888# 0.91128f
C33 drain_right.t5 a_n2094_n4888# 0.624036f
C34 drain_right.t9 a_n2094_n4888# 0.624036f
C35 drain_right.n8 a_n2094_n4888# 5.70507f
C36 drain_right.n9 a_n2094_n4888# 0.418633f
C37 drain_right.n10 a_n2094_n4888# 2.71912f
C38 drain_right.t16 a_n2094_n4888# 0.624036f
C39 drain_right.t4 a_n2094_n4888# 0.624036f
C40 drain_right.n11 a_n2094_n4888# 5.70859f
C41 drain_right.t1 a_n2094_n4888# 0.624036f
C42 drain_right.t23 a_n2094_n4888# 0.624036f
C43 drain_right.n12 a_n2094_n4888# 5.70507f
C44 drain_right.n13 a_n2094_n4888# 0.911296f
C45 drain_right.t18 a_n2094_n4888# 0.624036f
C46 drain_right.t3 a_n2094_n4888# 0.624036f
C47 drain_right.n14 a_n2094_n4888# 5.70507f
C48 drain_right.n15 a_n2094_n4888# 0.44946f
C49 drain_right.t0 a_n2094_n4888# 0.624036f
C50 drain_right.t22 a_n2094_n4888# 0.624036f
C51 drain_right.n16 a_n2094_n4888# 5.70507f
C52 drain_right.n17 a_n2094_n4888# 0.44946f
C53 drain_right.t13 a_n2094_n4888# 0.624036f
C54 drain_right.t6 a_n2094_n4888# 0.624036f
C55 drain_right.n18 a_n2094_n4888# 5.70507f
C56 drain_right.n19 a_n2094_n4888# 0.44946f
C57 drain_right.t21 a_n2094_n4888# 0.624036f
C58 drain_right.t12 a_n2094_n4888# 0.624036f
C59 drain_right.n20 a_n2094_n4888# 5.70507f
C60 drain_right.n21 a_n2094_n4888# 0.772603f
C61 minus.n0 a_n2094_n4888# 0.05178f
C62 minus.t2 a_n2094_n4888# 0.588554f
C63 minus.t11 a_n2094_n4888# 0.583347f
C64 minus.t10 a_n2094_n4888# 0.583347f
C65 minus.t17 a_n2094_n4888# 0.583347f
C66 minus.n1 a_n2094_n4888# 0.22202f
C67 minus.n2 a_n2094_n4888# 0.05178f
C68 minus.t23 a_n2094_n4888# 0.583347f
C69 minus.t1 a_n2094_n4888# 0.583347f
C70 minus.t5 a_n2094_n4888# 0.583347f
C71 minus.n3 a_n2094_n4888# 0.22202f
C72 minus.n4 a_n2094_n4888# 0.05178f
C73 minus.t20 a_n2094_n4888# 0.583347f
C74 minus.t22 a_n2094_n4888# 0.583347f
C75 minus.t0 a_n2094_n4888# 0.583347f
C76 minus.n5 a_n2094_n4888# 0.22202f
C77 minus.t19 a_n2094_n4888# 0.588554f
C78 minus.n6 a_n2094_n4888# 0.2387f
C79 minus.t7 a_n2094_n4888# 0.583347f
C80 minus.n7 a_n2094_n4888# 0.22202f
C81 minus.n8 a_n2094_n4888# 0.018135f
C82 minus.n9 a_n2094_n4888# 0.120399f
C83 minus.n10 a_n2094_n4888# 0.05178f
C84 minus.n11 a_n2094_n4888# 0.018135f
C85 minus.n12 a_n2094_n4888# 0.22202f
C86 minus.n13 a_n2094_n4888# 0.018135f
C87 minus.n14 a_n2094_n4888# 0.22202f
C88 minus.n15 a_n2094_n4888# 0.018135f
C89 minus.n16 a_n2094_n4888# 0.05178f
C90 minus.n17 a_n2094_n4888# 0.05178f
C91 minus.n18 a_n2094_n4888# 0.018135f
C92 minus.n19 a_n2094_n4888# 0.22202f
C93 minus.n20 a_n2094_n4888# 0.018135f
C94 minus.n21 a_n2094_n4888# 0.22202f
C95 minus.n22 a_n2094_n4888# 0.018135f
C96 minus.n23 a_n2094_n4888# 0.05178f
C97 minus.n24 a_n2094_n4888# 0.05178f
C98 minus.n25 a_n2094_n4888# 0.018135f
C99 minus.n26 a_n2094_n4888# 0.22202f
C100 minus.n27 a_n2094_n4888# 0.018135f
C101 minus.n28 a_n2094_n4888# 0.22202f
C102 minus.n29 a_n2094_n4888# 0.238619f
C103 minus.n30 a_n2094_n4888# 2.38155f
C104 minus.n31 a_n2094_n4888# 0.05178f
C105 minus.t3 a_n2094_n4888# 0.583347f
C106 minus.t9 a_n2094_n4888# 0.583347f
C107 minus.t16 a_n2094_n4888# 0.583347f
C108 minus.n32 a_n2094_n4888# 0.22202f
C109 minus.n33 a_n2094_n4888# 0.05178f
C110 minus.t14 a_n2094_n4888# 0.583347f
C111 minus.t18 a_n2094_n4888# 0.583347f
C112 minus.t15 a_n2094_n4888# 0.583347f
C113 minus.n34 a_n2094_n4888# 0.22202f
C114 minus.n35 a_n2094_n4888# 0.05178f
C115 minus.t21 a_n2094_n4888# 0.583347f
C116 minus.t12 a_n2094_n4888# 0.583347f
C117 minus.t4 a_n2094_n4888# 0.583347f
C118 minus.n36 a_n2094_n4888# 0.22202f
C119 minus.t6 a_n2094_n4888# 0.588554f
C120 minus.n37 a_n2094_n4888# 0.2387f
C121 minus.t13 a_n2094_n4888# 0.583347f
C122 minus.n38 a_n2094_n4888# 0.22202f
C123 minus.n39 a_n2094_n4888# 0.018135f
C124 minus.n40 a_n2094_n4888# 0.120399f
C125 minus.n41 a_n2094_n4888# 0.05178f
C126 minus.n42 a_n2094_n4888# 0.018135f
C127 minus.n43 a_n2094_n4888# 0.22202f
C128 minus.n44 a_n2094_n4888# 0.018135f
C129 minus.n45 a_n2094_n4888# 0.22202f
C130 minus.n46 a_n2094_n4888# 0.018135f
C131 minus.n47 a_n2094_n4888# 0.05178f
C132 minus.n48 a_n2094_n4888# 0.05178f
C133 minus.n49 a_n2094_n4888# 0.018135f
C134 minus.n50 a_n2094_n4888# 0.22202f
C135 minus.n51 a_n2094_n4888# 0.018135f
C136 minus.n52 a_n2094_n4888# 0.22202f
C137 minus.n53 a_n2094_n4888# 0.018135f
C138 minus.n54 a_n2094_n4888# 0.05178f
C139 minus.n55 a_n2094_n4888# 0.05178f
C140 minus.n56 a_n2094_n4888# 0.018135f
C141 minus.n57 a_n2094_n4888# 0.22202f
C142 minus.n58 a_n2094_n4888# 0.018135f
C143 minus.n59 a_n2094_n4888# 0.22202f
C144 minus.t8 a_n2094_n4888# 0.588554f
C145 minus.n60 a_n2094_n4888# 0.238619f
C146 minus.n61 a_n2094_n4888# 0.337197f
C147 minus.n62 a_n2094_n4888# 2.83536f
C148 drain_left.t4 a_n2094_n4888# 0.624328f
C149 drain_left.t9 a_n2094_n4888# 0.624328f
C150 drain_left.n0 a_n2094_n4888# 5.71128f
C151 drain_left.t14 a_n2094_n4888# 0.624328f
C152 drain_left.t13 a_n2094_n4888# 0.624328f
C153 drain_left.n1 a_n2094_n4888# 5.70775f
C154 drain_left.n2 a_n2094_n4888# 0.911707f
C155 drain_left.t8 a_n2094_n4888# 0.624328f
C156 drain_left.t3 a_n2094_n4888# 0.624328f
C157 drain_left.n3 a_n2094_n4888# 5.70775f
C158 drain_left.n4 a_n2094_n4888# 0.41883f
C159 drain_left.t20 a_n2094_n4888# 0.624328f
C160 drain_left.t23 a_n2094_n4888# 0.624328f
C161 drain_left.n5 a_n2094_n4888# 5.71128f
C162 drain_left.t7 a_n2094_n4888# 0.624328f
C163 drain_left.t22 a_n2094_n4888# 0.624328f
C164 drain_left.n6 a_n2094_n4888# 5.70775f
C165 drain_left.n7 a_n2094_n4888# 0.911707f
C166 drain_left.t6 a_n2094_n4888# 0.624328f
C167 drain_left.t0 a_n2094_n4888# 0.624328f
C168 drain_left.n8 a_n2094_n4888# 5.70775f
C169 drain_left.n9 a_n2094_n4888# 0.41883f
C170 drain_left.n10 a_n2094_n4888# 2.80229f
C171 drain_left.t15 a_n2094_n4888# 0.624328f
C172 drain_left.t18 a_n2094_n4888# 0.624328f
C173 drain_left.n11 a_n2094_n4888# 5.71127f
C174 drain_left.t1 a_n2094_n4888# 0.624328f
C175 drain_left.t10 a_n2094_n4888# 0.624328f
C176 drain_left.n12 a_n2094_n4888# 5.70774f
C177 drain_left.n13 a_n2094_n4888# 0.911723f
C178 drain_left.t11 a_n2094_n4888# 0.624328f
C179 drain_left.t16 a_n2094_n4888# 0.624328f
C180 drain_left.n14 a_n2094_n4888# 5.70774f
C181 drain_left.n15 a_n2094_n4888# 0.449671f
C182 drain_left.t19 a_n2094_n4888# 0.624328f
C183 drain_left.t2 a_n2094_n4888# 0.624328f
C184 drain_left.n16 a_n2094_n4888# 5.70774f
C185 drain_left.n17 a_n2094_n4888# 0.449671f
C186 drain_left.t12 a_n2094_n4888# 0.624328f
C187 drain_left.t17 a_n2094_n4888# 0.624328f
C188 drain_left.n18 a_n2094_n4888# 5.70774f
C189 drain_left.n19 a_n2094_n4888# 0.449671f
C190 drain_left.t21 a_n2094_n4888# 0.624328f
C191 drain_left.t5 a_n2094_n4888# 0.624328f
C192 drain_left.n20 a_n2094_n4888# 5.70774f
C193 drain_left.n21 a_n2094_n4888# 0.772965f
C194 source.t37 a_n2094_n4888# 6.20311f
C195 source.n0 a_n2094_n4888# 2.62335f
C196 source.t45 a_n2094_n4888# 0.542781f
C197 source.t31 a_n2094_n4888# 0.542781f
C198 source.n1 a_n2094_n4888# 4.8527f
C199 source.n2 a_n2094_n4888# 0.453779f
C200 source.t42 a_n2094_n4888# 0.542781f
C201 source.t36 a_n2094_n4888# 0.542781f
C202 source.n3 a_n2094_n4888# 4.8527f
C203 source.n4 a_n2094_n4888# 0.453779f
C204 source.t47 a_n2094_n4888# 0.542781f
C205 source.t44 a_n2094_n4888# 0.542781f
C206 source.n5 a_n2094_n4888# 4.8527f
C207 source.n6 a_n2094_n4888# 0.453779f
C208 source.t27 a_n2094_n4888# 0.542781f
C209 source.t34 a_n2094_n4888# 0.542781f
C210 source.n7 a_n2094_n4888# 4.8527f
C211 source.n8 a_n2094_n4888# 0.453779f
C212 source.t46 a_n2094_n4888# 0.542781f
C213 source.t25 a_n2094_n4888# 0.542781f
C214 source.n9 a_n2094_n4888# 4.8527f
C215 source.n10 a_n2094_n4888# 0.453779f
C216 source.t29 a_n2094_n4888# 6.20312f
C217 source.n11 a_n2094_n4888# 0.585096f
C218 source.t2 a_n2094_n4888# 6.20312f
C219 source.n12 a_n2094_n4888# 0.585096f
C220 source.t22 a_n2094_n4888# 0.542781f
C221 source.t11 a_n2094_n4888# 0.542781f
C222 source.n13 a_n2094_n4888# 4.8527f
C223 source.n14 a_n2094_n4888# 0.453779f
C224 source.t3 a_n2094_n4888# 0.542781f
C225 source.t14 a_n2094_n4888# 0.542781f
C226 source.n15 a_n2094_n4888# 4.8527f
C227 source.n16 a_n2094_n4888# 0.453779f
C228 source.t21 a_n2094_n4888# 0.542781f
C229 source.t17 a_n2094_n4888# 0.542781f
C230 source.n17 a_n2094_n4888# 4.8527f
C231 source.n18 a_n2094_n4888# 0.453779f
C232 source.t23 a_n2094_n4888# 0.542781f
C233 source.t19 a_n2094_n4888# 0.542781f
C234 source.n19 a_n2094_n4888# 4.8527f
C235 source.n20 a_n2094_n4888# 0.453779f
C236 source.t7 a_n2094_n4888# 0.542781f
C237 source.t4 a_n2094_n4888# 0.542781f
C238 source.n21 a_n2094_n4888# 4.8527f
C239 source.n22 a_n2094_n4888# 0.453779f
C240 source.t16 a_n2094_n4888# 6.20312f
C241 source.n23 a_n2094_n4888# 3.22791f
C242 source.t35 a_n2094_n4888# 6.20309f
C243 source.n24 a_n2094_n4888# 3.22795f
C244 source.t43 a_n2094_n4888# 0.542781f
C245 source.t40 a_n2094_n4888# 0.542781f
C246 source.n25 a_n2094_n4888# 4.8527f
C247 source.n26 a_n2094_n4888# 0.45377f
C248 source.t38 a_n2094_n4888# 0.542781f
C249 source.t24 a_n2094_n4888# 0.542781f
C250 source.n27 a_n2094_n4888# 4.8527f
C251 source.n28 a_n2094_n4888# 0.45377f
C252 source.t33 a_n2094_n4888# 0.542781f
C253 source.t39 a_n2094_n4888# 0.542781f
C254 source.n29 a_n2094_n4888# 4.8527f
C255 source.n30 a_n2094_n4888# 0.45377f
C256 source.t41 a_n2094_n4888# 0.542781f
C257 source.t26 a_n2094_n4888# 0.542781f
C258 source.n31 a_n2094_n4888# 4.8527f
C259 source.n32 a_n2094_n4888# 0.45377f
C260 source.t28 a_n2094_n4888# 0.542781f
C261 source.t30 a_n2094_n4888# 0.542781f
C262 source.n33 a_n2094_n4888# 4.8527f
C263 source.n34 a_n2094_n4888# 0.45377f
C264 source.t32 a_n2094_n4888# 6.20309f
C265 source.n35 a_n2094_n4888# 0.58513f
C266 source.t8 a_n2094_n4888# 6.20309f
C267 source.n36 a_n2094_n4888# 0.58513f
C268 source.t5 a_n2094_n4888# 0.542781f
C269 source.t20 a_n2094_n4888# 0.542781f
C270 source.n37 a_n2094_n4888# 4.8527f
C271 source.n38 a_n2094_n4888# 0.45377f
C272 source.t10 a_n2094_n4888# 0.542781f
C273 source.t9 a_n2094_n4888# 0.542781f
C274 source.n39 a_n2094_n4888# 4.8527f
C275 source.n40 a_n2094_n4888# 0.45377f
C276 source.t6 a_n2094_n4888# 0.542781f
C277 source.t12 a_n2094_n4888# 0.542781f
C278 source.n41 a_n2094_n4888# 4.8527f
C279 source.n42 a_n2094_n4888# 0.45377f
C280 source.t13 a_n2094_n4888# 0.542781f
C281 source.t18 a_n2094_n4888# 0.542781f
C282 source.n43 a_n2094_n4888# 4.8527f
C283 source.n44 a_n2094_n4888# 0.45377f
C284 source.t1 a_n2094_n4888# 0.542781f
C285 source.t15 a_n2094_n4888# 0.542781f
C286 source.n45 a_n2094_n4888# 4.8527f
C287 source.n46 a_n2094_n4888# 0.45377f
C288 source.t0 a_n2094_n4888# 6.20309f
C289 source.n47 a_n2094_n4888# 0.77135f
C290 source.n48 a_n2094_n4888# 3.0856f
C291 plus.n0 a_n2094_n4888# 0.05238f
C292 plus.t2 a_n2094_n4888# 0.590107f
C293 plus.t6 a_n2094_n4888# 0.590107f
C294 plus.t11 a_n2094_n4888# 0.590107f
C295 plus.n1 a_n2094_n4888# 0.224593f
C296 plus.n2 a_n2094_n4888# 0.05238f
C297 plus.t21 a_n2094_n4888# 0.590107f
C298 plus.t4 a_n2094_n4888# 0.590107f
C299 plus.t7 a_n2094_n4888# 0.590107f
C300 plus.n3 a_n2094_n4888# 0.224593f
C301 plus.n4 a_n2094_n4888# 0.05238f
C302 plus.t12 a_n2094_n4888# 0.590107f
C303 plus.t13 a_n2094_n4888# 0.590107f
C304 plus.t22 a_n2094_n4888# 0.590107f
C305 plus.n5 a_n2094_n4888# 0.224593f
C306 plus.t8 a_n2094_n4888# 0.595374f
C307 plus.n6 a_n2094_n4888# 0.241466f
C308 plus.t5 a_n2094_n4888# 0.590107f
C309 plus.n7 a_n2094_n4888# 0.224593f
C310 plus.n8 a_n2094_n4888# 0.018345f
C311 plus.n9 a_n2094_n4888# 0.121794f
C312 plus.n10 a_n2094_n4888# 0.05238f
C313 plus.n11 a_n2094_n4888# 0.018345f
C314 plus.n12 a_n2094_n4888# 0.224593f
C315 plus.n13 a_n2094_n4888# 0.018345f
C316 plus.n14 a_n2094_n4888# 0.224593f
C317 plus.n15 a_n2094_n4888# 0.018345f
C318 plus.n16 a_n2094_n4888# 0.05238f
C319 plus.n17 a_n2094_n4888# 0.05238f
C320 plus.n18 a_n2094_n4888# 0.018345f
C321 plus.n19 a_n2094_n4888# 0.224593f
C322 plus.n20 a_n2094_n4888# 0.018345f
C323 plus.n21 a_n2094_n4888# 0.224593f
C324 plus.n22 a_n2094_n4888# 0.018345f
C325 plus.n23 a_n2094_n4888# 0.05238f
C326 plus.n24 a_n2094_n4888# 0.05238f
C327 plus.n25 a_n2094_n4888# 0.018345f
C328 plus.n26 a_n2094_n4888# 0.224593f
C329 plus.n27 a_n2094_n4888# 0.018345f
C330 plus.n28 a_n2094_n4888# 0.224593f
C331 plus.t18 a_n2094_n4888# 0.595374f
C332 plus.n29 a_n2094_n4888# 0.241384f
C333 plus.n30 a_n2094_n4888# 0.794043f
C334 plus.n31 a_n2094_n4888# 0.05238f
C335 plus.t19 a_n2094_n4888# 0.595374f
C336 plus.t14 a_n2094_n4888# 0.590107f
C337 plus.t9 a_n2094_n4888# 0.590107f
C338 plus.t10 a_n2094_n4888# 0.590107f
C339 plus.n32 a_n2094_n4888# 0.224593f
C340 plus.n33 a_n2094_n4888# 0.05238f
C341 plus.t15 a_n2094_n4888# 0.590107f
C342 plus.t20 a_n2094_n4888# 0.590107f
C343 plus.t17 a_n2094_n4888# 0.590107f
C344 plus.n34 a_n2094_n4888# 0.224593f
C345 plus.n35 a_n2094_n4888# 0.05238f
C346 plus.t23 a_n2094_n4888# 0.590107f
C347 plus.t16 a_n2094_n4888# 0.590107f
C348 plus.t1 a_n2094_n4888# 0.590107f
C349 plus.n36 a_n2094_n4888# 0.224593f
C350 plus.t0 a_n2094_n4888# 0.595374f
C351 plus.n37 a_n2094_n4888# 0.241466f
C352 plus.t3 a_n2094_n4888# 0.590107f
C353 plus.n38 a_n2094_n4888# 0.224593f
C354 plus.n39 a_n2094_n4888# 0.018345f
C355 plus.n40 a_n2094_n4888# 0.121794f
C356 plus.n41 a_n2094_n4888# 0.05238f
C357 plus.n42 a_n2094_n4888# 0.018345f
C358 plus.n43 a_n2094_n4888# 0.224593f
C359 plus.n44 a_n2094_n4888# 0.018345f
C360 plus.n45 a_n2094_n4888# 0.224593f
C361 plus.n46 a_n2094_n4888# 0.018345f
C362 plus.n47 a_n2094_n4888# 0.05238f
C363 plus.n48 a_n2094_n4888# 0.05238f
C364 plus.n49 a_n2094_n4888# 0.018345f
C365 plus.n50 a_n2094_n4888# 0.224593f
C366 plus.n51 a_n2094_n4888# 0.018345f
C367 plus.n52 a_n2094_n4888# 0.224593f
C368 plus.n53 a_n2094_n4888# 0.018345f
C369 plus.n54 a_n2094_n4888# 0.05238f
C370 plus.n55 a_n2094_n4888# 0.05238f
C371 plus.n56 a_n2094_n4888# 0.018345f
C372 plus.n57 a_n2094_n4888# 0.224593f
C373 plus.n58 a_n2094_n4888# 0.018345f
C374 plus.n59 a_n2094_n4888# 0.224593f
C375 plus.n60 a_n2094_n4888# 0.241384f
C376 plus.n61 a_n2094_n4888# 1.9122f
.ends

