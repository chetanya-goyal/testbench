* NGSPICE file created from diffpair573.ext - technology: sky130A

.subckt diffpair573 minus drain_right drain_left source plus
X0 drain_left.t7 plus.t0 source.t13 a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X1 drain_left.t6 plus.t1 source.t14 a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X2 drain_right.t7 minus.t0 source.t4 a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X3 source.t10 plus.t2 drain_left.t5 a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X4 a_n1246_n4888# a_n1246_n4888# a_n1246_n4888# a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.2
X5 drain_left.t4 plus.t3 source.t11 a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X6 a_n1246_n4888# a_n1246_n4888# a_n1246_n4888# a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X7 source.t0 minus.t1 drain_right.t6 a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X8 source.t15 minus.t2 drain_right.t5 a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X9 source.t2 minus.t3 drain_right.t4 a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X10 drain_right.t3 minus.t4 source.t1 a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X11 drain_right.t2 minus.t5 source.t5 a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
X12 source.t8 plus.t4 drain_left.t3 a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X13 a_n1246_n4888# a_n1246_n4888# a_n1246_n4888# a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X14 drain_right.t1 minus.t6 source.t6 a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X15 drain_left.t2 plus.t5 source.t9 a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.2
X16 source.t3 minus.t7 drain_right.t0 a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X17 source.t7 plus.t6 drain_left.t1 a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.2
X18 a_n1246_n4888# a_n1246_n4888# a_n1246_n4888# a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.2
X19 source.t12 plus.t7 drain_left.t0 a_n1246_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.2
R0 plus.n1 plus.t4 2609.74
R1 plus.n5 plus.t5 2609.74
R2 plus.n8 plus.t0 2609.74
R3 plus.n12 plus.t6 2609.74
R4 plus.n2 plus.t3 2566.65
R5 plus.n4 plus.t7 2566.65
R6 plus.n9 plus.t2 2566.65
R7 plus.n11 plus.t1 2566.65
R8 plus.n1 plus.n0 161.489
R9 plus.n8 plus.n7 161.489
R10 plus.n3 plus.n0 161.3
R11 plus.n6 plus.n5 161.3
R12 plus.n10 plus.n7 161.3
R13 plus.n13 plus.n12 161.3
R14 plus.n3 plus.n2 38.7066
R15 plus.n4 plus.n3 38.7066
R16 plus.n11 plus.n10 38.7066
R17 plus.n10 plus.n9 38.7066
R18 plus.n2 plus.n1 34.3247
R19 plus.n5 plus.n4 34.3247
R20 plus.n12 plus.n11 34.3247
R21 plus.n9 plus.n8 34.3247
R22 plus plus.n13 30.696
R23 plus plus.n6 15.1179
R24 plus.n6 plus.n0 0.189894
R25 plus.n13 plus.n7 0.189894
R26 source.n0 source.t9 44.1297
R27 source.n3 source.t8 44.1296
R28 source.n4 source.t6 44.1296
R29 source.n7 source.t3 44.1296
R30 source.n15 source.t1 44.1295
R31 source.n12 source.t15 44.1295
R32 source.n11 source.t13 44.1295
R33 source.n8 source.t7 44.1295
R34 source.n2 source.n1 43.1397
R35 source.n6 source.n5 43.1397
R36 source.n14 source.n13 43.1396
R37 source.n10 source.n9 43.1396
R38 source.n8 source.n7 27.8052
R39 source.n16 source.n0 22.3138
R40 source.n16 source.n15 5.49188
R41 source.n13 source.t5 0.9905
R42 source.n13 source.t0 0.9905
R43 source.n9 source.t14 0.9905
R44 source.n9 source.t10 0.9905
R45 source.n1 source.t11 0.9905
R46 source.n1 source.t12 0.9905
R47 source.n5 source.t4 0.9905
R48 source.n5 source.t2 0.9905
R49 source.n4 source.n3 0.470328
R50 source.n12 source.n11 0.470328
R51 source.n7 source.n6 0.457397
R52 source.n6 source.n4 0.457397
R53 source.n3 source.n2 0.457397
R54 source.n2 source.n0 0.457397
R55 source.n10 source.n8 0.457397
R56 source.n11 source.n10 0.457397
R57 source.n14 source.n12 0.457397
R58 source.n15 source.n14 0.457397
R59 source source.n16 0.188
R60 drain_left.n5 drain_left.n3 60.2753
R61 drain_left.n2 drain_left.n1 59.9915
R62 drain_left.n2 drain_left.n0 59.9915
R63 drain_left.n5 drain_left.n4 59.8185
R64 drain_left drain_left.n2 35.0268
R65 drain_left drain_left.n5 6.11011
R66 drain_left.n1 drain_left.t5 0.9905
R67 drain_left.n1 drain_left.t7 0.9905
R68 drain_left.n0 drain_left.t1 0.9905
R69 drain_left.n0 drain_left.t6 0.9905
R70 drain_left.n4 drain_left.t0 0.9905
R71 drain_left.n4 drain_left.t2 0.9905
R72 drain_left.n3 drain_left.t3 0.9905
R73 drain_left.n3 drain_left.t4 0.9905
R74 minus.n5 minus.t7 2609.74
R75 minus.n1 minus.t6 2609.74
R76 minus.n12 minus.t4 2609.74
R77 minus.n8 minus.t2 2609.74
R78 minus.n4 minus.t0 2566.65
R79 minus.n2 minus.t3 2566.65
R80 minus.n11 minus.t1 2566.65
R81 minus.n9 minus.t5 2566.65
R82 minus.n1 minus.n0 161.489
R83 minus.n8 minus.n7 161.489
R84 minus.n6 minus.n5 161.3
R85 minus.n3 minus.n0 161.3
R86 minus.n13 minus.n12 161.3
R87 minus.n10 minus.n7 161.3
R88 minus.n14 minus.n6 39.8452
R89 minus.n4 minus.n3 38.7066
R90 minus.n3 minus.n2 38.7066
R91 minus.n10 minus.n9 38.7066
R92 minus.n11 minus.n10 38.7066
R93 minus.n5 minus.n4 34.3247
R94 minus.n2 minus.n1 34.3247
R95 minus.n9 minus.n8 34.3247
R96 minus.n12 minus.n11 34.3247
R97 minus.n14 minus.n13 6.44368
R98 minus.n6 minus.n0 0.189894
R99 minus.n13 minus.n7 0.189894
R100 minus minus.n14 0.188
R101 drain_right.n5 drain_right.n3 60.2753
R102 drain_right.n2 drain_right.n1 59.9915
R103 drain_right.n2 drain_right.n0 59.9915
R104 drain_right.n5 drain_right.n4 59.8185
R105 drain_right drain_right.n2 34.4736
R106 drain_right drain_right.n5 6.11011
R107 drain_right.n1 drain_right.t6 0.9905
R108 drain_right.n1 drain_right.t3 0.9905
R109 drain_right.n0 drain_right.t5 0.9905
R110 drain_right.n0 drain_right.t2 0.9905
R111 drain_right.n3 drain_right.t4 0.9905
R112 drain_right.n3 drain_right.t1 0.9905
R113 drain_right.n4 drain_right.t0 0.9905
R114 drain_right.n4 drain_right.t7 0.9905
C0 drain_right source 31.5835f
C1 drain_right plus 0.269775f
C2 drain_right minus 4.14863f
C3 source drain_left 31.5849f
C4 drain_left plus 4.26543f
C5 drain_left minus 0.17017f
C6 source plus 3.30369f
C7 source minus 3.28965f
C8 minus plus 6.18982f
C9 drain_right drain_left 0.58123f
C10 drain_right a_n1246_n4888# 7.87608f
C11 drain_left a_n1246_n4888# 8.082531f
C12 source a_n1246_n4888# 12.714375f
C13 minus a_n1246_n4888# 5.332683f
C14 plus a_n1246_n4888# 8.09458f
C15 drain_right.t5 a_n1246_n4888# 0.600785f
C16 drain_right.t2 a_n1246_n4888# 0.600785f
C17 drain_right.n0 a_n1246_n4888# 5.49371f
C18 drain_right.t6 a_n1246_n4888# 0.600785f
C19 drain_right.t3 a_n1246_n4888# 0.600785f
C20 drain_right.n1 a_n1246_n4888# 5.49371f
C21 drain_right.n2 a_n1246_n4888# 3.11636f
C22 drain_right.t4 a_n1246_n4888# 0.600785f
C23 drain_right.t1 a_n1246_n4888# 0.600785f
C24 drain_right.n3 a_n1246_n4888# 5.49589f
C25 drain_right.t0 a_n1246_n4888# 0.600785f
C26 drain_right.t7 a_n1246_n4888# 0.600785f
C27 drain_right.n4 a_n1246_n4888# 5.4925f
C28 drain_right.n5 a_n1246_n4888# 1.18844f
C29 minus.n0 a_n1246_n4888# 0.129856f
C30 minus.t7 a_n1246_n4888# 0.676091f
C31 minus.t0 a_n1246_n4888# 0.671872f
C32 minus.t3 a_n1246_n4888# 0.671872f
C33 minus.t6 a_n1246_n4888# 0.676091f
C34 minus.n1 a_n1246_n4888# 0.272279f
C35 minus.n2 a_n1246_n4888# 0.255712f
C36 minus.n3 a_n1246_n4888# 0.020887f
C37 minus.n4 a_n1246_n4888# 0.255712f
C38 minus.n5 a_n1246_n4888# 0.272196f
C39 minus.n6 a_n1246_n4888# 2.43977f
C40 minus.n7 a_n1246_n4888# 0.129856f
C41 minus.t1 a_n1246_n4888# 0.671872f
C42 minus.t5 a_n1246_n4888# 0.671872f
C43 minus.t2 a_n1246_n4888# 0.676091f
C44 minus.n8 a_n1246_n4888# 0.272279f
C45 minus.n9 a_n1246_n4888# 0.255712f
C46 minus.n10 a_n1246_n4888# 0.020887f
C47 minus.n11 a_n1246_n4888# 0.255712f
C48 minus.t4 a_n1246_n4888# 0.676091f
C49 minus.n12 a_n1246_n4888# 0.272196f
C50 minus.n13 a_n1246_n4888# 0.381961f
C51 minus.n14 a_n1246_n4888# 2.93397f
C52 drain_left.t1 a_n1246_n4888# 0.601644f
C53 drain_left.t6 a_n1246_n4888# 0.601644f
C54 drain_left.n0 a_n1246_n4888# 5.50157f
C55 drain_left.t5 a_n1246_n4888# 0.601644f
C56 drain_left.t7 a_n1246_n4888# 0.601644f
C57 drain_left.n1 a_n1246_n4888# 5.50157f
C58 drain_left.n2 a_n1246_n4888# 3.20081f
C59 drain_left.t3 a_n1246_n4888# 0.601644f
C60 drain_left.t4 a_n1246_n4888# 0.601644f
C61 drain_left.n3 a_n1246_n4888# 5.50376f
C62 drain_left.t0 a_n1246_n4888# 0.601644f
C63 drain_left.t2 a_n1246_n4888# 0.601644f
C64 drain_left.n4 a_n1246_n4888# 5.50036f
C65 drain_left.n5 a_n1246_n4888# 1.19014f
C66 source.t9 a_n1246_n4888# 4.78283f
C67 source.n0 a_n1246_n4888# 2.0227f
C68 source.t11 a_n1246_n4888# 0.418504f
C69 source.t12 a_n1246_n4888# 0.418504f
C70 source.n1 a_n1246_n4888# 3.74161f
C71 source.n2 a_n1246_n4888# 0.349881f
C72 source.t8 a_n1246_n4888# 4.78284f
C73 source.n3 a_n1246_n4888# 0.451131f
C74 source.t6 a_n1246_n4888# 4.78284f
C75 source.n4 a_n1246_n4888# 0.451131f
C76 source.t4 a_n1246_n4888# 0.418504f
C77 source.t2 a_n1246_n4888# 0.418504f
C78 source.n5 a_n1246_n4888# 3.74161f
C79 source.n6 a_n1246_n4888# 0.349881f
C80 source.t3 a_n1246_n4888# 4.78284f
C81 source.n7 a_n1246_n4888# 2.48884f
C82 source.t7 a_n1246_n4888# 4.78281f
C83 source.n8 a_n1246_n4888# 2.48887f
C84 source.t14 a_n1246_n4888# 0.418504f
C85 source.t10 a_n1246_n4888# 0.418504f
C86 source.n9 a_n1246_n4888# 3.74162f
C87 source.n10 a_n1246_n4888# 0.349873f
C88 source.t13 a_n1246_n4888# 4.78281f
C89 source.n11 a_n1246_n4888# 0.451157f
C90 source.t15 a_n1246_n4888# 4.78281f
C91 source.n12 a_n1246_n4888# 0.451157f
C92 source.t5 a_n1246_n4888# 0.418504f
C93 source.t0 a_n1246_n4888# 0.418504f
C94 source.n13 a_n1246_n4888# 3.74162f
C95 source.n14 a_n1246_n4888# 0.349873f
C96 source.t1 a_n1246_n4888# 4.78281f
C97 source.n15 a_n1246_n4888# 0.59474f
C98 source.n16 a_n1246_n4888# 2.37911f
C99 plus.n0 a_n1246_n4888# 0.132944f
C100 plus.t7 a_n1246_n4888# 0.687852f
C101 plus.t3 a_n1246_n4888# 0.687852f
C102 plus.t4 a_n1246_n4888# 0.692171f
C103 plus.n1 a_n1246_n4888# 0.278755f
C104 plus.n2 a_n1246_n4888# 0.261794f
C105 plus.n3 a_n1246_n4888# 0.021384f
C106 plus.n4 a_n1246_n4888# 0.261794f
C107 plus.t5 a_n1246_n4888# 0.692171f
C108 plus.n5 a_n1246_n4888# 0.278671f
C109 plus.n6 a_n1246_n4888# 0.919176f
C110 plus.n7 a_n1246_n4888# 0.132944f
C111 plus.t6 a_n1246_n4888# 0.692171f
C112 plus.t1 a_n1246_n4888# 0.687852f
C113 plus.t2 a_n1246_n4888# 0.687852f
C114 plus.t0 a_n1246_n4888# 0.692171f
C115 plus.n8 a_n1246_n4888# 0.278755f
C116 plus.n9 a_n1246_n4888# 0.261794f
C117 plus.n10 a_n1246_n4888# 0.021384f
C118 plus.n11 a_n1246_n4888# 0.261794f
C119 plus.n12 a_n1246_n4888# 0.278671f
C120 plus.n13 a_n1246_n4888# 1.95754f
.ends

