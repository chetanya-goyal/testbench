* NGSPICE file created from diffpair346.ext - technology: sky130A

.subckt diffpair346 minus drain_right drain_left source plus
X0 source.t27 plus.t0 drain_left.t1 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X1 source.t26 plus.t1 drain_left.t4 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X2 source.t0 minus.t0 drain_right.t13 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X3 drain_left.t13 plus.t2 source.t25 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X4 source.t11 minus.t1 drain_right.t12 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X5 drain_right.t11 minus.t2 source.t1 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X6 source.t5 minus.t3 drain_right.t10 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X7 drain_left.t5 plus.t3 source.t24 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X8 drain_left.t10 plus.t4 source.t23 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X9 source.t8 minus.t4 drain_right.t9 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X10 drain_left.t11 plus.t5 source.t22 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X11 drain_left.t8 plus.t6 source.t21 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X12 drain_left.t7 plus.t7 source.t20 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X13 a_n1644_n2688# a_n1644_n2688# a_n1644_n2688# a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.25
X14 source.t2 minus.t5 drain_right.t8 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X15 drain_left.t12 plus.t8 source.t19 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X16 source.t18 plus.t9 drain_left.t2 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X17 drain_right.t7 minus.t6 source.t10 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X18 drain_right.t6 minus.t7 source.t4 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X19 drain_right.t5 minus.t8 source.t6 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X20 drain_right.t4 minus.t9 source.t9 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X21 a_n1644_n2688# a_n1644_n2688# a_n1644_n2688# a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
X22 source.t17 plus.t10 drain_left.t0 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X23 drain_left.t9 plus.t11 source.t16 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.25
X24 source.t3 minus.t10 drain_right.t3 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X25 drain_right.t2 minus.t11 source.t12 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X26 source.t15 plus.t12 drain_left.t3 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X27 drain_right.t1 minus.t12 source.t13 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X28 drain_right.t0 minus.t13 source.t7 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.25
X29 a_n1644_n2688# a_n1644_n2688# a_n1644_n2688# a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
X30 source.t14 plus.t13 drain_left.t6 a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.25
X31 a_n1644_n2688# a_n1644_n2688# a_n1644_n2688# a_n1644_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.25
R0 plus.n3 plus.t4 1027.97
R1 plus.n15 plus.t5 1027.97
R2 plus.n20 plus.t11 1027.97
R3 plus.n32 plus.t8 1027.97
R4 plus.n1 plus.t0 992.92
R5 plus.n4 plus.t1 992.92
R6 plus.n6 plus.t7 992.92
R7 plus.n12 plus.t6 992.92
R8 plus.n14 plus.t13 992.92
R9 plus.n18 plus.t12 992.92
R10 plus.n21 plus.t9 992.92
R11 plus.n23 plus.t3 992.92
R12 plus.n29 plus.t2 992.92
R13 plus.n31 plus.t10 992.92
R14 plus.n3 plus.n2 161.489
R15 plus.n20 plus.n19 161.489
R16 plus.n5 plus.n2 161.3
R17 plus.n8 plus.n7 161.3
R18 plus.n9 plus.n1 161.3
R19 plus.n11 plus.n10 161.3
R20 plus.n13 plus.n0 161.3
R21 plus.n16 plus.n15 161.3
R22 plus.n22 plus.n19 161.3
R23 plus.n25 plus.n24 161.3
R24 plus.n26 plus.n18 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n17 161.3
R27 plus.n33 plus.n32 161.3
R28 plus.n7 plus.n1 73.0308
R29 plus.n11 plus.n1 73.0308
R30 plus.n28 plus.n18 73.0308
R31 plus.n24 plus.n18 73.0308
R32 plus.n6 plus.n5 61.346
R33 plus.n13 plus.n12 61.346
R34 plus.n30 plus.n29 61.346
R35 plus.n23 plus.n22 61.346
R36 plus.n4 plus.n3 49.6611
R37 plus.n15 plus.n14 49.6611
R38 plus.n32 plus.n31 49.6611
R39 plus.n21 plus.n20 49.6611
R40 plus plus.n33 28.0445
R41 plus.n5 plus.n4 23.3702
R42 plus.n14 plus.n13 23.3702
R43 plus.n31 plus.n30 23.3702
R44 plus.n22 plus.n21 23.3702
R45 plus.n7 plus.n6 11.6853
R46 plus.n12 plus.n11 11.6853
R47 plus.n29 plus.n28 11.6853
R48 plus.n24 plus.n23 11.6853
R49 plus plus.n16 10.9588
R50 plus.n8 plus.n2 0.189894
R51 plus.n9 plus.n8 0.189894
R52 plus.n10 plus.n9 0.189894
R53 plus.n10 plus.n0 0.189894
R54 plus.n16 plus.n0 0.189894
R55 plus.n33 plus.n17 0.189894
R56 plus.n27 plus.n17 0.189894
R57 plus.n27 plus.n26 0.189894
R58 plus.n26 plus.n25 0.189894
R59 plus.n25 plus.n19 0.189894
R60 drain_left.n7 drain_left.t10 68.2376
R61 drain_left.n1 drain_left.t12 68.2373
R62 drain_left.n4 drain_left.n2 66.0373
R63 drain_left.n9 drain_left.n8 65.5376
R64 drain_left.n7 drain_left.n6 65.5376
R65 drain_left.n11 drain_left.n10 65.5374
R66 drain_left.n4 drain_left.n3 65.5373
R67 drain_left.n1 drain_left.n0 65.5373
R68 drain_left drain_left.n5 27.9693
R69 drain_left drain_left.n11 6.15322
R70 drain_left.n2 drain_left.t2 2.2005
R71 drain_left.n2 drain_left.t9 2.2005
R72 drain_left.n3 drain_left.t3 2.2005
R73 drain_left.n3 drain_left.t5 2.2005
R74 drain_left.n0 drain_left.t0 2.2005
R75 drain_left.n0 drain_left.t13 2.2005
R76 drain_left.n10 drain_left.t6 2.2005
R77 drain_left.n10 drain_left.t11 2.2005
R78 drain_left.n8 drain_left.t1 2.2005
R79 drain_left.n8 drain_left.t8 2.2005
R80 drain_left.n6 drain_left.t4 2.2005
R81 drain_left.n6 drain_left.t7 2.2005
R82 drain_left.n9 drain_left.n7 0.5005
R83 drain_left.n11 drain_left.n9 0.5005
R84 drain_left.n5 drain_left.n1 0.320154
R85 drain_left.n5 drain_left.n4 0.070154
R86 source.n7 source.t9 51.0588
R87 source.n27 source.t4 51.0586
R88 source.n20 source.t16 51.0586
R89 source.n0 source.t22 51.0586
R90 source.n2 source.n1 48.8588
R91 source.n4 source.n3 48.8588
R92 source.n6 source.n5 48.8588
R93 source.n9 source.n8 48.8588
R94 source.n11 source.n10 48.8588
R95 source.n13 source.n12 48.8588
R96 source.n26 source.n25 48.8586
R97 source.n24 source.n23 48.8586
R98 source.n22 source.n21 48.8586
R99 source.n19 source.n18 48.8586
R100 source.n17 source.n16 48.8586
R101 source.n15 source.n14 48.8586
R102 source.n15 source.n13 20.015
R103 source.n28 source.n0 14.0021
R104 source.n28 source.n27 5.51343
R105 source.n25 source.t1 2.2005
R106 source.n25 source.t3 2.2005
R107 source.n23 source.t6 2.2005
R108 source.n23 source.t2 2.2005
R109 source.n21 source.t12 2.2005
R110 source.n21 source.t0 2.2005
R111 source.n18 source.t24 2.2005
R112 source.n18 source.t18 2.2005
R113 source.n16 source.t25 2.2005
R114 source.n16 source.t15 2.2005
R115 source.n14 source.t19 2.2005
R116 source.n14 source.t17 2.2005
R117 source.n1 source.t21 2.2005
R118 source.n1 source.t14 2.2005
R119 source.n3 source.t20 2.2005
R120 source.n3 source.t27 2.2005
R121 source.n5 source.t23 2.2005
R122 source.n5 source.t26 2.2005
R123 source.n8 source.t10 2.2005
R124 source.n8 source.t5 2.2005
R125 source.n10 source.t13 2.2005
R126 source.n10 source.t11 2.2005
R127 source.n12 source.t7 2.2005
R128 source.n12 source.t8 2.2005
R129 source.n7 source.n6 0.720328
R130 source.n22 source.n20 0.720328
R131 source.n13 source.n11 0.5005
R132 source.n11 source.n9 0.5005
R133 source.n9 source.n7 0.5005
R134 source.n6 source.n4 0.5005
R135 source.n4 source.n2 0.5005
R136 source.n2 source.n0 0.5005
R137 source.n17 source.n15 0.5005
R138 source.n19 source.n17 0.5005
R139 source.n20 source.n19 0.5005
R140 source.n24 source.n22 0.5005
R141 source.n26 source.n24 0.5005
R142 source.n27 source.n26 0.5005
R143 source source.n28 0.188
R144 minus.n15 minus.t13 1027.97
R145 minus.n3 minus.t9 1027.97
R146 minus.n32 minus.t7 1027.97
R147 minus.n20 minus.t11 1027.97
R148 minus.n1 minus.t1 992.92
R149 minus.n14 minus.t4 992.92
R150 minus.n12 minus.t12 992.92
R151 minus.n6 minus.t6 992.92
R152 minus.n4 minus.t3 992.92
R153 minus.n18 minus.t5 992.92
R154 minus.n31 minus.t10 992.92
R155 minus.n29 minus.t2 992.92
R156 minus.n23 minus.t8 992.92
R157 minus.n21 minus.t0 992.92
R158 minus.n3 minus.n2 161.489
R159 minus.n20 minus.n19 161.489
R160 minus.n16 minus.n15 161.3
R161 minus.n13 minus.n0 161.3
R162 minus.n11 minus.n10 161.3
R163 minus.n9 minus.n1 161.3
R164 minus.n8 minus.n7 161.3
R165 minus.n5 minus.n2 161.3
R166 minus.n33 minus.n32 161.3
R167 minus.n30 minus.n17 161.3
R168 minus.n28 minus.n27 161.3
R169 minus.n26 minus.n18 161.3
R170 minus.n25 minus.n24 161.3
R171 minus.n22 minus.n19 161.3
R172 minus.n11 minus.n1 73.0308
R173 minus.n7 minus.n1 73.0308
R174 minus.n24 minus.n18 73.0308
R175 minus.n28 minus.n18 73.0308
R176 minus.n13 minus.n12 61.346
R177 minus.n6 minus.n5 61.346
R178 minus.n23 minus.n22 61.346
R179 minus.n30 minus.n29 61.346
R180 minus.n15 minus.n14 49.6611
R181 minus.n4 minus.n3 49.6611
R182 minus.n21 minus.n20 49.6611
R183 minus.n32 minus.n31 49.6611
R184 minus.n34 minus.n16 33.027
R185 minus.n14 minus.n13 23.3702
R186 minus.n5 minus.n4 23.3702
R187 minus.n22 minus.n21 23.3702
R188 minus.n31 minus.n30 23.3702
R189 minus.n12 minus.n11 11.6853
R190 minus.n7 minus.n6 11.6853
R191 minus.n24 minus.n23 11.6853
R192 minus.n29 minus.n28 11.6853
R193 minus.n34 minus.n33 6.45126
R194 minus.n16 minus.n0 0.189894
R195 minus.n10 minus.n0 0.189894
R196 minus.n10 minus.n9 0.189894
R197 minus.n9 minus.n8 0.189894
R198 minus.n8 minus.n2 0.189894
R199 minus.n25 minus.n19 0.189894
R200 minus.n26 minus.n25 0.189894
R201 minus.n27 minus.n26 0.189894
R202 minus.n27 minus.n17 0.189894
R203 minus.n33 minus.n17 0.189894
R204 minus minus.n34 0.188
R205 drain_right.n1 drain_right.t2 68.2373
R206 drain_right.n11 drain_right.t0 67.7376
R207 drain_right.n8 drain_right.n6 66.0374
R208 drain_right.n4 drain_right.n2 66.0373
R209 drain_right.n8 drain_right.n7 65.5376
R210 drain_right.n10 drain_right.n9 65.5376
R211 drain_right.n4 drain_right.n3 65.5373
R212 drain_right.n1 drain_right.n0 65.5373
R213 drain_right drain_right.n5 27.4161
R214 drain_right drain_right.n11 5.90322
R215 drain_right.n2 drain_right.t3 2.2005
R216 drain_right.n2 drain_right.t6 2.2005
R217 drain_right.n3 drain_right.t8 2.2005
R218 drain_right.n3 drain_right.t11 2.2005
R219 drain_right.n0 drain_right.t13 2.2005
R220 drain_right.n0 drain_right.t5 2.2005
R221 drain_right.n6 drain_right.t10 2.2005
R222 drain_right.n6 drain_right.t4 2.2005
R223 drain_right.n7 drain_right.t12 2.2005
R224 drain_right.n7 drain_right.t7 2.2005
R225 drain_right.n9 drain_right.t9 2.2005
R226 drain_right.n9 drain_right.t1 2.2005
R227 drain_right.n11 drain_right.n10 0.5005
R228 drain_right.n10 drain_right.n8 0.5005
R229 drain_right.n5 drain_right.n1 0.320154
R230 drain_right.n5 drain_right.n4 0.070154
C0 source drain_left 23.4622f
C1 drain_right minus 3.58976f
C2 drain_right plus 0.314441f
C3 plus minus 4.65065f
C4 drain_right drain_left 0.8398f
C5 drain_right source 23.4536f
C6 minus drain_left 0.171605f
C7 plus drain_left 3.74592f
C8 minus source 3.34075f
C9 plus source 3.35529f
C10 drain_right a_n1644_n2688# 6.48726f
C11 drain_left a_n1644_n2688# 6.75287f
C12 source a_n1644_n2688# 5.097322f
C13 minus a_n1644_n2688# 6.184156f
C14 plus a_n1644_n2688# 7.99485f
C15 drain_right.t2 a_n1644_n2688# 2.56836f
C16 drain_right.t13 a_n1644_n2688# 0.230417f
C17 drain_right.t5 a_n1644_n2688# 0.230417f
C18 drain_right.n0 a_n1644_n2688# 2.01538f
C19 drain_right.n1 a_n1644_n2688# 0.747615f
C20 drain_right.t3 a_n1644_n2688# 0.230417f
C21 drain_right.t6 a_n1644_n2688# 0.230417f
C22 drain_right.n2 a_n1644_n2688# 2.01823f
C23 drain_right.t8 a_n1644_n2688# 0.230417f
C24 drain_right.t11 a_n1644_n2688# 0.230417f
C25 drain_right.n3 a_n1644_n2688# 2.01538f
C26 drain_right.n4 a_n1644_n2688# 0.703864f
C27 drain_right.n5 a_n1644_n2688# 1.22383f
C28 drain_right.t10 a_n1644_n2688# 0.230417f
C29 drain_right.t4 a_n1644_n2688# 0.230417f
C30 drain_right.n6 a_n1644_n2688# 2.01823f
C31 drain_right.t12 a_n1644_n2688# 0.230417f
C32 drain_right.t7 a_n1644_n2688# 0.230417f
C33 drain_right.n7 a_n1644_n2688# 2.01538f
C34 drain_right.n8 a_n1644_n2688# 0.738007f
C35 drain_right.t9 a_n1644_n2688# 0.230417f
C36 drain_right.t1 a_n1644_n2688# 0.230417f
C37 drain_right.n9 a_n1644_n2688# 2.01538f
C38 drain_right.n10 a_n1644_n2688# 0.363901f
C39 drain_right.t0 a_n1644_n2688# 2.56541f
C40 drain_right.n11 a_n1644_n2688# 0.669943f
C41 minus.n0 a_n1644_n2688# 0.052789f
C42 minus.t13 a_n1644_n2688# 0.341436f
C43 minus.t4 a_n1644_n2688# 0.336562f
C44 minus.t12 a_n1644_n2688# 0.336562f
C45 minus.t1 a_n1644_n2688# 0.336562f
C46 minus.n1 a_n1644_n2688# 0.160766f
C47 minus.n2 a_n1644_n2688# 0.112993f
C48 minus.t6 a_n1644_n2688# 0.336562f
C49 minus.t3 a_n1644_n2688# 0.336562f
C50 minus.t9 a_n1644_n2688# 0.341436f
C51 minus.n3 a_n1644_n2688# 0.158241f
C52 minus.n4 a_n1644_n2688# 0.143255f
C53 minus.n5 a_n1644_n2688# 0.020116f
C54 minus.n6 a_n1644_n2688# 0.143255f
C55 minus.n7 a_n1644_n2688# 0.020116f
C56 minus.n8 a_n1644_n2688# 0.052789f
C57 minus.n9 a_n1644_n2688# 0.052789f
C58 minus.n10 a_n1644_n2688# 0.052789f
C59 minus.n11 a_n1644_n2688# 0.020116f
C60 minus.n12 a_n1644_n2688# 0.143255f
C61 minus.n13 a_n1644_n2688# 0.020116f
C62 minus.n14 a_n1644_n2688# 0.143255f
C63 minus.n15 a_n1644_n2688# 0.158171f
C64 minus.n16 a_n1644_n2688# 1.60984f
C65 minus.n17 a_n1644_n2688# 0.052789f
C66 minus.t10 a_n1644_n2688# 0.336562f
C67 minus.t2 a_n1644_n2688# 0.336562f
C68 minus.t5 a_n1644_n2688# 0.336562f
C69 minus.n18 a_n1644_n2688# 0.160766f
C70 minus.n19 a_n1644_n2688# 0.112993f
C71 minus.t8 a_n1644_n2688# 0.336562f
C72 minus.t0 a_n1644_n2688# 0.336562f
C73 minus.t11 a_n1644_n2688# 0.341436f
C74 minus.n20 a_n1644_n2688# 0.158241f
C75 minus.n21 a_n1644_n2688# 0.143255f
C76 minus.n22 a_n1644_n2688# 0.020116f
C77 minus.n23 a_n1644_n2688# 0.143255f
C78 minus.n24 a_n1644_n2688# 0.020116f
C79 minus.n25 a_n1644_n2688# 0.052789f
C80 minus.n26 a_n1644_n2688# 0.052789f
C81 minus.n27 a_n1644_n2688# 0.052789f
C82 minus.n28 a_n1644_n2688# 0.020116f
C83 minus.n29 a_n1644_n2688# 0.143255f
C84 minus.n30 a_n1644_n2688# 0.020116f
C85 minus.n31 a_n1644_n2688# 0.143255f
C86 minus.t7 a_n1644_n2688# 0.341436f
C87 minus.n32 a_n1644_n2688# 0.158171f
C88 minus.n33 a_n1644_n2688# 0.339044f
C89 minus.n34 a_n1644_n2688# 1.97547f
C90 source.t22 a_n1644_n2688# 2.57936f
C91 source.n0 a_n1644_n2688# 1.47529f
C92 source.t21 a_n1644_n2688# 0.241888f
C93 source.t14 a_n1644_n2688# 0.241888f
C94 source.n1 a_n1644_n2688# 2.02493f
C95 source.n2 a_n1644_n2688# 0.426578f
C96 source.t20 a_n1644_n2688# 0.241888f
C97 source.t27 a_n1644_n2688# 0.241888f
C98 source.n3 a_n1644_n2688# 2.02493f
C99 source.n4 a_n1644_n2688# 0.426578f
C100 source.t23 a_n1644_n2688# 0.241888f
C101 source.t26 a_n1644_n2688# 0.241888f
C102 source.n5 a_n1644_n2688# 2.02493f
C103 source.n6 a_n1644_n2688# 0.450669f
C104 source.t9 a_n1644_n2688# 2.57937f
C105 source.n7 a_n1644_n2688# 0.555922f
C106 source.t10 a_n1644_n2688# 0.241888f
C107 source.t5 a_n1644_n2688# 0.241888f
C108 source.n8 a_n1644_n2688# 2.02493f
C109 source.n9 a_n1644_n2688# 0.426578f
C110 source.t13 a_n1644_n2688# 0.241888f
C111 source.t11 a_n1644_n2688# 0.241888f
C112 source.n10 a_n1644_n2688# 2.02493f
C113 source.n11 a_n1644_n2688# 0.426578f
C114 source.t7 a_n1644_n2688# 0.241888f
C115 source.t8 a_n1644_n2688# 0.241888f
C116 source.n12 a_n1644_n2688# 2.02493f
C117 source.n13 a_n1644_n2688# 1.91747f
C118 source.t19 a_n1644_n2688# 0.241888f
C119 source.t17 a_n1644_n2688# 0.241888f
C120 source.n14 a_n1644_n2688# 2.02492f
C121 source.n15 a_n1644_n2688# 1.91748f
C122 source.t25 a_n1644_n2688# 0.241888f
C123 source.t15 a_n1644_n2688# 0.241888f
C124 source.n16 a_n1644_n2688# 2.02492f
C125 source.n17 a_n1644_n2688# 0.426584f
C126 source.t24 a_n1644_n2688# 0.241888f
C127 source.t18 a_n1644_n2688# 0.241888f
C128 source.n18 a_n1644_n2688# 2.02492f
C129 source.n19 a_n1644_n2688# 0.426584f
C130 source.t16 a_n1644_n2688# 2.57936f
C131 source.n20 a_n1644_n2688# 0.555928f
C132 source.t12 a_n1644_n2688# 0.241888f
C133 source.t0 a_n1644_n2688# 0.241888f
C134 source.n21 a_n1644_n2688# 2.02492f
C135 source.n22 a_n1644_n2688# 0.450675f
C136 source.t6 a_n1644_n2688# 0.241888f
C137 source.t2 a_n1644_n2688# 0.241888f
C138 source.n23 a_n1644_n2688# 2.02492f
C139 source.n24 a_n1644_n2688# 0.426584f
C140 source.t1 a_n1644_n2688# 0.241888f
C141 source.t3 a_n1644_n2688# 0.241888f
C142 source.n25 a_n1644_n2688# 2.02492f
C143 source.n26 a_n1644_n2688# 0.426584f
C144 source.t4 a_n1644_n2688# 2.57936f
C145 source.n27 a_n1644_n2688# 0.716741f
C146 source.n28 a_n1644_n2688# 1.76803f
C147 drain_left.t12 a_n1644_n2688# 2.56584f
C148 drain_left.t0 a_n1644_n2688# 0.230191f
C149 drain_left.t13 a_n1644_n2688# 0.230191f
C150 drain_left.n0 a_n1644_n2688# 2.0134f
C151 drain_left.n1 a_n1644_n2688# 0.746881f
C152 drain_left.t2 a_n1644_n2688# 0.230191f
C153 drain_left.t9 a_n1644_n2688# 0.230191f
C154 drain_left.n2 a_n1644_n2688# 2.01625f
C155 drain_left.t3 a_n1644_n2688# 0.230191f
C156 drain_left.t5 a_n1644_n2688# 0.230191f
C157 drain_left.n3 a_n1644_n2688# 2.0134f
C158 drain_left.n4 a_n1644_n2688# 0.703173f
C159 drain_left.n5 a_n1644_n2688# 1.28948f
C160 drain_left.t10 a_n1644_n2688# 2.56584f
C161 drain_left.t4 a_n1644_n2688# 0.230191f
C162 drain_left.t7 a_n1644_n2688# 0.230191f
C163 drain_left.n6 a_n1644_n2688# 2.0134f
C164 drain_left.n7 a_n1644_n2688# 0.763334f
C165 drain_left.t1 a_n1644_n2688# 0.230191f
C166 drain_left.t8 a_n1644_n2688# 0.230191f
C167 drain_left.n8 a_n1644_n2688# 2.0134f
C168 drain_left.n9 a_n1644_n2688# 0.363544f
C169 drain_left.t6 a_n1644_n2688# 0.230191f
C170 drain_left.t11 a_n1644_n2688# 0.230191f
C171 drain_left.n10 a_n1644_n2688# 2.0134f
C172 drain_left.n11 a_n1644_n2688# 0.630714f
C173 plus.n0 a_n1644_n2688# 0.054198f
C174 plus.t13 a_n1644_n2688# 0.345545f
C175 plus.t6 a_n1644_n2688# 0.345545f
C176 plus.t0 a_n1644_n2688# 0.345545f
C177 plus.n1 a_n1644_n2688# 0.165057f
C178 plus.n2 a_n1644_n2688# 0.116009f
C179 plus.t7 a_n1644_n2688# 0.345545f
C180 plus.t1 a_n1644_n2688# 0.345545f
C181 plus.t4 a_n1644_n2688# 0.350549f
C182 plus.n3 a_n1644_n2688# 0.162465f
C183 plus.n4 a_n1644_n2688# 0.147078f
C184 plus.n5 a_n1644_n2688# 0.020652f
C185 plus.n6 a_n1644_n2688# 0.147078f
C186 plus.n7 a_n1644_n2688# 0.020652f
C187 plus.n8 a_n1644_n2688# 0.054198f
C188 plus.n9 a_n1644_n2688# 0.054198f
C189 plus.n10 a_n1644_n2688# 0.054198f
C190 plus.n11 a_n1644_n2688# 0.020652f
C191 plus.n12 a_n1644_n2688# 0.147078f
C192 plus.n13 a_n1644_n2688# 0.020652f
C193 plus.n14 a_n1644_n2688# 0.147078f
C194 plus.t5 a_n1644_n2688# 0.350549f
C195 plus.n15 a_n1644_n2688# 0.162392f
C196 plus.n16 a_n1644_n2688# 0.525967f
C197 plus.n17 a_n1644_n2688# 0.054198f
C198 plus.t8 a_n1644_n2688# 0.350549f
C199 plus.t10 a_n1644_n2688# 0.345545f
C200 plus.t2 a_n1644_n2688# 0.345545f
C201 plus.t12 a_n1644_n2688# 0.345545f
C202 plus.n18 a_n1644_n2688# 0.165057f
C203 plus.n19 a_n1644_n2688# 0.116009f
C204 plus.t3 a_n1644_n2688# 0.345545f
C205 plus.t9 a_n1644_n2688# 0.345545f
C206 plus.t11 a_n1644_n2688# 0.350549f
C207 plus.n20 a_n1644_n2688# 0.162465f
C208 plus.n21 a_n1644_n2688# 0.147078f
C209 plus.n22 a_n1644_n2688# 0.020652f
C210 plus.n23 a_n1644_n2688# 0.147078f
C211 plus.n24 a_n1644_n2688# 0.020652f
C212 plus.n25 a_n1644_n2688# 0.054198f
C213 plus.n26 a_n1644_n2688# 0.054198f
C214 plus.n27 a_n1644_n2688# 0.054198f
C215 plus.n28 a_n1644_n2688# 0.020652f
C216 plus.n29 a_n1644_n2688# 0.147078f
C217 plus.n30 a_n1644_n2688# 0.020652f
C218 plus.n31 a_n1644_n2688# 0.147078f
C219 plus.n32 a_n1644_n2688# 0.162392f
C220 plus.n33 a_n1644_n2688# 1.43954f
.ends

