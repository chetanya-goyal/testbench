* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t27 minus.t0 drain_right.t2 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X1 drain_right.t11 minus.t1 source.t26 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X2 a_n2044_n1288# a_n2044_n1288# a_n2044_n1288# a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.5
X3 source.t25 minus.t2 drain_right.t3 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X4 source.t1 plus.t0 drain_left.t13 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X5 a_n2044_n1288# a_n2044_n1288# a_n2044_n1288# a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X6 a_n2044_n1288# a_n2044_n1288# a_n2044_n1288# a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X7 source.t3 plus.t1 drain_left.t12 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X8 source.t24 minus.t3 drain_right.t5 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X9 drain_left.t11 plus.t2 source.t8 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X10 source.t5 plus.t3 drain_left.t10 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X11 drain_right.t6 minus.t4 source.t23 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X12 drain_left.t9 plus.t4 source.t12 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X13 drain_right.t1 minus.t5 source.t22 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X14 drain_right.t10 minus.t6 source.t21 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X15 drain_right.t0 minus.t7 source.t20 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X16 source.t13 plus.t5 drain_left.t8 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X17 drain_left.t7 plus.t6 source.t4 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X18 a_n2044_n1288# a_n2044_n1288# a_n2044_n1288# a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X19 drain_left.t6 plus.t7 source.t7 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X20 source.t19 minus.t8 drain_right.t9 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X21 drain_right.t7 minus.t9 source.t18 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X22 source.t10 plus.t8 drain_left.t5 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X23 drain_right.t4 minus.t10 source.t17 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X24 source.t16 minus.t11 drain_right.t8 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X25 drain_left.t4 plus.t9 source.t6 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X26 drain_right.t12 minus.t12 source.t15 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X27 drain_left.t3 plus.t10 source.t9 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X28 source.t14 minus.t13 drain_right.t13 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X29 drain_left.t2 plus.t11 source.t0 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X30 drain_left.t1 plus.t12 source.t11 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X31 source.t2 plus.t13 drain_left.t0 a_n2044_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
R0 minus.n4 minus.t9 195.948
R1 minus.n20 minus.t12 195.948
R2 minus.n3 minus.t3 174.966
R3 minus.n7 minus.t6 174.966
R4 minus.n8 minus.t11 174.966
R5 minus.n1 minus.t5 174.966
R6 minus.n13 minus.t8 174.966
R7 minus.n14 minus.t1 174.966
R8 minus.n19 minus.t0 174.966
R9 minus.n23 minus.t10 174.966
R10 minus.n24 minus.t13 174.966
R11 minus.n17 minus.t7 174.966
R12 minus.n29 minus.t2 174.966
R13 minus.n30 minus.t4 174.966
R14 minus.n15 minus.n14 161.3
R15 minus.n13 minus.n0 161.3
R16 minus.n12 minus.n11 161.3
R17 minus.n10 minus.n1 161.3
R18 minus.n7 minus.n2 161.3
R19 minus.n6 minus.n5 161.3
R20 minus.n31 minus.n30 161.3
R21 minus.n29 minus.n16 161.3
R22 minus.n28 minus.n27 161.3
R23 minus.n26 minus.n17 161.3
R24 minus.n23 minus.n18 161.3
R25 minus.n22 minus.n21 161.3
R26 minus.n9 minus.n8 80.6037
R27 minus.n25 minus.n24 80.6037
R28 minus.n5 minus.n4 70.4033
R29 minus.n21 minus.n20 70.4033
R30 minus.n8 minus.n7 48.2005
R31 minus.n8 minus.n1 48.2005
R32 minus.n14 minus.n13 48.2005
R33 minus.n24 minus.n23 48.2005
R34 minus.n24 minus.n17 48.2005
R35 minus.n30 minus.n29 48.2005
R36 minus.n32 minus.n15 29.3812
R37 minus.n7 minus.n6 24.8308
R38 minus.n12 minus.n1 24.8308
R39 minus.n23 minus.n22 24.8308
R40 minus.n28 minus.n17 24.8308
R41 minus.n6 minus.n3 23.3702
R42 minus.n13 minus.n12 23.3702
R43 minus.n22 minus.n19 23.3702
R44 minus.n29 minus.n28 23.3702
R45 minus.n4 minus.n3 20.9576
R46 minus.n20 minus.n19 20.9576
R47 minus.n32 minus.n31 6.5933
R48 minus.n10 minus.n9 0.285035
R49 minus.n9 minus.n2 0.285035
R50 minus.n25 minus.n18 0.285035
R51 minus.n26 minus.n25 0.285035
R52 minus.n15 minus.n0 0.189894
R53 minus.n11 minus.n0 0.189894
R54 minus.n11 minus.n10 0.189894
R55 minus.n5 minus.n2 0.189894
R56 minus.n21 minus.n18 0.189894
R57 minus.n27 minus.n26 0.189894
R58 minus.n27 minus.n16 0.189894
R59 minus.n31 minus.n16 0.189894
R60 minus minus.n32 0.188
R61 drain_right.n2 drain_right.n0 289.615
R62 drain_right.n20 drain_right.n18 289.615
R63 drain_right.n3 drain_right.n2 185
R64 drain_right.n21 drain_right.n20 185
R65 drain_right.t12 drain_right.n1 167.117
R66 drain_right.t11 drain_right.n19 167.117
R67 drain_right.n15 drain_right.n13 101.511
R68 drain_right.n11 drain_right.n9 101.511
R69 drain_right.n15 drain_right.n14 100.796
R70 drain_right.n17 drain_right.n16 100.796
R71 drain_right.n11 drain_right.n10 100.796
R72 drain_right.n8 drain_right.n7 100.796
R73 drain_right.n2 drain_right.t12 52.3082
R74 drain_right.n20 drain_right.t11 52.3082
R75 drain_right.n8 drain_right.n6 48.8039
R76 drain_right.n25 drain_right.n24 48.0884
R77 drain_right drain_right.n12 23.3523
R78 drain_right.n9 drain_right.t3 9.9005
R79 drain_right.n9 drain_right.t6 9.9005
R80 drain_right.n10 drain_right.t13 9.9005
R81 drain_right.n10 drain_right.t0 9.9005
R82 drain_right.n7 drain_right.t2 9.9005
R83 drain_right.n7 drain_right.t4 9.9005
R84 drain_right.n13 drain_right.t5 9.9005
R85 drain_right.n13 drain_right.t7 9.9005
R86 drain_right.n14 drain_right.t8 9.9005
R87 drain_right.n14 drain_right.t10 9.9005
R88 drain_right.n16 drain_right.t9 9.9005
R89 drain_right.n16 drain_right.t1 9.9005
R90 drain_right.n3 drain_right.n1 9.71174
R91 drain_right.n21 drain_right.n19 9.71174
R92 drain_right.n6 drain_right.n5 9.45567
R93 drain_right.n24 drain_right.n23 9.45567
R94 drain_right.n5 drain_right.n4 9.3005
R95 drain_right.n23 drain_right.n22 9.3005
R96 drain_right.n6 drain_right.n0 8.14595
R97 drain_right.n24 drain_right.n18 8.14595
R98 drain_right.n4 drain_right.n3 7.3702
R99 drain_right.n22 drain_right.n21 7.3702
R100 drain_right drain_right.n25 6.01097
R101 drain_right.n4 drain_right.n0 5.81868
R102 drain_right.n22 drain_right.n18 5.81868
R103 drain_right.n5 drain_right.n1 3.44771
R104 drain_right.n23 drain_right.n19 3.44771
R105 drain_right.n25 drain_right.n17 0.716017
R106 drain_right.n17 drain_right.n15 0.716017
R107 drain_right.n12 drain_right.n8 0.481792
R108 drain_right.n12 drain_right.n11 0.124033
R109 source.n50 source.n48 289.615
R110 source.n36 source.n34 289.615
R111 source.n2 source.n0 289.615
R112 source.n16 source.n14 289.615
R113 source.n51 source.n50 185
R114 source.n37 source.n36 185
R115 source.n3 source.n2 185
R116 source.n17 source.n16 185
R117 source.t23 source.n49 167.117
R118 source.t11 source.n35 167.117
R119 source.t7 source.n1 167.117
R120 source.t18 source.n15 167.117
R121 source.n9 source.n8 84.1169
R122 source.n11 source.n10 84.1169
R123 source.n13 source.n12 84.1169
R124 source.n23 source.n22 84.1169
R125 source.n25 source.n24 84.1169
R126 source.n27 source.n26 84.1169
R127 source.n47 source.n46 84.1168
R128 source.n45 source.n44 84.1168
R129 source.n43 source.n42 84.1168
R130 source.n33 source.n32 84.1168
R131 source.n31 source.n30 84.1168
R132 source.n29 source.n28 84.1168
R133 source.n50 source.t23 52.3082
R134 source.n36 source.t11 52.3082
R135 source.n2 source.t7 52.3082
R136 source.n16 source.t18 52.3082
R137 source.n55 source.n54 31.4096
R138 source.n41 source.n40 31.4096
R139 source.n7 source.n6 31.4096
R140 source.n21 source.n20 31.4096
R141 source.n29 source.n27 15.143
R142 source.n46 source.t20 9.9005
R143 source.n46 source.t25 9.9005
R144 source.n44 source.t17 9.9005
R145 source.n44 source.t14 9.9005
R146 source.n42 source.t15 9.9005
R147 source.n42 source.t27 9.9005
R148 source.n32 source.t6 9.9005
R149 source.n32 source.t3 9.9005
R150 source.n30 source.t4 9.9005
R151 source.n30 source.t5 9.9005
R152 source.n28 source.t12 9.9005
R153 source.n28 source.t1 9.9005
R154 source.n8 source.t9 9.9005
R155 source.n8 source.t2 9.9005
R156 source.n10 source.t0 9.9005
R157 source.n10 source.t13 9.9005
R158 source.n12 source.t8 9.9005
R159 source.n12 source.t10 9.9005
R160 source.n22 source.t21 9.9005
R161 source.n22 source.t24 9.9005
R162 source.n24 source.t22 9.9005
R163 source.n24 source.t16 9.9005
R164 source.n26 source.t26 9.9005
R165 source.n26 source.t19 9.9005
R166 source.n51 source.n49 9.71174
R167 source.n37 source.n35 9.71174
R168 source.n3 source.n1 9.71174
R169 source.n17 source.n15 9.71174
R170 source.n54 source.n53 9.45567
R171 source.n40 source.n39 9.45567
R172 source.n6 source.n5 9.45567
R173 source.n20 source.n19 9.45567
R174 source.n53 source.n52 9.3005
R175 source.n39 source.n38 9.3005
R176 source.n5 source.n4 9.3005
R177 source.n19 source.n18 9.3005
R178 source.n56 source.n7 8.8068
R179 source.n54 source.n48 8.14595
R180 source.n40 source.n34 8.14595
R181 source.n6 source.n0 8.14595
R182 source.n20 source.n14 8.14595
R183 source.n52 source.n51 7.3702
R184 source.n38 source.n37 7.3702
R185 source.n4 source.n3 7.3702
R186 source.n18 source.n17 7.3702
R187 source.n52 source.n48 5.81868
R188 source.n38 source.n34 5.81868
R189 source.n4 source.n0 5.81868
R190 source.n18 source.n14 5.81868
R191 source.n56 source.n55 5.62119
R192 source.n53 source.n49 3.44771
R193 source.n39 source.n35 3.44771
R194 source.n5 source.n1 3.44771
R195 source.n19 source.n15 3.44771
R196 source.n21 source.n13 0.828086
R197 source.n43 source.n41 0.828086
R198 source.n27 source.n25 0.716017
R199 source.n25 source.n23 0.716017
R200 source.n23 source.n21 0.716017
R201 source.n13 source.n11 0.716017
R202 source.n11 source.n9 0.716017
R203 source.n9 source.n7 0.716017
R204 source.n31 source.n29 0.716017
R205 source.n33 source.n31 0.716017
R206 source.n41 source.n33 0.716017
R207 source.n45 source.n43 0.716017
R208 source.n47 source.n45 0.716017
R209 source.n55 source.n47 0.716017
R210 source source.n56 0.188
R211 plus.n4 plus.t2 195.948
R212 plus.n20 plus.t12 195.948
R213 plus.n14 plus.t7 174.966
R214 plus.n13 plus.t13 174.966
R215 plus.n1 plus.t10 174.966
R216 plus.n8 plus.t5 174.966
R217 plus.n7 plus.t11 174.966
R218 plus.n3 plus.t8 174.966
R219 plus.n30 plus.t4 174.966
R220 plus.n29 plus.t0 174.966
R221 plus.n17 plus.t6 174.966
R222 plus.n24 plus.t3 174.966
R223 plus.n23 plus.t9 174.966
R224 plus.n19 plus.t1 174.966
R225 plus.n6 plus.n5 161.3
R226 plus.n7 plus.n2 161.3
R227 plus.n10 plus.n1 161.3
R228 plus.n12 plus.n11 161.3
R229 plus.n13 plus.n0 161.3
R230 plus.n15 plus.n14 161.3
R231 plus.n22 plus.n21 161.3
R232 plus.n23 plus.n18 161.3
R233 plus.n26 plus.n17 161.3
R234 plus.n28 plus.n27 161.3
R235 plus.n29 plus.n16 161.3
R236 plus.n31 plus.n30 161.3
R237 plus.n9 plus.n8 80.6037
R238 plus.n25 plus.n24 80.6037
R239 plus.n5 plus.n4 70.4033
R240 plus.n21 plus.n20 70.4033
R241 plus.n14 plus.n13 48.2005
R242 plus.n8 plus.n1 48.2005
R243 plus.n8 plus.n7 48.2005
R244 plus.n30 plus.n29 48.2005
R245 plus.n24 plus.n17 48.2005
R246 plus.n24 plus.n23 48.2005
R247 plus plus.n31 27.0502
R248 plus.n12 plus.n1 24.8308
R249 plus.n7 plus.n6 24.8308
R250 plus.n28 plus.n17 24.8308
R251 plus.n23 plus.n22 24.8308
R252 plus.n13 plus.n12 23.3702
R253 plus.n6 plus.n3 23.3702
R254 plus.n29 plus.n28 23.3702
R255 plus.n22 plus.n19 23.3702
R256 plus.n4 plus.n3 20.9576
R257 plus.n20 plus.n19 20.9576
R258 plus plus.n15 8.44936
R259 plus.n9 plus.n2 0.285035
R260 plus.n10 plus.n9 0.285035
R261 plus.n26 plus.n25 0.285035
R262 plus.n25 plus.n18 0.285035
R263 plus.n5 plus.n2 0.189894
R264 plus.n11 plus.n10 0.189894
R265 plus.n11 plus.n0 0.189894
R266 plus.n15 plus.n0 0.189894
R267 plus.n31 plus.n16 0.189894
R268 plus.n27 plus.n16 0.189894
R269 plus.n27 plus.n26 0.189894
R270 plus.n21 plus.n18 0.189894
R271 drain_left.n2 drain_left.n0 289.615
R272 drain_left.n15 drain_left.n13 289.615
R273 drain_left.n3 drain_left.n2 185
R274 drain_left.n16 drain_left.n15 185
R275 drain_left.t9 drain_left.n1 167.117
R276 drain_left.t11 drain_left.n14 167.117
R277 drain_left.n11 drain_left.n9 101.511
R278 drain_left.n25 drain_left.n24 100.796
R279 drain_left.n23 drain_left.n22 100.796
R280 drain_left.n21 drain_left.n20 100.796
R281 drain_left.n11 drain_left.n10 100.796
R282 drain_left.n8 drain_left.n7 100.796
R283 drain_left.n2 drain_left.t9 52.3082
R284 drain_left.n15 drain_left.t11 52.3082
R285 drain_left.n8 drain_left.n6 48.8039
R286 drain_left.n21 drain_left.n19 48.8039
R287 drain_left drain_left.n12 23.9055
R288 drain_left.n9 drain_left.t12 9.9005
R289 drain_left.n9 drain_left.t1 9.9005
R290 drain_left.n10 drain_left.t10 9.9005
R291 drain_left.n10 drain_left.t4 9.9005
R292 drain_left.n7 drain_left.t13 9.9005
R293 drain_left.n7 drain_left.t7 9.9005
R294 drain_left.n24 drain_left.t0 9.9005
R295 drain_left.n24 drain_left.t6 9.9005
R296 drain_left.n22 drain_left.t8 9.9005
R297 drain_left.n22 drain_left.t3 9.9005
R298 drain_left.n20 drain_left.t5 9.9005
R299 drain_left.n20 drain_left.t2 9.9005
R300 drain_left.n3 drain_left.n1 9.71174
R301 drain_left.n16 drain_left.n14 9.71174
R302 drain_left.n6 drain_left.n5 9.45567
R303 drain_left.n19 drain_left.n18 9.45567
R304 drain_left.n5 drain_left.n4 9.3005
R305 drain_left.n18 drain_left.n17 9.3005
R306 drain_left.n6 drain_left.n0 8.14595
R307 drain_left.n19 drain_left.n13 8.14595
R308 drain_left.n4 drain_left.n3 7.3702
R309 drain_left.n17 drain_left.n16 7.3702
R310 drain_left drain_left.n25 6.36873
R311 drain_left.n4 drain_left.n0 5.81868
R312 drain_left.n17 drain_left.n13 5.81868
R313 drain_left.n5 drain_left.n1 3.44771
R314 drain_left.n18 drain_left.n14 3.44771
R315 drain_left.n23 drain_left.n21 0.716017
R316 drain_left.n25 drain_left.n23 0.716017
R317 drain_left.n12 drain_left.n8 0.481792
R318 drain_left.n12 drain_left.n11 0.124033
C0 source plus 2.03002f
C1 drain_right minus 1.66163f
C2 source drain_left 6.07827f
C3 drain_left plus 1.86097f
C4 source minus 2.01597f
C5 plus minus 3.8518f
C6 source drain_right 6.07708f
C7 drain_right plus 0.362987f
C8 drain_left minus 0.178852f
C9 drain_left drain_right 1.05573f
C10 drain_right a_n2044_n1288# 4.093f
C11 drain_left a_n2044_n1288# 4.37054f
C12 source a_n2044_n1288# 2.669246f
C13 minus a_n2044_n1288# 7.228437f
C14 plus a_n2044_n1288# 8.157229f
C15 drain_left.n0 a_n2044_n1288# 0.029987f
C16 drain_left.n1 a_n2044_n1288# 0.06635f
C17 drain_left.t9 a_n2044_n1288# 0.049792f
C18 drain_left.n2 a_n2044_n1288# 0.051928f
C19 drain_left.n3 a_n2044_n1288# 0.01674f
C20 drain_left.n4 a_n2044_n1288# 0.01104f
C21 drain_left.n5 a_n2044_n1288# 0.146251f
C22 drain_left.n6 a_n2044_n1288# 0.048333f
C23 drain_left.t13 a_n2044_n1288# 0.032471f
C24 drain_left.t7 a_n2044_n1288# 0.032471f
C25 drain_left.n7 a_n2044_n1288# 0.203991f
C26 drain_left.n8 a_n2044_n1288# 0.322492f
C27 drain_left.t12 a_n2044_n1288# 0.032471f
C28 drain_left.t1 a_n2044_n1288# 0.032471f
C29 drain_left.n9 a_n2044_n1288# 0.205826f
C30 drain_left.t10 a_n2044_n1288# 0.032471f
C31 drain_left.t4 a_n2044_n1288# 0.032471f
C32 drain_left.n10 a_n2044_n1288# 0.203991f
C33 drain_left.n11 a_n2044_n1288# 0.475079f
C34 drain_left.n12 a_n2044_n1288# 0.634511f
C35 drain_left.n13 a_n2044_n1288# 0.029987f
C36 drain_left.n14 a_n2044_n1288# 0.06635f
C37 drain_left.t11 a_n2044_n1288# 0.049792f
C38 drain_left.n15 a_n2044_n1288# 0.051928f
C39 drain_left.n16 a_n2044_n1288# 0.01674f
C40 drain_left.n17 a_n2044_n1288# 0.01104f
C41 drain_left.n18 a_n2044_n1288# 0.146251f
C42 drain_left.n19 a_n2044_n1288# 0.048333f
C43 drain_left.t5 a_n2044_n1288# 0.032471f
C44 drain_left.t2 a_n2044_n1288# 0.032471f
C45 drain_left.n20 a_n2044_n1288# 0.203992f
C46 drain_left.n21 a_n2044_n1288# 0.337007f
C47 drain_left.t8 a_n2044_n1288# 0.032471f
C48 drain_left.t3 a_n2044_n1288# 0.032471f
C49 drain_left.n22 a_n2044_n1288# 0.203992f
C50 drain_left.n23 a_n2044_n1288# 0.251985f
C51 drain_left.t0 a_n2044_n1288# 0.032471f
C52 drain_left.t6 a_n2044_n1288# 0.032471f
C53 drain_left.n24 a_n2044_n1288# 0.203992f
C54 drain_left.n25 a_n2044_n1288# 0.428497f
C55 plus.n0 a_n2044_n1288# 0.037599f
C56 plus.t7 a_n2044_n1288# 0.116433f
C57 plus.t13 a_n2044_n1288# 0.116433f
C58 plus.t10 a_n2044_n1288# 0.116433f
C59 plus.n1 a_n2044_n1288# 0.087812f
C60 plus.n2 a_n2044_n1288# 0.050171f
C61 plus.t5 a_n2044_n1288# 0.116433f
C62 plus.t11 a_n2044_n1288# 0.116433f
C63 plus.t8 a_n2044_n1288# 0.116433f
C64 plus.n3 a_n2044_n1288# 0.08758f
C65 plus.t2 a_n2044_n1288# 0.12542f
C66 plus.n4 a_n2044_n1288# 0.075173f
C67 plus.n5 a_n2044_n1288# 0.123634f
C68 plus.n6 a_n2044_n1288# 0.008532f
C69 plus.n7 a_n2044_n1288# 0.087812f
C70 plus.n8 a_n2044_n1288# 0.092403f
C71 plus.n9 a_n2044_n1288# 0.050053f
C72 plus.n10 a_n2044_n1288# 0.050171f
C73 plus.n11 a_n2044_n1288# 0.037599f
C74 plus.n12 a_n2044_n1288# 0.008532f
C75 plus.n13 a_n2044_n1288# 0.08758f
C76 plus.n14 a_n2044_n1288# 0.083871f
C77 plus.n15 a_n2044_n1288# 0.277466f
C78 plus.n16 a_n2044_n1288# 0.037599f
C79 plus.t4 a_n2044_n1288# 0.116433f
C80 plus.t0 a_n2044_n1288# 0.116433f
C81 plus.t6 a_n2044_n1288# 0.116433f
C82 plus.n17 a_n2044_n1288# 0.087812f
C83 plus.n18 a_n2044_n1288# 0.050171f
C84 plus.t3 a_n2044_n1288# 0.116433f
C85 plus.t9 a_n2044_n1288# 0.116433f
C86 plus.t1 a_n2044_n1288# 0.116433f
C87 plus.n19 a_n2044_n1288# 0.08758f
C88 plus.t12 a_n2044_n1288# 0.12542f
C89 plus.n20 a_n2044_n1288# 0.075173f
C90 plus.n21 a_n2044_n1288# 0.123634f
C91 plus.n22 a_n2044_n1288# 0.008532f
C92 plus.n23 a_n2044_n1288# 0.087812f
C93 plus.n24 a_n2044_n1288# 0.092403f
C94 plus.n25 a_n2044_n1288# 0.050053f
C95 plus.n26 a_n2044_n1288# 0.050171f
C96 plus.n27 a_n2044_n1288# 0.037599f
C97 plus.n28 a_n2044_n1288# 0.008532f
C98 plus.n29 a_n2044_n1288# 0.08758f
C99 plus.n30 a_n2044_n1288# 0.083871f
C100 plus.n31 a_n2044_n1288# 0.903119f
C101 source.n0 a_n2044_n1288# 0.049532f
C102 source.n1 a_n2044_n1288# 0.109594f
C103 source.t7 a_n2044_n1288# 0.082245f
C104 source.n2 a_n2044_n1288# 0.085773f
C105 source.n3 a_n2044_n1288# 0.02765f
C106 source.n4 a_n2044_n1288# 0.018236f
C107 source.n5 a_n2044_n1288# 0.241573f
C108 source.n6 a_n2044_n1288# 0.054298f
C109 source.n7 a_n2044_n1288# 0.54583f
C110 source.t9 a_n2044_n1288# 0.053634f
C111 source.t2 a_n2044_n1288# 0.053634f
C112 source.n8 a_n2044_n1288# 0.286727f
C113 source.n9 a_n2044_n1288# 0.420318f
C114 source.t0 a_n2044_n1288# 0.053634f
C115 source.t13 a_n2044_n1288# 0.053634f
C116 source.n10 a_n2044_n1288# 0.286727f
C117 source.n11 a_n2044_n1288# 0.420318f
C118 source.t8 a_n2044_n1288# 0.053634f
C119 source.t10 a_n2044_n1288# 0.053634f
C120 source.n12 a_n2044_n1288# 0.286727f
C121 source.n13 a_n2044_n1288# 0.432572f
C122 source.n14 a_n2044_n1288# 0.049532f
C123 source.n15 a_n2044_n1288# 0.109594f
C124 source.t18 a_n2044_n1288# 0.082245f
C125 source.n16 a_n2044_n1288# 0.085773f
C126 source.n17 a_n2044_n1288# 0.02765f
C127 source.n18 a_n2044_n1288# 0.018236f
C128 source.n19 a_n2044_n1288# 0.241573f
C129 source.n20 a_n2044_n1288# 0.054298f
C130 source.n21 a_n2044_n1288# 0.196674f
C131 source.t21 a_n2044_n1288# 0.053634f
C132 source.t24 a_n2044_n1288# 0.053634f
C133 source.n22 a_n2044_n1288# 0.286727f
C134 source.n23 a_n2044_n1288# 0.420318f
C135 source.t22 a_n2044_n1288# 0.053634f
C136 source.t16 a_n2044_n1288# 0.053634f
C137 source.n24 a_n2044_n1288# 0.286727f
C138 source.n25 a_n2044_n1288# 0.420318f
C139 source.t26 a_n2044_n1288# 0.053634f
C140 source.t19 a_n2044_n1288# 0.053634f
C141 source.n26 a_n2044_n1288# 0.286727f
C142 source.n27 a_n2044_n1288# 1.18061f
C143 source.t12 a_n2044_n1288# 0.053634f
C144 source.t1 a_n2044_n1288# 0.053634f
C145 source.n28 a_n2044_n1288# 0.286726f
C146 source.n29 a_n2044_n1288# 1.18061f
C147 source.t4 a_n2044_n1288# 0.053634f
C148 source.t5 a_n2044_n1288# 0.053634f
C149 source.n30 a_n2044_n1288# 0.286726f
C150 source.n31 a_n2044_n1288# 0.420319f
C151 source.t6 a_n2044_n1288# 0.053634f
C152 source.t3 a_n2044_n1288# 0.053634f
C153 source.n32 a_n2044_n1288# 0.286726f
C154 source.n33 a_n2044_n1288# 0.420319f
C155 source.n34 a_n2044_n1288# 0.049532f
C156 source.n35 a_n2044_n1288# 0.109594f
C157 source.t11 a_n2044_n1288# 0.082245f
C158 source.n36 a_n2044_n1288# 0.085773f
C159 source.n37 a_n2044_n1288# 0.02765f
C160 source.n38 a_n2044_n1288# 0.018236f
C161 source.n39 a_n2044_n1288# 0.241573f
C162 source.n40 a_n2044_n1288# 0.054298f
C163 source.n41 a_n2044_n1288# 0.196674f
C164 source.t15 a_n2044_n1288# 0.053634f
C165 source.t27 a_n2044_n1288# 0.053634f
C166 source.n42 a_n2044_n1288# 0.286726f
C167 source.n43 a_n2044_n1288# 0.432574f
C168 source.t17 a_n2044_n1288# 0.053634f
C169 source.t14 a_n2044_n1288# 0.053634f
C170 source.n44 a_n2044_n1288# 0.286726f
C171 source.n45 a_n2044_n1288# 0.420319f
C172 source.t20 a_n2044_n1288# 0.053634f
C173 source.t25 a_n2044_n1288# 0.053634f
C174 source.n46 a_n2044_n1288# 0.286726f
C175 source.n47 a_n2044_n1288# 0.420319f
C176 source.n48 a_n2044_n1288# 0.049532f
C177 source.n49 a_n2044_n1288# 0.109594f
C178 source.t23 a_n2044_n1288# 0.082245f
C179 source.n50 a_n2044_n1288# 0.085773f
C180 source.n51 a_n2044_n1288# 0.02765f
C181 source.n52 a_n2044_n1288# 0.018236f
C182 source.n53 a_n2044_n1288# 0.241573f
C183 source.n54 a_n2044_n1288# 0.054298f
C184 source.n55 a_n2044_n1288# 0.364104f
C185 source.n56 a_n2044_n1288# 0.84714f
C186 drain_right.n0 a_n2044_n1288# 0.030387f
C187 drain_right.n1 a_n2044_n1288# 0.067235f
C188 drain_right.t12 a_n2044_n1288# 0.050457f
C189 drain_right.n2 a_n2044_n1288# 0.052621f
C190 drain_right.n3 a_n2044_n1288# 0.016963f
C191 drain_right.n4 a_n2044_n1288# 0.011187f
C192 drain_right.n5 a_n2044_n1288# 0.148204f
C193 drain_right.n6 a_n2044_n1288# 0.048978f
C194 drain_right.t2 a_n2044_n1288# 0.032904f
C195 drain_right.t4 a_n2044_n1288# 0.032904f
C196 drain_right.n7 a_n2044_n1288# 0.206715f
C197 drain_right.n8 a_n2044_n1288# 0.326797f
C198 drain_right.t3 a_n2044_n1288# 0.032904f
C199 drain_right.t6 a_n2044_n1288# 0.032904f
C200 drain_right.n9 a_n2044_n1288# 0.208574f
C201 drain_right.t13 a_n2044_n1288# 0.032904f
C202 drain_right.t0 a_n2044_n1288# 0.032904f
C203 drain_right.n10 a_n2044_n1288# 0.206715f
C204 drain_right.n11 a_n2044_n1288# 0.481422f
C205 drain_right.n12 a_n2044_n1288# 0.602274f
C206 drain_right.t5 a_n2044_n1288# 0.032904f
C207 drain_right.t7 a_n2044_n1288# 0.032904f
C208 drain_right.n13 a_n2044_n1288# 0.208575f
C209 drain_right.t8 a_n2044_n1288# 0.032904f
C210 drain_right.t10 a_n2044_n1288# 0.032904f
C211 drain_right.n14 a_n2044_n1288# 0.206716f
C212 drain_right.n15 a_n2044_n1288# 0.517226f
C213 drain_right.t9 a_n2044_n1288# 0.032904f
C214 drain_right.t1 a_n2044_n1288# 0.032904f
C215 drain_right.n16 a_n2044_n1288# 0.206716f
C216 drain_right.n17 a_n2044_n1288# 0.25535f
C217 drain_right.n18 a_n2044_n1288# 0.030387f
C218 drain_right.n19 a_n2044_n1288# 0.067235f
C219 drain_right.t11 a_n2044_n1288# 0.050457f
C220 drain_right.n20 a_n2044_n1288# 0.052621f
C221 drain_right.n21 a_n2044_n1288# 0.016963f
C222 drain_right.n22 a_n2044_n1288# 0.011187f
C223 drain_right.n23 a_n2044_n1288# 0.148204f
C224 drain_right.n24 a_n2044_n1288# 0.047696f
C225 drain_right.n25 a_n2044_n1288# 0.269996f
C226 minus.n0 a_n2044_n1288# 0.03712f
C227 minus.t5 a_n2044_n1288# 0.114952f
C228 minus.n1 a_n2044_n1288# 0.086695f
C229 minus.n2 a_n2044_n1288# 0.049533f
C230 minus.t3 a_n2044_n1288# 0.114952f
C231 minus.n3 a_n2044_n1288# 0.086466f
C232 minus.t9 a_n2044_n1288# 0.123824f
C233 minus.n4 a_n2044_n1288# 0.074217f
C234 minus.n5 a_n2044_n1288# 0.122061f
C235 minus.n6 a_n2044_n1288# 0.008423f
C236 minus.t6 a_n2044_n1288# 0.114952f
C237 minus.n7 a_n2044_n1288# 0.086695f
C238 minus.t11 a_n2044_n1288# 0.114952f
C239 minus.n8 a_n2044_n1288# 0.091227f
C240 minus.n9 a_n2044_n1288# 0.049417f
C241 minus.n10 a_n2044_n1288# 0.049533f
C242 minus.n11 a_n2044_n1288# 0.03712f
C243 minus.n12 a_n2044_n1288# 0.008423f
C244 minus.t8 a_n2044_n1288# 0.114952f
C245 minus.n13 a_n2044_n1288# 0.086466f
C246 minus.t1 a_n2044_n1288# 0.114952f
C247 minus.n14 a_n2044_n1288# 0.082804f
C248 minus.n15 a_n2044_n1288# 0.935008f
C249 minus.n16 a_n2044_n1288# 0.03712f
C250 minus.t7 a_n2044_n1288# 0.114952f
C251 minus.n17 a_n2044_n1288# 0.086695f
C252 minus.n18 a_n2044_n1288# 0.049533f
C253 minus.t0 a_n2044_n1288# 0.114952f
C254 minus.n19 a_n2044_n1288# 0.086466f
C255 minus.t12 a_n2044_n1288# 0.123824f
C256 minus.n20 a_n2044_n1288# 0.074217f
C257 minus.n21 a_n2044_n1288# 0.122061f
C258 minus.n22 a_n2044_n1288# 0.008423f
C259 minus.t10 a_n2044_n1288# 0.114952f
C260 minus.n23 a_n2044_n1288# 0.086695f
C261 minus.t13 a_n2044_n1288# 0.114952f
C262 minus.n24 a_n2044_n1288# 0.091227f
C263 minus.n25 a_n2044_n1288# 0.049417f
C264 minus.n26 a_n2044_n1288# 0.049533f
C265 minus.n27 a_n2044_n1288# 0.03712f
C266 minus.n28 a_n2044_n1288# 0.008423f
C267 minus.t2 a_n2044_n1288# 0.114952f
C268 minus.n29 a_n2044_n1288# 0.086466f
C269 minus.t4 a_n2044_n1288# 0.114952f
C270 minus.n30 a_n2044_n1288# 0.082804f
C271 minus.n31 a_n2044_n1288# 0.250808f
C272 minus.n32 a_n2044_n1288# 1.15034f
.ends

