* NGSPICE file created from diffpair602.ext - technology: sky130A

.subckt diffpair602 minus drain_right drain_left source plus
X0 drain_left.t5 plus.t0 source.t10 a_n1380_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X1 source.t9 plus.t1 drain_left.t4 a_n1380_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X2 source.t5 minus.t0 drain_right.t5 a_n1380_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X3 drain_left.t3 plus.t2 source.t11 a_n1380_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X4 source.t1 minus.t1 drain_right.t4 a_n1380_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X5 drain_right.t3 minus.t2 source.t3 a_n1380_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X6 drain_right.t2 minus.t3 source.t4 a_n1380_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X7 a_n1380_n4888# a_n1380_n4888# a_n1380_n4888# a_n1380_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.5
X8 a_n1380_n4888# a_n1380_n4888# a_n1380_n4888# a_n1380_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X9 drain_left.t2 plus.t3 source.t7 a_n1380_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.5
X10 a_n1380_n4888# a_n1380_n4888# a_n1380_n4888# a_n1380_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
X11 drain_right.t1 minus.t4 source.t0 a_n1380_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X12 drain_right.t0 minus.t5 source.t2 a_n1380_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X13 source.t8 plus.t4 drain_left.t1 a_n1380_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.5
X14 drain_left.t0 plus.t5 source.t6 a_n1380_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.5
X15 a_n1380_n4888# a_n1380_n4888# a_n1380_n4888# a_n1380_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.5
R0 plus.n0 plus.t2 1069.39
R1 plus.n4 plus.t0 1069.39
R2 plus.n2 plus.t5 1042.57
R3 plus.n1 plus.t4 1042.57
R4 plus.n6 plus.t3 1042.57
R5 plus.n5 plus.t1 1042.57
R6 plus.n3 plus.n2 161.3
R7 plus.n7 plus.n6 161.3
R8 plus.n2 plus.n1 48.2005
R9 plus.n6 plus.n5 48.2005
R10 plus.n3 plus.n0 45.1367
R11 plus.n7 plus.n4 45.1367
R12 plus plus.n7 31.2926
R13 plus plus.n3 15.2069
R14 plus.n1 plus.n0 13.3799
R15 plus.n5 plus.n4 13.3799
R16 source.n0 source.t6 44.1297
R17 source.n3 source.t0 44.1296
R18 source.n11 source.t2 44.1295
R19 source.n8 source.t10 44.1295
R20 source.n2 source.n1 43.1397
R21 source.n5 source.n4 43.1397
R22 source.n10 source.n9 43.1396
R23 source.n7 source.n6 43.1396
R24 source.n7 source.n5 28.7794
R25 source.n12 source.n0 22.4432
R26 source.n12 source.n11 5.62119
R27 source.n9 source.t3 0.9905
R28 source.n9 source.t1 0.9905
R29 source.n6 source.t7 0.9905
R30 source.n6 source.t9 0.9905
R31 source.n1 source.t11 0.9905
R32 source.n1 source.t8 0.9905
R33 source.n4 source.t4 0.9905
R34 source.n4 source.t5 0.9905
R35 source.n3 source.n2 0.828086
R36 source.n10 source.n8 0.828086
R37 source.n5 source.n3 0.716017
R38 source.n2 source.n0 0.716017
R39 source.n8 source.n7 0.716017
R40 source.n11 source.n10 0.716017
R41 source source.n12 0.188
R42 drain_left.n3 drain_left.t3 61.5239
R43 drain_left.n1 drain_left.t2 61.2896
R44 drain_left.n1 drain_left.n0 59.9419
R45 drain_left.n3 drain_left.n2 59.8185
R46 drain_left drain_left.n1 35.3954
R47 drain_left drain_left.n3 6.36873
R48 drain_left.n0 drain_left.t4 0.9905
R49 drain_left.n0 drain_left.t5 0.9905
R50 drain_left.n2 drain_left.t1 0.9905
R51 drain_left.n2 drain_left.t0 0.9905
R52 minus.n0 minus.t4 1069.39
R53 minus.n4 minus.t2 1069.39
R54 minus.n1 minus.t0 1042.57
R55 minus.n2 minus.t3 1042.57
R56 minus.n5 minus.t1 1042.57
R57 minus.n6 minus.t5 1042.57
R58 minus.n3 minus.n2 161.3
R59 minus.n7 minus.n6 161.3
R60 minus.n2 minus.n1 48.2005
R61 minus.n6 minus.n5 48.2005
R62 minus.n3 minus.n0 45.1367
R63 minus.n7 minus.n4 45.1367
R64 minus.n8 minus.n3 40.4418
R65 minus.n1 minus.n0 13.3799
R66 minus.n5 minus.n4 13.3799
R67 minus.n8 minus.n7 6.5327
R68 minus minus.n8 0.188
R69 drain_right.n1 drain_right.t3 61.2896
R70 drain_right.n3 drain_right.t2 60.8084
R71 drain_right.n3 drain_right.n2 60.534
R72 drain_right.n1 drain_right.n0 59.9419
R73 drain_right drain_right.n1 34.8421
R74 drain_right drain_right.n3 6.01097
R75 drain_right.n0 drain_right.t4 0.9905
R76 drain_right.n0 drain_right.t0 0.9905
R77 drain_right.n2 drain_right.t5 0.9905
R78 drain_right.n2 drain_right.t1 0.9905
C0 source drain_right 17.9269f
C1 minus drain_right 5.87159f
C2 minus source 5.15284f
C3 drain_left plus 5.99805f
C4 drain_left drain_right 0.6421f
C5 drain_left source 17.9419f
C6 drain_right plus 0.288098f
C7 minus drain_left 0.171162f
C8 source plus 5.16783f
C9 minus plus 6.35056f
C10 drain_right a_n1380_n4888# 8.47608f
C11 drain_left a_n1380_n4888# 8.677509f
C12 source a_n1380_n4888# 9.139956f
C13 minus a_n1380_n4888# 5.82279f
C14 plus a_n1380_n4888# 8.21609f
C15 drain_right.t3 a_n1380_n4888# 4.5489f
C16 drain_right.t4 a_n1380_n4888# 0.388826f
C17 drain_right.t0 a_n1380_n4888# 0.388826f
C18 drain_right.n0 a_n1380_n4888# 3.55533f
C19 drain_right.n1 a_n1380_n4888# 2.13863f
C20 drain_right.t5 a_n1380_n4888# 0.388826f
C21 drain_right.t1 a_n1380_n4888# 0.388826f
C22 drain_right.n2 a_n1380_n4888# 3.55864f
C23 drain_right.t2 a_n1380_n4888# 4.54636f
C24 drain_right.n3 a_n1380_n4888# 0.88582f
C25 minus.t4 a_n1380_n4888# 1.47222f
C26 minus.n0 a_n1380_n4888# 0.535164f
C27 minus.t0 a_n1380_n4888# 1.45848f
C28 minus.n1 a_n1380_n4888# 0.559569f
C29 minus.t3 a_n1380_n4888# 1.45848f
C30 minus.n2 a_n1380_n4888# 0.547882f
C31 minus.n3 a_n1380_n4888# 2.31619f
C32 minus.t2 a_n1380_n4888# 1.47222f
C33 minus.n4 a_n1380_n4888# 0.535164f
C34 minus.t1 a_n1380_n4888# 1.45848f
C35 minus.n5 a_n1380_n4888# 0.559569f
C36 minus.t5 a_n1380_n4888# 1.45848f
C37 minus.n6 a_n1380_n4888# 0.547882f
C38 minus.n7 a_n1380_n4888# 0.499227f
C39 minus.n8 a_n1380_n4888# 2.58717f
C40 drain_left.t2 a_n1380_n4888# 4.54962f
C41 drain_left.t4 a_n1380_n4888# 0.388887f
C42 drain_left.t5 a_n1380_n4888# 0.388887f
C43 drain_left.n0 a_n1380_n4888# 3.55589f
C44 drain_left.n1 a_n1380_n4888# 2.19057f
C45 drain_left.t3 a_n1380_n4888# 4.55107f
C46 drain_left.t1 a_n1380_n4888# 0.388887f
C47 drain_left.t0 a_n1380_n4888# 0.388887f
C48 drain_left.n2 a_n1380_n4888# 3.55529f
C49 drain_left.n3 a_n1380_n4888# 0.87161f
C50 source.t6 a_n1380_n4888# 4.47504f
C51 source.n0 a_n1380_n4888# 1.92508f
C52 source.t11 a_n1380_n4888# 0.391573f
C53 source.t8 a_n1380_n4888# 0.391573f
C54 source.n1 a_n1380_n4888# 3.50083f
C55 source.n2 a_n1380_n4888# 0.377605f
C56 source.t0 a_n1380_n4888# 4.47505f
C57 source.n3 a_n1380_n4888# 0.471307f
C58 source.t4 a_n1380_n4888# 0.391573f
C59 source.t5 a_n1380_n4888# 0.391573f
C60 source.n4 a_n1380_n4888# 3.50083f
C61 source.n5 a_n1380_n4888# 2.33339f
C62 source.t7 a_n1380_n4888# 0.391573f
C63 source.t9 a_n1380_n4888# 0.391573f
C64 source.n6 a_n1380_n4888# 3.50083f
C65 source.n7 a_n1380_n4888# 2.33339f
C66 source.t10 a_n1380_n4888# 4.475029f
C67 source.n8 a_n1380_n4888# 0.471332f
C68 source.t3 a_n1380_n4888# 0.391573f
C69 source.t1 a_n1380_n4888# 0.391573f
C70 source.n9 a_n1380_n4888# 3.50083f
C71 source.n10 a_n1380_n4888# 0.377598f
C72 source.t2 a_n1380_n4888# 4.475029f
C73 source.n11 a_n1380_n4888# 0.593569f
C74 source.n12 a_n1380_n4888# 2.23895f
C75 plus.t2 a_n1380_n4888# 1.4895f
C76 plus.n0 a_n1380_n4888# 0.541444f
C77 plus.t5 a_n1380_n4888# 1.4756f
C78 plus.t4 a_n1380_n4888# 1.4756f
C79 plus.n1 a_n1380_n4888# 0.566136f
C80 plus.n2 a_n1380_n4888# 0.554312f
C81 plus.n3 a_n1380_n4888# 0.955536f
C82 plus.t0 a_n1380_n4888# 1.4895f
C83 plus.n4 a_n1380_n4888# 0.541444f
C84 plus.t3 a_n1380_n4888# 1.4756f
C85 plus.t1 a_n1380_n4888# 1.4756f
C86 plus.n5 a_n1380_n4888# 0.566135f
C87 plus.n6 a_n1380_n4888# 0.554312f
C88 plus.n7 a_n1380_n4888# 1.87649f
.ends

