* NGSPICE file created from diffpair662.ext - technology: sky130A

.subckt diffpair662 minus drain_right drain_left source plus
X0 source.t11 plus.t0 drain_left.t2 a_n1180_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.25
X1 drain_right.t5 minus.t0 source.t2 a_n1180_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.25
X2 source.t3 minus.t1 drain_right.t4 a_n1180_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.25
X3 drain_left.t3 plus.t1 source.t10 a_n1180_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.25
X4 source.t1 minus.t2 drain_right.t3 a_n1180_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.25
X5 drain_left.t4 plus.t2 source.t9 a_n1180_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.25
X6 drain_left.t1 plus.t3 source.t8 a_n1180_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.25
X7 a_n1180_n5888# a_n1180_n5888# a_n1180_n5888# a_n1180_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.25
X8 drain_right.t2 minus.t3 source.t0 a_n1180_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.25
X9 a_n1180_n5888# a_n1180_n5888# a_n1180_n5888# a_n1180_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.25
X10 drain_right.t1 minus.t4 source.t5 a_n1180_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.25
X11 a_n1180_n5888# a_n1180_n5888# a_n1180_n5888# a_n1180_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.25
X12 source.t7 plus.t4 drain_left.t5 a_n1180_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.25
X13 drain_right.t0 minus.t5 source.t4 a_n1180_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.25
X14 a_n1180_n5888# a_n1180_n5888# a_n1180_n5888# a_n1180_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.25
X15 drain_left.t0 plus.t5 source.t6 a_n1180_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.25
R0 plus.n0 plus.t1 2583.52
R1 plus.n2 plus.t2 2583.52
R2 plus.n4 plus.t5 2583.52
R3 plus.n6 plus.t3 2583.52
R4 plus.n1 plus.t0 2535.32
R5 plus.n5 plus.t4 2535.32
R6 plus.n3 plus.n0 161.489
R7 plus.n7 plus.n4 161.489
R8 plus.n3 plus.n2 161.3
R9 plus.n7 plus.n6 161.3
R10 plus.n1 plus.n0 36.5157
R11 plus.n2 plus.n1 36.5157
R12 plus.n6 plus.n5 36.5157
R13 plus.n5 plus.n4 36.5157
R14 plus plus.n7 32.3816
R15 plus plus.n3 17.0535
R16 drain_left.n134 drain_left.n0 289.615
R17 drain_left.n275 drain_left.n141 289.615
R18 drain_left.n44 drain_left.n43 185
R19 drain_left.n49 drain_left.n48 185
R20 drain_left.n51 drain_left.n50 185
R21 drain_left.n40 drain_left.n39 185
R22 drain_left.n57 drain_left.n56 185
R23 drain_left.n59 drain_left.n58 185
R24 drain_left.n36 drain_left.n35 185
R25 drain_left.n66 drain_left.n65 185
R26 drain_left.n67 drain_left.n34 185
R27 drain_left.n69 drain_left.n68 185
R28 drain_left.n32 drain_left.n31 185
R29 drain_left.n75 drain_left.n74 185
R30 drain_left.n77 drain_left.n76 185
R31 drain_left.n28 drain_left.n27 185
R32 drain_left.n83 drain_left.n82 185
R33 drain_left.n85 drain_left.n84 185
R34 drain_left.n24 drain_left.n23 185
R35 drain_left.n91 drain_left.n90 185
R36 drain_left.n93 drain_left.n92 185
R37 drain_left.n20 drain_left.n19 185
R38 drain_left.n99 drain_left.n98 185
R39 drain_left.n101 drain_left.n100 185
R40 drain_left.n16 drain_left.n15 185
R41 drain_left.n107 drain_left.n106 185
R42 drain_left.n110 drain_left.n109 185
R43 drain_left.n108 drain_left.n12 185
R44 drain_left.n115 drain_left.n11 185
R45 drain_left.n117 drain_left.n116 185
R46 drain_left.n119 drain_left.n118 185
R47 drain_left.n8 drain_left.n7 185
R48 drain_left.n125 drain_left.n124 185
R49 drain_left.n127 drain_left.n126 185
R50 drain_left.n4 drain_left.n3 185
R51 drain_left.n133 drain_left.n132 185
R52 drain_left.n135 drain_left.n134 185
R53 drain_left.n276 drain_left.n275 185
R54 drain_left.n274 drain_left.n273 185
R55 drain_left.n145 drain_left.n144 185
R56 drain_left.n268 drain_left.n267 185
R57 drain_left.n266 drain_left.n265 185
R58 drain_left.n149 drain_left.n148 185
R59 drain_left.n260 drain_left.n259 185
R60 drain_left.n258 drain_left.n257 185
R61 drain_left.n256 drain_left.n152 185
R62 drain_left.n156 drain_left.n153 185
R63 drain_left.n251 drain_left.n250 185
R64 drain_left.n249 drain_left.n248 185
R65 drain_left.n158 drain_left.n157 185
R66 drain_left.n243 drain_left.n242 185
R67 drain_left.n241 drain_left.n240 185
R68 drain_left.n162 drain_left.n161 185
R69 drain_left.n235 drain_left.n234 185
R70 drain_left.n233 drain_left.n232 185
R71 drain_left.n166 drain_left.n165 185
R72 drain_left.n227 drain_left.n226 185
R73 drain_left.n225 drain_left.n224 185
R74 drain_left.n170 drain_left.n169 185
R75 drain_left.n219 drain_left.n218 185
R76 drain_left.n217 drain_left.n216 185
R77 drain_left.n174 drain_left.n173 185
R78 drain_left.n211 drain_left.n210 185
R79 drain_left.n209 drain_left.n176 185
R80 drain_left.n208 drain_left.n207 185
R81 drain_left.n179 drain_left.n177 185
R82 drain_left.n202 drain_left.n201 185
R83 drain_left.n200 drain_left.n199 185
R84 drain_left.n183 drain_left.n182 185
R85 drain_left.n194 drain_left.n193 185
R86 drain_left.n192 drain_left.n191 185
R87 drain_left.n187 drain_left.n186 185
R88 drain_left.n45 drain_left.t1 149.524
R89 drain_left.n188 drain_left.t3 149.524
R90 drain_left.n49 drain_left.n43 104.615
R91 drain_left.n50 drain_left.n49 104.615
R92 drain_left.n50 drain_left.n39 104.615
R93 drain_left.n57 drain_left.n39 104.615
R94 drain_left.n58 drain_left.n57 104.615
R95 drain_left.n58 drain_left.n35 104.615
R96 drain_left.n66 drain_left.n35 104.615
R97 drain_left.n67 drain_left.n66 104.615
R98 drain_left.n68 drain_left.n67 104.615
R99 drain_left.n68 drain_left.n31 104.615
R100 drain_left.n75 drain_left.n31 104.615
R101 drain_left.n76 drain_left.n75 104.615
R102 drain_left.n76 drain_left.n27 104.615
R103 drain_left.n83 drain_left.n27 104.615
R104 drain_left.n84 drain_left.n83 104.615
R105 drain_left.n84 drain_left.n23 104.615
R106 drain_left.n91 drain_left.n23 104.615
R107 drain_left.n92 drain_left.n91 104.615
R108 drain_left.n92 drain_left.n19 104.615
R109 drain_left.n99 drain_left.n19 104.615
R110 drain_left.n100 drain_left.n99 104.615
R111 drain_left.n100 drain_left.n15 104.615
R112 drain_left.n107 drain_left.n15 104.615
R113 drain_left.n109 drain_left.n107 104.615
R114 drain_left.n109 drain_left.n108 104.615
R115 drain_left.n108 drain_left.n11 104.615
R116 drain_left.n117 drain_left.n11 104.615
R117 drain_left.n118 drain_left.n117 104.615
R118 drain_left.n118 drain_left.n7 104.615
R119 drain_left.n125 drain_left.n7 104.615
R120 drain_left.n126 drain_left.n125 104.615
R121 drain_left.n126 drain_left.n3 104.615
R122 drain_left.n133 drain_left.n3 104.615
R123 drain_left.n134 drain_left.n133 104.615
R124 drain_left.n275 drain_left.n274 104.615
R125 drain_left.n274 drain_left.n144 104.615
R126 drain_left.n267 drain_left.n144 104.615
R127 drain_left.n267 drain_left.n266 104.615
R128 drain_left.n266 drain_left.n148 104.615
R129 drain_left.n259 drain_left.n148 104.615
R130 drain_left.n259 drain_left.n258 104.615
R131 drain_left.n258 drain_left.n152 104.615
R132 drain_left.n156 drain_left.n152 104.615
R133 drain_left.n250 drain_left.n156 104.615
R134 drain_left.n250 drain_left.n249 104.615
R135 drain_left.n249 drain_left.n157 104.615
R136 drain_left.n242 drain_left.n157 104.615
R137 drain_left.n242 drain_left.n241 104.615
R138 drain_left.n241 drain_left.n161 104.615
R139 drain_left.n234 drain_left.n161 104.615
R140 drain_left.n234 drain_left.n233 104.615
R141 drain_left.n233 drain_left.n165 104.615
R142 drain_left.n226 drain_left.n165 104.615
R143 drain_left.n226 drain_left.n225 104.615
R144 drain_left.n225 drain_left.n169 104.615
R145 drain_left.n218 drain_left.n169 104.615
R146 drain_left.n218 drain_left.n217 104.615
R147 drain_left.n217 drain_left.n173 104.615
R148 drain_left.n210 drain_left.n173 104.615
R149 drain_left.n210 drain_left.n209 104.615
R150 drain_left.n209 drain_left.n208 104.615
R151 drain_left.n208 drain_left.n177 104.615
R152 drain_left.n201 drain_left.n177 104.615
R153 drain_left.n201 drain_left.n200 104.615
R154 drain_left.n200 drain_left.n182 104.615
R155 drain_left.n193 drain_left.n182 104.615
R156 drain_left.n193 drain_left.n192 104.615
R157 drain_left.n192 drain_left.n186 104.615
R158 drain_left.n140 drain_left.n139 58.7851
R159 drain_left.n281 drain_left.n280 58.7153
R160 drain_left.t1 drain_left.n43 52.3082
R161 drain_left.t3 drain_left.n186 52.3082
R162 drain_left.n281 drain_left.n279 47.8126
R163 drain_left.n140 drain_left.n138 47.6323
R164 drain_left drain_left.n140 38.5906
R165 drain_left.n69 drain_left.n34 13.1884
R166 drain_left.n116 drain_left.n115 13.1884
R167 drain_left.n257 drain_left.n256 13.1884
R168 drain_left.n211 drain_left.n176 13.1884
R169 drain_left.n65 drain_left.n64 12.8005
R170 drain_left.n70 drain_left.n32 12.8005
R171 drain_left.n114 drain_left.n12 12.8005
R172 drain_left.n119 drain_left.n10 12.8005
R173 drain_left.n260 drain_left.n151 12.8005
R174 drain_left.n255 drain_left.n153 12.8005
R175 drain_left.n212 drain_left.n174 12.8005
R176 drain_left.n207 drain_left.n178 12.8005
R177 drain_left.n63 drain_left.n36 12.0247
R178 drain_left.n74 drain_left.n73 12.0247
R179 drain_left.n111 drain_left.n110 12.0247
R180 drain_left.n120 drain_left.n8 12.0247
R181 drain_left.n261 drain_left.n149 12.0247
R182 drain_left.n252 drain_left.n251 12.0247
R183 drain_left.n216 drain_left.n215 12.0247
R184 drain_left.n206 drain_left.n179 12.0247
R185 drain_left.n60 drain_left.n59 11.249
R186 drain_left.n77 drain_left.n30 11.249
R187 drain_left.n106 drain_left.n14 11.249
R188 drain_left.n124 drain_left.n123 11.249
R189 drain_left.n265 drain_left.n264 11.249
R190 drain_left.n248 drain_left.n155 11.249
R191 drain_left.n219 drain_left.n172 11.249
R192 drain_left.n203 drain_left.n202 11.249
R193 drain_left.n56 drain_left.n38 10.4732
R194 drain_left.n78 drain_left.n28 10.4732
R195 drain_left.n105 drain_left.n16 10.4732
R196 drain_left.n127 drain_left.n6 10.4732
R197 drain_left.n268 drain_left.n147 10.4732
R198 drain_left.n247 drain_left.n158 10.4732
R199 drain_left.n220 drain_left.n170 10.4732
R200 drain_left.n199 drain_left.n181 10.4732
R201 drain_left.n45 drain_left.n44 10.2747
R202 drain_left.n188 drain_left.n187 10.2747
R203 drain_left.n55 drain_left.n40 9.69747
R204 drain_left.n82 drain_left.n81 9.69747
R205 drain_left.n102 drain_left.n101 9.69747
R206 drain_left.n128 drain_left.n4 9.69747
R207 drain_left.n269 drain_left.n145 9.69747
R208 drain_left.n244 drain_left.n243 9.69747
R209 drain_left.n224 drain_left.n223 9.69747
R210 drain_left.n198 drain_left.n183 9.69747
R211 drain_left.n138 drain_left.n137 9.45567
R212 drain_left.n279 drain_left.n278 9.45567
R213 drain_left.n2 drain_left.n1 9.3005
R214 drain_left.n131 drain_left.n130 9.3005
R215 drain_left.n129 drain_left.n128 9.3005
R216 drain_left.n6 drain_left.n5 9.3005
R217 drain_left.n123 drain_left.n122 9.3005
R218 drain_left.n121 drain_left.n120 9.3005
R219 drain_left.n10 drain_left.n9 9.3005
R220 drain_left.n89 drain_left.n88 9.3005
R221 drain_left.n87 drain_left.n86 9.3005
R222 drain_left.n26 drain_left.n25 9.3005
R223 drain_left.n81 drain_left.n80 9.3005
R224 drain_left.n79 drain_left.n78 9.3005
R225 drain_left.n30 drain_left.n29 9.3005
R226 drain_left.n73 drain_left.n72 9.3005
R227 drain_left.n71 drain_left.n70 9.3005
R228 drain_left.n47 drain_left.n46 9.3005
R229 drain_left.n42 drain_left.n41 9.3005
R230 drain_left.n53 drain_left.n52 9.3005
R231 drain_left.n55 drain_left.n54 9.3005
R232 drain_left.n38 drain_left.n37 9.3005
R233 drain_left.n61 drain_left.n60 9.3005
R234 drain_left.n63 drain_left.n62 9.3005
R235 drain_left.n64 drain_left.n33 9.3005
R236 drain_left.n22 drain_left.n21 9.3005
R237 drain_left.n95 drain_left.n94 9.3005
R238 drain_left.n97 drain_left.n96 9.3005
R239 drain_left.n18 drain_left.n17 9.3005
R240 drain_left.n103 drain_left.n102 9.3005
R241 drain_left.n105 drain_left.n104 9.3005
R242 drain_left.n14 drain_left.n13 9.3005
R243 drain_left.n112 drain_left.n111 9.3005
R244 drain_left.n114 drain_left.n113 9.3005
R245 drain_left.n137 drain_left.n136 9.3005
R246 drain_left.n190 drain_left.n189 9.3005
R247 drain_left.n185 drain_left.n184 9.3005
R248 drain_left.n196 drain_left.n195 9.3005
R249 drain_left.n198 drain_left.n197 9.3005
R250 drain_left.n181 drain_left.n180 9.3005
R251 drain_left.n204 drain_left.n203 9.3005
R252 drain_left.n206 drain_left.n205 9.3005
R253 drain_left.n178 drain_left.n175 9.3005
R254 drain_left.n237 drain_left.n236 9.3005
R255 drain_left.n239 drain_left.n238 9.3005
R256 drain_left.n160 drain_left.n159 9.3005
R257 drain_left.n245 drain_left.n244 9.3005
R258 drain_left.n247 drain_left.n246 9.3005
R259 drain_left.n155 drain_left.n154 9.3005
R260 drain_left.n253 drain_left.n252 9.3005
R261 drain_left.n255 drain_left.n254 9.3005
R262 drain_left.n278 drain_left.n277 9.3005
R263 drain_left.n143 drain_left.n142 9.3005
R264 drain_left.n272 drain_left.n271 9.3005
R265 drain_left.n270 drain_left.n269 9.3005
R266 drain_left.n147 drain_left.n146 9.3005
R267 drain_left.n264 drain_left.n263 9.3005
R268 drain_left.n262 drain_left.n261 9.3005
R269 drain_left.n151 drain_left.n150 9.3005
R270 drain_left.n164 drain_left.n163 9.3005
R271 drain_left.n231 drain_left.n230 9.3005
R272 drain_left.n229 drain_left.n228 9.3005
R273 drain_left.n168 drain_left.n167 9.3005
R274 drain_left.n223 drain_left.n222 9.3005
R275 drain_left.n221 drain_left.n220 9.3005
R276 drain_left.n172 drain_left.n171 9.3005
R277 drain_left.n215 drain_left.n214 9.3005
R278 drain_left.n213 drain_left.n212 9.3005
R279 drain_left.n52 drain_left.n51 8.92171
R280 drain_left.n85 drain_left.n26 8.92171
R281 drain_left.n98 drain_left.n18 8.92171
R282 drain_left.n132 drain_left.n131 8.92171
R283 drain_left.n273 drain_left.n272 8.92171
R284 drain_left.n240 drain_left.n160 8.92171
R285 drain_left.n227 drain_left.n168 8.92171
R286 drain_left.n195 drain_left.n194 8.92171
R287 drain_left.n48 drain_left.n42 8.14595
R288 drain_left.n86 drain_left.n24 8.14595
R289 drain_left.n97 drain_left.n20 8.14595
R290 drain_left.n135 drain_left.n2 8.14595
R291 drain_left.n276 drain_left.n143 8.14595
R292 drain_left.n239 drain_left.n162 8.14595
R293 drain_left.n228 drain_left.n166 8.14595
R294 drain_left.n191 drain_left.n185 8.14595
R295 drain_left.n47 drain_left.n44 7.3702
R296 drain_left.n90 drain_left.n89 7.3702
R297 drain_left.n94 drain_left.n93 7.3702
R298 drain_left.n136 drain_left.n0 7.3702
R299 drain_left.n277 drain_left.n141 7.3702
R300 drain_left.n236 drain_left.n235 7.3702
R301 drain_left.n232 drain_left.n231 7.3702
R302 drain_left.n190 drain_left.n187 7.3702
R303 drain_left.n90 drain_left.n22 6.59444
R304 drain_left.n93 drain_left.n22 6.59444
R305 drain_left.n138 drain_left.n0 6.59444
R306 drain_left.n279 drain_left.n141 6.59444
R307 drain_left.n235 drain_left.n164 6.59444
R308 drain_left.n232 drain_left.n164 6.59444
R309 drain_left drain_left.n281 6.15322
R310 drain_left.n48 drain_left.n47 5.81868
R311 drain_left.n89 drain_left.n24 5.81868
R312 drain_left.n94 drain_left.n20 5.81868
R313 drain_left.n136 drain_left.n135 5.81868
R314 drain_left.n277 drain_left.n276 5.81868
R315 drain_left.n236 drain_left.n162 5.81868
R316 drain_left.n231 drain_left.n166 5.81868
R317 drain_left.n191 drain_left.n190 5.81868
R318 drain_left.n51 drain_left.n42 5.04292
R319 drain_left.n86 drain_left.n85 5.04292
R320 drain_left.n98 drain_left.n97 5.04292
R321 drain_left.n132 drain_left.n2 5.04292
R322 drain_left.n273 drain_left.n143 5.04292
R323 drain_left.n240 drain_left.n239 5.04292
R324 drain_left.n228 drain_left.n227 5.04292
R325 drain_left.n194 drain_left.n185 5.04292
R326 drain_left.n52 drain_left.n40 4.26717
R327 drain_left.n82 drain_left.n26 4.26717
R328 drain_left.n101 drain_left.n18 4.26717
R329 drain_left.n131 drain_left.n4 4.26717
R330 drain_left.n272 drain_left.n145 4.26717
R331 drain_left.n243 drain_left.n160 4.26717
R332 drain_left.n224 drain_left.n168 4.26717
R333 drain_left.n195 drain_left.n183 4.26717
R334 drain_left.n56 drain_left.n55 3.49141
R335 drain_left.n81 drain_left.n28 3.49141
R336 drain_left.n102 drain_left.n16 3.49141
R337 drain_left.n128 drain_left.n127 3.49141
R338 drain_left.n269 drain_left.n268 3.49141
R339 drain_left.n244 drain_left.n158 3.49141
R340 drain_left.n223 drain_left.n170 3.49141
R341 drain_left.n199 drain_left.n198 3.49141
R342 drain_left.n189 drain_left.n188 2.84303
R343 drain_left.n46 drain_left.n45 2.84303
R344 drain_left.n59 drain_left.n38 2.71565
R345 drain_left.n78 drain_left.n77 2.71565
R346 drain_left.n106 drain_left.n105 2.71565
R347 drain_left.n124 drain_left.n6 2.71565
R348 drain_left.n265 drain_left.n147 2.71565
R349 drain_left.n248 drain_left.n247 2.71565
R350 drain_left.n220 drain_left.n219 2.71565
R351 drain_left.n202 drain_left.n181 2.71565
R352 drain_left.n60 drain_left.n36 1.93989
R353 drain_left.n74 drain_left.n30 1.93989
R354 drain_left.n110 drain_left.n14 1.93989
R355 drain_left.n123 drain_left.n8 1.93989
R356 drain_left.n264 drain_left.n149 1.93989
R357 drain_left.n251 drain_left.n155 1.93989
R358 drain_left.n216 drain_left.n172 1.93989
R359 drain_left.n203 drain_left.n179 1.93989
R360 drain_left.n65 drain_left.n63 1.16414
R361 drain_left.n73 drain_left.n32 1.16414
R362 drain_left.n111 drain_left.n12 1.16414
R363 drain_left.n120 drain_left.n119 1.16414
R364 drain_left.n261 drain_left.n260 1.16414
R365 drain_left.n252 drain_left.n153 1.16414
R366 drain_left.n215 drain_left.n174 1.16414
R367 drain_left.n207 drain_left.n206 1.16414
R368 drain_left.n139 drain_left.t5 0.7925
R369 drain_left.n139 drain_left.t0 0.7925
R370 drain_left.n280 drain_left.t2 0.7925
R371 drain_left.n280 drain_left.t4 0.7925
R372 drain_left.n64 drain_left.n34 0.388379
R373 drain_left.n70 drain_left.n69 0.388379
R374 drain_left.n115 drain_left.n114 0.388379
R375 drain_left.n116 drain_left.n10 0.388379
R376 drain_left.n257 drain_left.n151 0.388379
R377 drain_left.n256 drain_left.n255 0.388379
R378 drain_left.n212 drain_left.n211 0.388379
R379 drain_left.n178 drain_left.n176 0.388379
R380 drain_left.n46 drain_left.n41 0.155672
R381 drain_left.n53 drain_left.n41 0.155672
R382 drain_left.n54 drain_left.n53 0.155672
R383 drain_left.n54 drain_left.n37 0.155672
R384 drain_left.n61 drain_left.n37 0.155672
R385 drain_left.n62 drain_left.n61 0.155672
R386 drain_left.n62 drain_left.n33 0.155672
R387 drain_left.n71 drain_left.n33 0.155672
R388 drain_left.n72 drain_left.n71 0.155672
R389 drain_left.n72 drain_left.n29 0.155672
R390 drain_left.n79 drain_left.n29 0.155672
R391 drain_left.n80 drain_left.n79 0.155672
R392 drain_left.n80 drain_left.n25 0.155672
R393 drain_left.n87 drain_left.n25 0.155672
R394 drain_left.n88 drain_left.n87 0.155672
R395 drain_left.n88 drain_left.n21 0.155672
R396 drain_left.n95 drain_left.n21 0.155672
R397 drain_left.n96 drain_left.n95 0.155672
R398 drain_left.n96 drain_left.n17 0.155672
R399 drain_left.n103 drain_left.n17 0.155672
R400 drain_left.n104 drain_left.n103 0.155672
R401 drain_left.n104 drain_left.n13 0.155672
R402 drain_left.n112 drain_left.n13 0.155672
R403 drain_left.n113 drain_left.n112 0.155672
R404 drain_left.n113 drain_left.n9 0.155672
R405 drain_left.n121 drain_left.n9 0.155672
R406 drain_left.n122 drain_left.n121 0.155672
R407 drain_left.n122 drain_left.n5 0.155672
R408 drain_left.n129 drain_left.n5 0.155672
R409 drain_left.n130 drain_left.n129 0.155672
R410 drain_left.n130 drain_left.n1 0.155672
R411 drain_left.n137 drain_left.n1 0.155672
R412 drain_left.n278 drain_left.n142 0.155672
R413 drain_left.n271 drain_left.n142 0.155672
R414 drain_left.n271 drain_left.n270 0.155672
R415 drain_left.n270 drain_left.n146 0.155672
R416 drain_left.n263 drain_left.n146 0.155672
R417 drain_left.n263 drain_left.n262 0.155672
R418 drain_left.n262 drain_left.n150 0.155672
R419 drain_left.n254 drain_left.n150 0.155672
R420 drain_left.n254 drain_left.n253 0.155672
R421 drain_left.n253 drain_left.n154 0.155672
R422 drain_left.n246 drain_left.n154 0.155672
R423 drain_left.n246 drain_left.n245 0.155672
R424 drain_left.n245 drain_left.n159 0.155672
R425 drain_left.n238 drain_left.n159 0.155672
R426 drain_left.n238 drain_left.n237 0.155672
R427 drain_left.n237 drain_left.n163 0.155672
R428 drain_left.n230 drain_left.n163 0.155672
R429 drain_left.n230 drain_left.n229 0.155672
R430 drain_left.n229 drain_left.n167 0.155672
R431 drain_left.n222 drain_left.n167 0.155672
R432 drain_left.n222 drain_left.n221 0.155672
R433 drain_left.n221 drain_left.n171 0.155672
R434 drain_left.n214 drain_left.n171 0.155672
R435 drain_left.n214 drain_left.n213 0.155672
R436 drain_left.n213 drain_left.n175 0.155672
R437 drain_left.n205 drain_left.n175 0.155672
R438 drain_left.n205 drain_left.n204 0.155672
R439 drain_left.n204 drain_left.n180 0.155672
R440 drain_left.n197 drain_left.n180 0.155672
R441 drain_left.n197 drain_left.n196 0.155672
R442 drain_left.n196 drain_left.n184 0.155672
R443 drain_left.n189 drain_left.n184 0.155672
R444 source.n562 source.n428 289.615
R445 source.n420 source.n286 289.615
R446 source.n134 source.n0 289.615
R447 source.n276 source.n142 289.615
R448 source.n472 source.n471 185
R449 source.n477 source.n476 185
R450 source.n479 source.n478 185
R451 source.n468 source.n467 185
R452 source.n485 source.n484 185
R453 source.n487 source.n486 185
R454 source.n464 source.n463 185
R455 source.n494 source.n493 185
R456 source.n495 source.n462 185
R457 source.n497 source.n496 185
R458 source.n460 source.n459 185
R459 source.n503 source.n502 185
R460 source.n505 source.n504 185
R461 source.n456 source.n455 185
R462 source.n511 source.n510 185
R463 source.n513 source.n512 185
R464 source.n452 source.n451 185
R465 source.n519 source.n518 185
R466 source.n521 source.n520 185
R467 source.n448 source.n447 185
R468 source.n527 source.n526 185
R469 source.n529 source.n528 185
R470 source.n444 source.n443 185
R471 source.n535 source.n534 185
R472 source.n538 source.n537 185
R473 source.n536 source.n440 185
R474 source.n543 source.n439 185
R475 source.n545 source.n544 185
R476 source.n547 source.n546 185
R477 source.n436 source.n435 185
R478 source.n553 source.n552 185
R479 source.n555 source.n554 185
R480 source.n432 source.n431 185
R481 source.n561 source.n560 185
R482 source.n563 source.n562 185
R483 source.n330 source.n329 185
R484 source.n335 source.n334 185
R485 source.n337 source.n336 185
R486 source.n326 source.n325 185
R487 source.n343 source.n342 185
R488 source.n345 source.n344 185
R489 source.n322 source.n321 185
R490 source.n352 source.n351 185
R491 source.n353 source.n320 185
R492 source.n355 source.n354 185
R493 source.n318 source.n317 185
R494 source.n361 source.n360 185
R495 source.n363 source.n362 185
R496 source.n314 source.n313 185
R497 source.n369 source.n368 185
R498 source.n371 source.n370 185
R499 source.n310 source.n309 185
R500 source.n377 source.n376 185
R501 source.n379 source.n378 185
R502 source.n306 source.n305 185
R503 source.n385 source.n384 185
R504 source.n387 source.n386 185
R505 source.n302 source.n301 185
R506 source.n393 source.n392 185
R507 source.n396 source.n395 185
R508 source.n394 source.n298 185
R509 source.n401 source.n297 185
R510 source.n403 source.n402 185
R511 source.n405 source.n404 185
R512 source.n294 source.n293 185
R513 source.n411 source.n410 185
R514 source.n413 source.n412 185
R515 source.n290 source.n289 185
R516 source.n419 source.n418 185
R517 source.n421 source.n420 185
R518 source.n135 source.n134 185
R519 source.n133 source.n132 185
R520 source.n4 source.n3 185
R521 source.n127 source.n126 185
R522 source.n125 source.n124 185
R523 source.n8 source.n7 185
R524 source.n119 source.n118 185
R525 source.n117 source.n116 185
R526 source.n115 source.n11 185
R527 source.n15 source.n12 185
R528 source.n110 source.n109 185
R529 source.n108 source.n107 185
R530 source.n17 source.n16 185
R531 source.n102 source.n101 185
R532 source.n100 source.n99 185
R533 source.n21 source.n20 185
R534 source.n94 source.n93 185
R535 source.n92 source.n91 185
R536 source.n25 source.n24 185
R537 source.n86 source.n85 185
R538 source.n84 source.n83 185
R539 source.n29 source.n28 185
R540 source.n78 source.n77 185
R541 source.n76 source.n75 185
R542 source.n33 source.n32 185
R543 source.n70 source.n69 185
R544 source.n68 source.n35 185
R545 source.n67 source.n66 185
R546 source.n38 source.n36 185
R547 source.n61 source.n60 185
R548 source.n59 source.n58 185
R549 source.n42 source.n41 185
R550 source.n53 source.n52 185
R551 source.n51 source.n50 185
R552 source.n46 source.n45 185
R553 source.n277 source.n276 185
R554 source.n275 source.n274 185
R555 source.n146 source.n145 185
R556 source.n269 source.n268 185
R557 source.n267 source.n266 185
R558 source.n150 source.n149 185
R559 source.n261 source.n260 185
R560 source.n259 source.n258 185
R561 source.n257 source.n153 185
R562 source.n157 source.n154 185
R563 source.n252 source.n251 185
R564 source.n250 source.n249 185
R565 source.n159 source.n158 185
R566 source.n244 source.n243 185
R567 source.n242 source.n241 185
R568 source.n163 source.n162 185
R569 source.n236 source.n235 185
R570 source.n234 source.n233 185
R571 source.n167 source.n166 185
R572 source.n228 source.n227 185
R573 source.n226 source.n225 185
R574 source.n171 source.n170 185
R575 source.n220 source.n219 185
R576 source.n218 source.n217 185
R577 source.n175 source.n174 185
R578 source.n212 source.n211 185
R579 source.n210 source.n177 185
R580 source.n209 source.n208 185
R581 source.n180 source.n178 185
R582 source.n203 source.n202 185
R583 source.n201 source.n200 185
R584 source.n184 source.n183 185
R585 source.n195 source.n194 185
R586 source.n193 source.n192 185
R587 source.n188 source.n187 185
R588 source.n473 source.t4 149.524
R589 source.n331 source.t6 149.524
R590 source.n47 source.t9 149.524
R591 source.n189 source.t5 149.524
R592 source.n477 source.n471 104.615
R593 source.n478 source.n477 104.615
R594 source.n478 source.n467 104.615
R595 source.n485 source.n467 104.615
R596 source.n486 source.n485 104.615
R597 source.n486 source.n463 104.615
R598 source.n494 source.n463 104.615
R599 source.n495 source.n494 104.615
R600 source.n496 source.n495 104.615
R601 source.n496 source.n459 104.615
R602 source.n503 source.n459 104.615
R603 source.n504 source.n503 104.615
R604 source.n504 source.n455 104.615
R605 source.n511 source.n455 104.615
R606 source.n512 source.n511 104.615
R607 source.n512 source.n451 104.615
R608 source.n519 source.n451 104.615
R609 source.n520 source.n519 104.615
R610 source.n520 source.n447 104.615
R611 source.n527 source.n447 104.615
R612 source.n528 source.n527 104.615
R613 source.n528 source.n443 104.615
R614 source.n535 source.n443 104.615
R615 source.n537 source.n535 104.615
R616 source.n537 source.n536 104.615
R617 source.n536 source.n439 104.615
R618 source.n545 source.n439 104.615
R619 source.n546 source.n545 104.615
R620 source.n546 source.n435 104.615
R621 source.n553 source.n435 104.615
R622 source.n554 source.n553 104.615
R623 source.n554 source.n431 104.615
R624 source.n561 source.n431 104.615
R625 source.n562 source.n561 104.615
R626 source.n335 source.n329 104.615
R627 source.n336 source.n335 104.615
R628 source.n336 source.n325 104.615
R629 source.n343 source.n325 104.615
R630 source.n344 source.n343 104.615
R631 source.n344 source.n321 104.615
R632 source.n352 source.n321 104.615
R633 source.n353 source.n352 104.615
R634 source.n354 source.n353 104.615
R635 source.n354 source.n317 104.615
R636 source.n361 source.n317 104.615
R637 source.n362 source.n361 104.615
R638 source.n362 source.n313 104.615
R639 source.n369 source.n313 104.615
R640 source.n370 source.n369 104.615
R641 source.n370 source.n309 104.615
R642 source.n377 source.n309 104.615
R643 source.n378 source.n377 104.615
R644 source.n378 source.n305 104.615
R645 source.n385 source.n305 104.615
R646 source.n386 source.n385 104.615
R647 source.n386 source.n301 104.615
R648 source.n393 source.n301 104.615
R649 source.n395 source.n393 104.615
R650 source.n395 source.n394 104.615
R651 source.n394 source.n297 104.615
R652 source.n403 source.n297 104.615
R653 source.n404 source.n403 104.615
R654 source.n404 source.n293 104.615
R655 source.n411 source.n293 104.615
R656 source.n412 source.n411 104.615
R657 source.n412 source.n289 104.615
R658 source.n419 source.n289 104.615
R659 source.n420 source.n419 104.615
R660 source.n134 source.n133 104.615
R661 source.n133 source.n3 104.615
R662 source.n126 source.n3 104.615
R663 source.n126 source.n125 104.615
R664 source.n125 source.n7 104.615
R665 source.n118 source.n7 104.615
R666 source.n118 source.n117 104.615
R667 source.n117 source.n11 104.615
R668 source.n15 source.n11 104.615
R669 source.n109 source.n15 104.615
R670 source.n109 source.n108 104.615
R671 source.n108 source.n16 104.615
R672 source.n101 source.n16 104.615
R673 source.n101 source.n100 104.615
R674 source.n100 source.n20 104.615
R675 source.n93 source.n20 104.615
R676 source.n93 source.n92 104.615
R677 source.n92 source.n24 104.615
R678 source.n85 source.n24 104.615
R679 source.n85 source.n84 104.615
R680 source.n84 source.n28 104.615
R681 source.n77 source.n28 104.615
R682 source.n77 source.n76 104.615
R683 source.n76 source.n32 104.615
R684 source.n69 source.n32 104.615
R685 source.n69 source.n68 104.615
R686 source.n68 source.n67 104.615
R687 source.n67 source.n36 104.615
R688 source.n60 source.n36 104.615
R689 source.n60 source.n59 104.615
R690 source.n59 source.n41 104.615
R691 source.n52 source.n41 104.615
R692 source.n52 source.n51 104.615
R693 source.n51 source.n45 104.615
R694 source.n276 source.n275 104.615
R695 source.n275 source.n145 104.615
R696 source.n268 source.n145 104.615
R697 source.n268 source.n267 104.615
R698 source.n267 source.n149 104.615
R699 source.n260 source.n149 104.615
R700 source.n260 source.n259 104.615
R701 source.n259 source.n153 104.615
R702 source.n157 source.n153 104.615
R703 source.n251 source.n157 104.615
R704 source.n251 source.n250 104.615
R705 source.n250 source.n158 104.615
R706 source.n243 source.n158 104.615
R707 source.n243 source.n242 104.615
R708 source.n242 source.n162 104.615
R709 source.n235 source.n162 104.615
R710 source.n235 source.n234 104.615
R711 source.n234 source.n166 104.615
R712 source.n227 source.n166 104.615
R713 source.n227 source.n226 104.615
R714 source.n226 source.n170 104.615
R715 source.n219 source.n170 104.615
R716 source.n219 source.n218 104.615
R717 source.n218 source.n174 104.615
R718 source.n211 source.n174 104.615
R719 source.n211 source.n210 104.615
R720 source.n210 source.n209 104.615
R721 source.n209 source.n178 104.615
R722 source.n202 source.n178 104.615
R723 source.n202 source.n201 104.615
R724 source.n201 source.n183 104.615
R725 source.n194 source.n183 104.615
R726 source.n194 source.n193 104.615
R727 source.n193 source.n187 104.615
R728 source.t4 source.n471 52.3082
R729 source.t6 source.n329 52.3082
R730 source.t9 source.n45 52.3082
R731 source.t5 source.n187 52.3082
R732 source.n427 source.n426 42.0366
R733 source.n285 source.n284 42.0366
R734 source.n141 source.n140 42.0366
R735 source.n283 source.n282 42.0366
R736 source.n285 source.n283 32.1362
R737 source.n567 source.n566 30.6338
R738 source.n425 source.n424 30.6338
R739 source.n139 source.n138 30.6338
R740 source.n281 source.n280 30.6338
R741 source.n568 source.n139 26.1233
R742 source.n497 source.n462 13.1884
R743 source.n544 source.n543 13.1884
R744 source.n355 source.n320 13.1884
R745 source.n402 source.n401 13.1884
R746 source.n116 source.n115 13.1884
R747 source.n70 source.n35 13.1884
R748 source.n258 source.n257 13.1884
R749 source.n212 source.n177 13.1884
R750 source.n493 source.n492 12.8005
R751 source.n498 source.n460 12.8005
R752 source.n542 source.n440 12.8005
R753 source.n547 source.n438 12.8005
R754 source.n351 source.n350 12.8005
R755 source.n356 source.n318 12.8005
R756 source.n400 source.n298 12.8005
R757 source.n405 source.n296 12.8005
R758 source.n119 source.n10 12.8005
R759 source.n114 source.n12 12.8005
R760 source.n71 source.n33 12.8005
R761 source.n66 source.n37 12.8005
R762 source.n261 source.n152 12.8005
R763 source.n256 source.n154 12.8005
R764 source.n213 source.n175 12.8005
R765 source.n208 source.n179 12.8005
R766 source.n491 source.n464 12.0247
R767 source.n502 source.n501 12.0247
R768 source.n539 source.n538 12.0247
R769 source.n548 source.n436 12.0247
R770 source.n349 source.n322 12.0247
R771 source.n360 source.n359 12.0247
R772 source.n397 source.n396 12.0247
R773 source.n406 source.n294 12.0247
R774 source.n120 source.n8 12.0247
R775 source.n111 source.n110 12.0247
R776 source.n75 source.n74 12.0247
R777 source.n65 source.n38 12.0247
R778 source.n262 source.n150 12.0247
R779 source.n253 source.n252 12.0247
R780 source.n217 source.n216 12.0247
R781 source.n207 source.n180 12.0247
R782 source.n488 source.n487 11.249
R783 source.n505 source.n458 11.249
R784 source.n534 source.n442 11.249
R785 source.n552 source.n551 11.249
R786 source.n346 source.n345 11.249
R787 source.n363 source.n316 11.249
R788 source.n392 source.n300 11.249
R789 source.n410 source.n409 11.249
R790 source.n124 source.n123 11.249
R791 source.n107 source.n14 11.249
R792 source.n78 source.n31 11.249
R793 source.n62 source.n61 11.249
R794 source.n266 source.n265 11.249
R795 source.n249 source.n156 11.249
R796 source.n220 source.n173 11.249
R797 source.n204 source.n203 11.249
R798 source.n484 source.n466 10.4732
R799 source.n506 source.n456 10.4732
R800 source.n533 source.n444 10.4732
R801 source.n555 source.n434 10.4732
R802 source.n342 source.n324 10.4732
R803 source.n364 source.n314 10.4732
R804 source.n391 source.n302 10.4732
R805 source.n413 source.n292 10.4732
R806 source.n127 source.n6 10.4732
R807 source.n106 source.n17 10.4732
R808 source.n79 source.n29 10.4732
R809 source.n58 source.n40 10.4732
R810 source.n269 source.n148 10.4732
R811 source.n248 source.n159 10.4732
R812 source.n221 source.n171 10.4732
R813 source.n200 source.n182 10.4732
R814 source.n473 source.n472 10.2747
R815 source.n331 source.n330 10.2747
R816 source.n47 source.n46 10.2747
R817 source.n189 source.n188 10.2747
R818 source.n483 source.n468 9.69747
R819 source.n510 source.n509 9.69747
R820 source.n530 source.n529 9.69747
R821 source.n556 source.n432 9.69747
R822 source.n341 source.n326 9.69747
R823 source.n368 source.n367 9.69747
R824 source.n388 source.n387 9.69747
R825 source.n414 source.n290 9.69747
R826 source.n128 source.n4 9.69747
R827 source.n103 source.n102 9.69747
R828 source.n83 source.n82 9.69747
R829 source.n57 source.n42 9.69747
R830 source.n270 source.n146 9.69747
R831 source.n245 source.n244 9.69747
R832 source.n225 source.n224 9.69747
R833 source.n199 source.n184 9.69747
R834 source.n566 source.n565 9.45567
R835 source.n424 source.n423 9.45567
R836 source.n138 source.n137 9.45567
R837 source.n280 source.n279 9.45567
R838 source.n430 source.n429 9.3005
R839 source.n559 source.n558 9.3005
R840 source.n557 source.n556 9.3005
R841 source.n434 source.n433 9.3005
R842 source.n551 source.n550 9.3005
R843 source.n549 source.n548 9.3005
R844 source.n438 source.n437 9.3005
R845 source.n517 source.n516 9.3005
R846 source.n515 source.n514 9.3005
R847 source.n454 source.n453 9.3005
R848 source.n509 source.n508 9.3005
R849 source.n507 source.n506 9.3005
R850 source.n458 source.n457 9.3005
R851 source.n501 source.n500 9.3005
R852 source.n499 source.n498 9.3005
R853 source.n475 source.n474 9.3005
R854 source.n470 source.n469 9.3005
R855 source.n481 source.n480 9.3005
R856 source.n483 source.n482 9.3005
R857 source.n466 source.n465 9.3005
R858 source.n489 source.n488 9.3005
R859 source.n491 source.n490 9.3005
R860 source.n492 source.n461 9.3005
R861 source.n450 source.n449 9.3005
R862 source.n523 source.n522 9.3005
R863 source.n525 source.n524 9.3005
R864 source.n446 source.n445 9.3005
R865 source.n531 source.n530 9.3005
R866 source.n533 source.n532 9.3005
R867 source.n442 source.n441 9.3005
R868 source.n540 source.n539 9.3005
R869 source.n542 source.n541 9.3005
R870 source.n565 source.n564 9.3005
R871 source.n288 source.n287 9.3005
R872 source.n417 source.n416 9.3005
R873 source.n415 source.n414 9.3005
R874 source.n292 source.n291 9.3005
R875 source.n409 source.n408 9.3005
R876 source.n407 source.n406 9.3005
R877 source.n296 source.n295 9.3005
R878 source.n375 source.n374 9.3005
R879 source.n373 source.n372 9.3005
R880 source.n312 source.n311 9.3005
R881 source.n367 source.n366 9.3005
R882 source.n365 source.n364 9.3005
R883 source.n316 source.n315 9.3005
R884 source.n359 source.n358 9.3005
R885 source.n357 source.n356 9.3005
R886 source.n333 source.n332 9.3005
R887 source.n328 source.n327 9.3005
R888 source.n339 source.n338 9.3005
R889 source.n341 source.n340 9.3005
R890 source.n324 source.n323 9.3005
R891 source.n347 source.n346 9.3005
R892 source.n349 source.n348 9.3005
R893 source.n350 source.n319 9.3005
R894 source.n308 source.n307 9.3005
R895 source.n381 source.n380 9.3005
R896 source.n383 source.n382 9.3005
R897 source.n304 source.n303 9.3005
R898 source.n389 source.n388 9.3005
R899 source.n391 source.n390 9.3005
R900 source.n300 source.n299 9.3005
R901 source.n398 source.n397 9.3005
R902 source.n400 source.n399 9.3005
R903 source.n423 source.n422 9.3005
R904 source.n49 source.n48 9.3005
R905 source.n44 source.n43 9.3005
R906 source.n55 source.n54 9.3005
R907 source.n57 source.n56 9.3005
R908 source.n40 source.n39 9.3005
R909 source.n63 source.n62 9.3005
R910 source.n65 source.n64 9.3005
R911 source.n37 source.n34 9.3005
R912 source.n96 source.n95 9.3005
R913 source.n98 source.n97 9.3005
R914 source.n19 source.n18 9.3005
R915 source.n104 source.n103 9.3005
R916 source.n106 source.n105 9.3005
R917 source.n14 source.n13 9.3005
R918 source.n112 source.n111 9.3005
R919 source.n114 source.n113 9.3005
R920 source.n137 source.n136 9.3005
R921 source.n2 source.n1 9.3005
R922 source.n131 source.n130 9.3005
R923 source.n129 source.n128 9.3005
R924 source.n6 source.n5 9.3005
R925 source.n123 source.n122 9.3005
R926 source.n121 source.n120 9.3005
R927 source.n10 source.n9 9.3005
R928 source.n23 source.n22 9.3005
R929 source.n90 source.n89 9.3005
R930 source.n88 source.n87 9.3005
R931 source.n27 source.n26 9.3005
R932 source.n82 source.n81 9.3005
R933 source.n80 source.n79 9.3005
R934 source.n31 source.n30 9.3005
R935 source.n74 source.n73 9.3005
R936 source.n72 source.n71 9.3005
R937 source.n191 source.n190 9.3005
R938 source.n186 source.n185 9.3005
R939 source.n197 source.n196 9.3005
R940 source.n199 source.n198 9.3005
R941 source.n182 source.n181 9.3005
R942 source.n205 source.n204 9.3005
R943 source.n207 source.n206 9.3005
R944 source.n179 source.n176 9.3005
R945 source.n238 source.n237 9.3005
R946 source.n240 source.n239 9.3005
R947 source.n161 source.n160 9.3005
R948 source.n246 source.n245 9.3005
R949 source.n248 source.n247 9.3005
R950 source.n156 source.n155 9.3005
R951 source.n254 source.n253 9.3005
R952 source.n256 source.n255 9.3005
R953 source.n279 source.n278 9.3005
R954 source.n144 source.n143 9.3005
R955 source.n273 source.n272 9.3005
R956 source.n271 source.n270 9.3005
R957 source.n148 source.n147 9.3005
R958 source.n265 source.n264 9.3005
R959 source.n263 source.n262 9.3005
R960 source.n152 source.n151 9.3005
R961 source.n165 source.n164 9.3005
R962 source.n232 source.n231 9.3005
R963 source.n230 source.n229 9.3005
R964 source.n169 source.n168 9.3005
R965 source.n224 source.n223 9.3005
R966 source.n222 source.n221 9.3005
R967 source.n173 source.n172 9.3005
R968 source.n216 source.n215 9.3005
R969 source.n214 source.n213 9.3005
R970 source.n480 source.n479 8.92171
R971 source.n513 source.n454 8.92171
R972 source.n526 source.n446 8.92171
R973 source.n560 source.n559 8.92171
R974 source.n338 source.n337 8.92171
R975 source.n371 source.n312 8.92171
R976 source.n384 source.n304 8.92171
R977 source.n418 source.n417 8.92171
R978 source.n132 source.n131 8.92171
R979 source.n99 source.n19 8.92171
R980 source.n86 source.n27 8.92171
R981 source.n54 source.n53 8.92171
R982 source.n274 source.n273 8.92171
R983 source.n241 source.n161 8.92171
R984 source.n228 source.n169 8.92171
R985 source.n196 source.n195 8.92171
R986 source.n476 source.n470 8.14595
R987 source.n514 source.n452 8.14595
R988 source.n525 source.n448 8.14595
R989 source.n563 source.n430 8.14595
R990 source.n334 source.n328 8.14595
R991 source.n372 source.n310 8.14595
R992 source.n383 source.n306 8.14595
R993 source.n421 source.n288 8.14595
R994 source.n135 source.n2 8.14595
R995 source.n98 source.n21 8.14595
R996 source.n87 source.n25 8.14595
R997 source.n50 source.n44 8.14595
R998 source.n277 source.n144 8.14595
R999 source.n240 source.n163 8.14595
R1000 source.n229 source.n167 8.14595
R1001 source.n192 source.n186 8.14595
R1002 source.n475 source.n472 7.3702
R1003 source.n518 source.n517 7.3702
R1004 source.n522 source.n521 7.3702
R1005 source.n564 source.n428 7.3702
R1006 source.n333 source.n330 7.3702
R1007 source.n376 source.n375 7.3702
R1008 source.n380 source.n379 7.3702
R1009 source.n422 source.n286 7.3702
R1010 source.n136 source.n0 7.3702
R1011 source.n95 source.n94 7.3702
R1012 source.n91 source.n90 7.3702
R1013 source.n49 source.n46 7.3702
R1014 source.n278 source.n142 7.3702
R1015 source.n237 source.n236 7.3702
R1016 source.n233 source.n232 7.3702
R1017 source.n191 source.n188 7.3702
R1018 source.n518 source.n450 6.59444
R1019 source.n521 source.n450 6.59444
R1020 source.n566 source.n428 6.59444
R1021 source.n376 source.n308 6.59444
R1022 source.n379 source.n308 6.59444
R1023 source.n424 source.n286 6.59444
R1024 source.n138 source.n0 6.59444
R1025 source.n94 source.n23 6.59444
R1026 source.n91 source.n23 6.59444
R1027 source.n280 source.n142 6.59444
R1028 source.n236 source.n165 6.59444
R1029 source.n233 source.n165 6.59444
R1030 source.n476 source.n475 5.81868
R1031 source.n517 source.n452 5.81868
R1032 source.n522 source.n448 5.81868
R1033 source.n564 source.n563 5.81868
R1034 source.n334 source.n333 5.81868
R1035 source.n375 source.n310 5.81868
R1036 source.n380 source.n306 5.81868
R1037 source.n422 source.n421 5.81868
R1038 source.n136 source.n135 5.81868
R1039 source.n95 source.n21 5.81868
R1040 source.n90 source.n25 5.81868
R1041 source.n50 source.n49 5.81868
R1042 source.n278 source.n277 5.81868
R1043 source.n237 source.n163 5.81868
R1044 source.n232 source.n167 5.81868
R1045 source.n192 source.n191 5.81868
R1046 source.n568 source.n567 5.51343
R1047 source.n479 source.n470 5.04292
R1048 source.n514 source.n513 5.04292
R1049 source.n526 source.n525 5.04292
R1050 source.n560 source.n430 5.04292
R1051 source.n337 source.n328 5.04292
R1052 source.n372 source.n371 5.04292
R1053 source.n384 source.n383 5.04292
R1054 source.n418 source.n288 5.04292
R1055 source.n132 source.n2 5.04292
R1056 source.n99 source.n98 5.04292
R1057 source.n87 source.n86 5.04292
R1058 source.n53 source.n44 5.04292
R1059 source.n274 source.n144 5.04292
R1060 source.n241 source.n240 5.04292
R1061 source.n229 source.n228 5.04292
R1062 source.n195 source.n186 5.04292
R1063 source.n480 source.n468 4.26717
R1064 source.n510 source.n454 4.26717
R1065 source.n529 source.n446 4.26717
R1066 source.n559 source.n432 4.26717
R1067 source.n338 source.n326 4.26717
R1068 source.n368 source.n312 4.26717
R1069 source.n387 source.n304 4.26717
R1070 source.n417 source.n290 4.26717
R1071 source.n131 source.n4 4.26717
R1072 source.n102 source.n19 4.26717
R1073 source.n83 source.n27 4.26717
R1074 source.n54 source.n42 4.26717
R1075 source.n273 source.n146 4.26717
R1076 source.n244 source.n161 4.26717
R1077 source.n225 source.n169 4.26717
R1078 source.n196 source.n184 4.26717
R1079 source.n484 source.n483 3.49141
R1080 source.n509 source.n456 3.49141
R1081 source.n530 source.n444 3.49141
R1082 source.n556 source.n555 3.49141
R1083 source.n342 source.n341 3.49141
R1084 source.n367 source.n314 3.49141
R1085 source.n388 source.n302 3.49141
R1086 source.n414 source.n413 3.49141
R1087 source.n128 source.n127 3.49141
R1088 source.n103 source.n17 3.49141
R1089 source.n82 source.n29 3.49141
R1090 source.n58 source.n57 3.49141
R1091 source.n270 source.n269 3.49141
R1092 source.n245 source.n159 3.49141
R1093 source.n224 source.n171 3.49141
R1094 source.n200 source.n199 3.49141
R1095 source.n48 source.n47 2.84303
R1096 source.n190 source.n189 2.84303
R1097 source.n474 source.n473 2.84303
R1098 source.n332 source.n331 2.84303
R1099 source.n487 source.n466 2.71565
R1100 source.n506 source.n505 2.71565
R1101 source.n534 source.n533 2.71565
R1102 source.n552 source.n434 2.71565
R1103 source.n345 source.n324 2.71565
R1104 source.n364 source.n363 2.71565
R1105 source.n392 source.n391 2.71565
R1106 source.n410 source.n292 2.71565
R1107 source.n124 source.n6 2.71565
R1108 source.n107 source.n106 2.71565
R1109 source.n79 source.n78 2.71565
R1110 source.n61 source.n40 2.71565
R1111 source.n266 source.n148 2.71565
R1112 source.n249 source.n248 2.71565
R1113 source.n221 source.n220 2.71565
R1114 source.n203 source.n182 2.71565
R1115 source.n488 source.n464 1.93989
R1116 source.n502 source.n458 1.93989
R1117 source.n538 source.n442 1.93989
R1118 source.n551 source.n436 1.93989
R1119 source.n346 source.n322 1.93989
R1120 source.n360 source.n316 1.93989
R1121 source.n396 source.n300 1.93989
R1122 source.n409 source.n294 1.93989
R1123 source.n123 source.n8 1.93989
R1124 source.n110 source.n14 1.93989
R1125 source.n75 source.n31 1.93989
R1126 source.n62 source.n38 1.93989
R1127 source.n265 source.n150 1.93989
R1128 source.n252 source.n156 1.93989
R1129 source.n217 source.n173 1.93989
R1130 source.n204 source.n180 1.93989
R1131 source.n493 source.n491 1.16414
R1132 source.n501 source.n460 1.16414
R1133 source.n539 source.n440 1.16414
R1134 source.n548 source.n547 1.16414
R1135 source.n351 source.n349 1.16414
R1136 source.n359 source.n318 1.16414
R1137 source.n397 source.n298 1.16414
R1138 source.n406 source.n405 1.16414
R1139 source.n120 source.n119 1.16414
R1140 source.n111 source.n12 1.16414
R1141 source.n74 source.n33 1.16414
R1142 source.n66 source.n65 1.16414
R1143 source.n262 source.n261 1.16414
R1144 source.n253 source.n154 1.16414
R1145 source.n216 source.n175 1.16414
R1146 source.n208 source.n207 1.16414
R1147 source.n426 source.t2 0.7925
R1148 source.n426 source.t1 0.7925
R1149 source.n284 source.t8 0.7925
R1150 source.n284 source.t7 0.7925
R1151 source.n140 source.t10 0.7925
R1152 source.n140 source.t11 0.7925
R1153 source.n282 source.t0 0.7925
R1154 source.n282 source.t3 0.7925
R1155 source.n281 source.n141 0.720328
R1156 source.n427 source.n425 0.720328
R1157 source.n283 source.n281 0.5005
R1158 source.n141 source.n139 0.5005
R1159 source.n425 source.n285 0.5005
R1160 source.n567 source.n427 0.5005
R1161 source.n492 source.n462 0.388379
R1162 source.n498 source.n497 0.388379
R1163 source.n543 source.n542 0.388379
R1164 source.n544 source.n438 0.388379
R1165 source.n350 source.n320 0.388379
R1166 source.n356 source.n355 0.388379
R1167 source.n401 source.n400 0.388379
R1168 source.n402 source.n296 0.388379
R1169 source.n116 source.n10 0.388379
R1170 source.n115 source.n114 0.388379
R1171 source.n71 source.n70 0.388379
R1172 source.n37 source.n35 0.388379
R1173 source.n258 source.n152 0.388379
R1174 source.n257 source.n256 0.388379
R1175 source.n213 source.n212 0.388379
R1176 source.n179 source.n177 0.388379
R1177 source source.n568 0.188
R1178 source.n474 source.n469 0.155672
R1179 source.n481 source.n469 0.155672
R1180 source.n482 source.n481 0.155672
R1181 source.n482 source.n465 0.155672
R1182 source.n489 source.n465 0.155672
R1183 source.n490 source.n489 0.155672
R1184 source.n490 source.n461 0.155672
R1185 source.n499 source.n461 0.155672
R1186 source.n500 source.n499 0.155672
R1187 source.n500 source.n457 0.155672
R1188 source.n507 source.n457 0.155672
R1189 source.n508 source.n507 0.155672
R1190 source.n508 source.n453 0.155672
R1191 source.n515 source.n453 0.155672
R1192 source.n516 source.n515 0.155672
R1193 source.n516 source.n449 0.155672
R1194 source.n523 source.n449 0.155672
R1195 source.n524 source.n523 0.155672
R1196 source.n524 source.n445 0.155672
R1197 source.n531 source.n445 0.155672
R1198 source.n532 source.n531 0.155672
R1199 source.n532 source.n441 0.155672
R1200 source.n540 source.n441 0.155672
R1201 source.n541 source.n540 0.155672
R1202 source.n541 source.n437 0.155672
R1203 source.n549 source.n437 0.155672
R1204 source.n550 source.n549 0.155672
R1205 source.n550 source.n433 0.155672
R1206 source.n557 source.n433 0.155672
R1207 source.n558 source.n557 0.155672
R1208 source.n558 source.n429 0.155672
R1209 source.n565 source.n429 0.155672
R1210 source.n332 source.n327 0.155672
R1211 source.n339 source.n327 0.155672
R1212 source.n340 source.n339 0.155672
R1213 source.n340 source.n323 0.155672
R1214 source.n347 source.n323 0.155672
R1215 source.n348 source.n347 0.155672
R1216 source.n348 source.n319 0.155672
R1217 source.n357 source.n319 0.155672
R1218 source.n358 source.n357 0.155672
R1219 source.n358 source.n315 0.155672
R1220 source.n365 source.n315 0.155672
R1221 source.n366 source.n365 0.155672
R1222 source.n366 source.n311 0.155672
R1223 source.n373 source.n311 0.155672
R1224 source.n374 source.n373 0.155672
R1225 source.n374 source.n307 0.155672
R1226 source.n381 source.n307 0.155672
R1227 source.n382 source.n381 0.155672
R1228 source.n382 source.n303 0.155672
R1229 source.n389 source.n303 0.155672
R1230 source.n390 source.n389 0.155672
R1231 source.n390 source.n299 0.155672
R1232 source.n398 source.n299 0.155672
R1233 source.n399 source.n398 0.155672
R1234 source.n399 source.n295 0.155672
R1235 source.n407 source.n295 0.155672
R1236 source.n408 source.n407 0.155672
R1237 source.n408 source.n291 0.155672
R1238 source.n415 source.n291 0.155672
R1239 source.n416 source.n415 0.155672
R1240 source.n416 source.n287 0.155672
R1241 source.n423 source.n287 0.155672
R1242 source.n137 source.n1 0.155672
R1243 source.n130 source.n1 0.155672
R1244 source.n130 source.n129 0.155672
R1245 source.n129 source.n5 0.155672
R1246 source.n122 source.n5 0.155672
R1247 source.n122 source.n121 0.155672
R1248 source.n121 source.n9 0.155672
R1249 source.n113 source.n9 0.155672
R1250 source.n113 source.n112 0.155672
R1251 source.n112 source.n13 0.155672
R1252 source.n105 source.n13 0.155672
R1253 source.n105 source.n104 0.155672
R1254 source.n104 source.n18 0.155672
R1255 source.n97 source.n18 0.155672
R1256 source.n97 source.n96 0.155672
R1257 source.n96 source.n22 0.155672
R1258 source.n89 source.n22 0.155672
R1259 source.n89 source.n88 0.155672
R1260 source.n88 source.n26 0.155672
R1261 source.n81 source.n26 0.155672
R1262 source.n81 source.n80 0.155672
R1263 source.n80 source.n30 0.155672
R1264 source.n73 source.n30 0.155672
R1265 source.n73 source.n72 0.155672
R1266 source.n72 source.n34 0.155672
R1267 source.n64 source.n34 0.155672
R1268 source.n64 source.n63 0.155672
R1269 source.n63 source.n39 0.155672
R1270 source.n56 source.n39 0.155672
R1271 source.n56 source.n55 0.155672
R1272 source.n55 source.n43 0.155672
R1273 source.n48 source.n43 0.155672
R1274 source.n279 source.n143 0.155672
R1275 source.n272 source.n143 0.155672
R1276 source.n272 source.n271 0.155672
R1277 source.n271 source.n147 0.155672
R1278 source.n264 source.n147 0.155672
R1279 source.n264 source.n263 0.155672
R1280 source.n263 source.n151 0.155672
R1281 source.n255 source.n151 0.155672
R1282 source.n255 source.n254 0.155672
R1283 source.n254 source.n155 0.155672
R1284 source.n247 source.n155 0.155672
R1285 source.n247 source.n246 0.155672
R1286 source.n246 source.n160 0.155672
R1287 source.n239 source.n160 0.155672
R1288 source.n239 source.n238 0.155672
R1289 source.n238 source.n164 0.155672
R1290 source.n231 source.n164 0.155672
R1291 source.n231 source.n230 0.155672
R1292 source.n230 source.n168 0.155672
R1293 source.n223 source.n168 0.155672
R1294 source.n223 source.n222 0.155672
R1295 source.n222 source.n172 0.155672
R1296 source.n215 source.n172 0.155672
R1297 source.n215 source.n214 0.155672
R1298 source.n214 source.n176 0.155672
R1299 source.n206 source.n176 0.155672
R1300 source.n206 source.n205 0.155672
R1301 source.n205 source.n181 0.155672
R1302 source.n198 source.n181 0.155672
R1303 source.n198 source.n197 0.155672
R1304 source.n197 source.n185 0.155672
R1305 source.n190 source.n185 0.155672
R1306 minus.n2 minus.t3 2583.52
R1307 minus.n0 minus.t4 2583.52
R1308 minus.n6 minus.t5 2583.52
R1309 minus.n4 minus.t0 2583.52
R1310 minus.n1 minus.t1 2535.32
R1311 minus.n5 minus.t2 2535.32
R1312 minus.n3 minus.n0 161.489
R1313 minus.n7 minus.n4 161.489
R1314 minus.n3 minus.n2 161.3
R1315 minus.n7 minus.n6 161.3
R1316 minus.n8 minus.n3 43.4247
R1317 minus.n2 minus.n1 36.5157
R1318 minus.n1 minus.n0 36.5157
R1319 minus.n5 minus.n4 36.5157
R1320 minus.n6 minus.n5 36.5157
R1321 minus.n8 minus.n7 6.48535
R1322 minus minus.n8 0.188
R1323 drain_right.n134 drain_right.n0 289.615
R1324 drain_right.n276 drain_right.n142 289.615
R1325 drain_right.n44 drain_right.n43 185
R1326 drain_right.n49 drain_right.n48 185
R1327 drain_right.n51 drain_right.n50 185
R1328 drain_right.n40 drain_right.n39 185
R1329 drain_right.n57 drain_right.n56 185
R1330 drain_right.n59 drain_right.n58 185
R1331 drain_right.n36 drain_right.n35 185
R1332 drain_right.n66 drain_right.n65 185
R1333 drain_right.n67 drain_right.n34 185
R1334 drain_right.n69 drain_right.n68 185
R1335 drain_right.n32 drain_right.n31 185
R1336 drain_right.n75 drain_right.n74 185
R1337 drain_right.n77 drain_right.n76 185
R1338 drain_right.n28 drain_right.n27 185
R1339 drain_right.n83 drain_right.n82 185
R1340 drain_right.n85 drain_right.n84 185
R1341 drain_right.n24 drain_right.n23 185
R1342 drain_right.n91 drain_right.n90 185
R1343 drain_right.n93 drain_right.n92 185
R1344 drain_right.n20 drain_right.n19 185
R1345 drain_right.n99 drain_right.n98 185
R1346 drain_right.n101 drain_right.n100 185
R1347 drain_right.n16 drain_right.n15 185
R1348 drain_right.n107 drain_right.n106 185
R1349 drain_right.n110 drain_right.n109 185
R1350 drain_right.n108 drain_right.n12 185
R1351 drain_right.n115 drain_right.n11 185
R1352 drain_right.n117 drain_right.n116 185
R1353 drain_right.n119 drain_right.n118 185
R1354 drain_right.n8 drain_right.n7 185
R1355 drain_right.n125 drain_right.n124 185
R1356 drain_right.n127 drain_right.n126 185
R1357 drain_right.n4 drain_right.n3 185
R1358 drain_right.n133 drain_right.n132 185
R1359 drain_right.n135 drain_right.n134 185
R1360 drain_right.n277 drain_right.n276 185
R1361 drain_right.n275 drain_right.n274 185
R1362 drain_right.n146 drain_right.n145 185
R1363 drain_right.n269 drain_right.n268 185
R1364 drain_right.n267 drain_right.n266 185
R1365 drain_right.n150 drain_right.n149 185
R1366 drain_right.n261 drain_right.n260 185
R1367 drain_right.n259 drain_right.n258 185
R1368 drain_right.n257 drain_right.n153 185
R1369 drain_right.n157 drain_right.n154 185
R1370 drain_right.n252 drain_right.n251 185
R1371 drain_right.n250 drain_right.n249 185
R1372 drain_right.n159 drain_right.n158 185
R1373 drain_right.n244 drain_right.n243 185
R1374 drain_right.n242 drain_right.n241 185
R1375 drain_right.n163 drain_right.n162 185
R1376 drain_right.n236 drain_right.n235 185
R1377 drain_right.n234 drain_right.n233 185
R1378 drain_right.n167 drain_right.n166 185
R1379 drain_right.n228 drain_right.n227 185
R1380 drain_right.n226 drain_right.n225 185
R1381 drain_right.n171 drain_right.n170 185
R1382 drain_right.n220 drain_right.n219 185
R1383 drain_right.n218 drain_right.n217 185
R1384 drain_right.n175 drain_right.n174 185
R1385 drain_right.n212 drain_right.n211 185
R1386 drain_right.n210 drain_right.n177 185
R1387 drain_right.n209 drain_right.n208 185
R1388 drain_right.n180 drain_right.n178 185
R1389 drain_right.n203 drain_right.n202 185
R1390 drain_right.n201 drain_right.n200 185
R1391 drain_right.n184 drain_right.n183 185
R1392 drain_right.n195 drain_right.n194 185
R1393 drain_right.n193 drain_right.n192 185
R1394 drain_right.n188 drain_right.n187 185
R1395 drain_right.n45 drain_right.t5 149.524
R1396 drain_right.n189 drain_right.t2 149.524
R1397 drain_right.n49 drain_right.n43 104.615
R1398 drain_right.n50 drain_right.n49 104.615
R1399 drain_right.n50 drain_right.n39 104.615
R1400 drain_right.n57 drain_right.n39 104.615
R1401 drain_right.n58 drain_right.n57 104.615
R1402 drain_right.n58 drain_right.n35 104.615
R1403 drain_right.n66 drain_right.n35 104.615
R1404 drain_right.n67 drain_right.n66 104.615
R1405 drain_right.n68 drain_right.n67 104.615
R1406 drain_right.n68 drain_right.n31 104.615
R1407 drain_right.n75 drain_right.n31 104.615
R1408 drain_right.n76 drain_right.n75 104.615
R1409 drain_right.n76 drain_right.n27 104.615
R1410 drain_right.n83 drain_right.n27 104.615
R1411 drain_right.n84 drain_right.n83 104.615
R1412 drain_right.n84 drain_right.n23 104.615
R1413 drain_right.n91 drain_right.n23 104.615
R1414 drain_right.n92 drain_right.n91 104.615
R1415 drain_right.n92 drain_right.n19 104.615
R1416 drain_right.n99 drain_right.n19 104.615
R1417 drain_right.n100 drain_right.n99 104.615
R1418 drain_right.n100 drain_right.n15 104.615
R1419 drain_right.n107 drain_right.n15 104.615
R1420 drain_right.n109 drain_right.n107 104.615
R1421 drain_right.n109 drain_right.n108 104.615
R1422 drain_right.n108 drain_right.n11 104.615
R1423 drain_right.n117 drain_right.n11 104.615
R1424 drain_right.n118 drain_right.n117 104.615
R1425 drain_right.n118 drain_right.n7 104.615
R1426 drain_right.n125 drain_right.n7 104.615
R1427 drain_right.n126 drain_right.n125 104.615
R1428 drain_right.n126 drain_right.n3 104.615
R1429 drain_right.n133 drain_right.n3 104.615
R1430 drain_right.n134 drain_right.n133 104.615
R1431 drain_right.n276 drain_right.n275 104.615
R1432 drain_right.n275 drain_right.n145 104.615
R1433 drain_right.n268 drain_right.n145 104.615
R1434 drain_right.n268 drain_right.n267 104.615
R1435 drain_right.n267 drain_right.n149 104.615
R1436 drain_right.n260 drain_right.n149 104.615
R1437 drain_right.n260 drain_right.n259 104.615
R1438 drain_right.n259 drain_right.n153 104.615
R1439 drain_right.n157 drain_right.n153 104.615
R1440 drain_right.n251 drain_right.n157 104.615
R1441 drain_right.n251 drain_right.n250 104.615
R1442 drain_right.n250 drain_right.n158 104.615
R1443 drain_right.n243 drain_right.n158 104.615
R1444 drain_right.n243 drain_right.n242 104.615
R1445 drain_right.n242 drain_right.n162 104.615
R1446 drain_right.n235 drain_right.n162 104.615
R1447 drain_right.n235 drain_right.n234 104.615
R1448 drain_right.n234 drain_right.n166 104.615
R1449 drain_right.n227 drain_right.n166 104.615
R1450 drain_right.n227 drain_right.n226 104.615
R1451 drain_right.n226 drain_right.n170 104.615
R1452 drain_right.n219 drain_right.n170 104.615
R1453 drain_right.n219 drain_right.n218 104.615
R1454 drain_right.n218 drain_right.n174 104.615
R1455 drain_right.n211 drain_right.n174 104.615
R1456 drain_right.n211 drain_right.n210 104.615
R1457 drain_right.n210 drain_right.n209 104.615
R1458 drain_right.n209 drain_right.n178 104.615
R1459 drain_right.n202 drain_right.n178 104.615
R1460 drain_right.n202 drain_right.n201 104.615
R1461 drain_right.n201 drain_right.n183 104.615
R1462 drain_right.n194 drain_right.n183 104.615
R1463 drain_right.n194 drain_right.n193 104.615
R1464 drain_right.n193 drain_right.n187 104.615
R1465 drain_right.n281 drain_right.n141 59.2153
R1466 drain_right.n140 drain_right.n139 58.7851
R1467 drain_right.t5 drain_right.n43 52.3082
R1468 drain_right.t2 drain_right.n187 52.3082
R1469 drain_right.n140 drain_right.n138 47.6323
R1470 drain_right.n281 drain_right.n280 47.3126
R1471 drain_right drain_right.n140 38.0373
R1472 drain_right.n69 drain_right.n34 13.1884
R1473 drain_right.n116 drain_right.n115 13.1884
R1474 drain_right.n258 drain_right.n257 13.1884
R1475 drain_right.n212 drain_right.n177 13.1884
R1476 drain_right.n65 drain_right.n64 12.8005
R1477 drain_right.n70 drain_right.n32 12.8005
R1478 drain_right.n114 drain_right.n12 12.8005
R1479 drain_right.n119 drain_right.n10 12.8005
R1480 drain_right.n261 drain_right.n152 12.8005
R1481 drain_right.n256 drain_right.n154 12.8005
R1482 drain_right.n213 drain_right.n175 12.8005
R1483 drain_right.n208 drain_right.n179 12.8005
R1484 drain_right.n63 drain_right.n36 12.0247
R1485 drain_right.n74 drain_right.n73 12.0247
R1486 drain_right.n111 drain_right.n110 12.0247
R1487 drain_right.n120 drain_right.n8 12.0247
R1488 drain_right.n262 drain_right.n150 12.0247
R1489 drain_right.n253 drain_right.n252 12.0247
R1490 drain_right.n217 drain_right.n216 12.0247
R1491 drain_right.n207 drain_right.n180 12.0247
R1492 drain_right.n60 drain_right.n59 11.249
R1493 drain_right.n77 drain_right.n30 11.249
R1494 drain_right.n106 drain_right.n14 11.249
R1495 drain_right.n124 drain_right.n123 11.249
R1496 drain_right.n266 drain_right.n265 11.249
R1497 drain_right.n249 drain_right.n156 11.249
R1498 drain_right.n220 drain_right.n173 11.249
R1499 drain_right.n204 drain_right.n203 11.249
R1500 drain_right.n56 drain_right.n38 10.4732
R1501 drain_right.n78 drain_right.n28 10.4732
R1502 drain_right.n105 drain_right.n16 10.4732
R1503 drain_right.n127 drain_right.n6 10.4732
R1504 drain_right.n269 drain_right.n148 10.4732
R1505 drain_right.n248 drain_right.n159 10.4732
R1506 drain_right.n221 drain_right.n171 10.4732
R1507 drain_right.n200 drain_right.n182 10.4732
R1508 drain_right.n45 drain_right.n44 10.2747
R1509 drain_right.n189 drain_right.n188 10.2747
R1510 drain_right.n55 drain_right.n40 9.69747
R1511 drain_right.n82 drain_right.n81 9.69747
R1512 drain_right.n102 drain_right.n101 9.69747
R1513 drain_right.n128 drain_right.n4 9.69747
R1514 drain_right.n270 drain_right.n146 9.69747
R1515 drain_right.n245 drain_right.n244 9.69747
R1516 drain_right.n225 drain_right.n224 9.69747
R1517 drain_right.n199 drain_right.n184 9.69747
R1518 drain_right.n138 drain_right.n137 9.45567
R1519 drain_right.n280 drain_right.n279 9.45567
R1520 drain_right.n2 drain_right.n1 9.3005
R1521 drain_right.n131 drain_right.n130 9.3005
R1522 drain_right.n129 drain_right.n128 9.3005
R1523 drain_right.n6 drain_right.n5 9.3005
R1524 drain_right.n123 drain_right.n122 9.3005
R1525 drain_right.n121 drain_right.n120 9.3005
R1526 drain_right.n10 drain_right.n9 9.3005
R1527 drain_right.n89 drain_right.n88 9.3005
R1528 drain_right.n87 drain_right.n86 9.3005
R1529 drain_right.n26 drain_right.n25 9.3005
R1530 drain_right.n81 drain_right.n80 9.3005
R1531 drain_right.n79 drain_right.n78 9.3005
R1532 drain_right.n30 drain_right.n29 9.3005
R1533 drain_right.n73 drain_right.n72 9.3005
R1534 drain_right.n71 drain_right.n70 9.3005
R1535 drain_right.n47 drain_right.n46 9.3005
R1536 drain_right.n42 drain_right.n41 9.3005
R1537 drain_right.n53 drain_right.n52 9.3005
R1538 drain_right.n55 drain_right.n54 9.3005
R1539 drain_right.n38 drain_right.n37 9.3005
R1540 drain_right.n61 drain_right.n60 9.3005
R1541 drain_right.n63 drain_right.n62 9.3005
R1542 drain_right.n64 drain_right.n33 9.3005
R1543 drain_right.n22 drain_right.n21 9.3005
R1544 drain_right.n95 drain_right.n94 9.3005
R1545 drain_right.n97 drain_right.n96 9.3005
R1546 drain_right.n18 drain_right.n17 9.3005
R1547 drain_right.n103 drain_right.n102 9.3005
R1548 drain_right.n105 drain_right.n104 9.3005
R1549 drain_right.n14 drain_right.n13 9.3005
R1550 drain_right.n112 drain_right.n111 9.3005
R1551 drain_right.n114 drain_right.n113 9.3005
R1552 drain_right.n137 drain_right.n136 9.3005
R1553 drain_right.n191 drain_right.n190 9.3005
R1554 drain_right.n186 drain_right.n185 9.3005
R1555 drain_right.n197 drain_right.n196 9.3005
R1556 drain_right.n199 drain_right.n198 9.3005
R1557 drain_right.n182 drain_right.n181 9.3005
R1558 drain_right.n205 drain_right.n204 9.3005
R1559 drain_right.n207 drain_right.n206 9.3005
R1560 drain_right.n179 drain_right.n176 9.3005
R1561 drain_right.n238 drain_right.n237 9.3005
R1562 drain_right.n240 drain_right.n239 9.3005
R1563 drain_right.n161 drain_right.n160 9.3005
R1564 drain_right.n246 drain_right.n245 9.3005
R1565 drain_right.n248 drain_right.n247 9.3005
R1566 drain_right.n156 drain_right.n155 9.3005
R1567 drain_right.n254 drain_right.n253 9.3005
R1568 drain_right.n256 drain_right.n255 9.3005
R1569 drain_right.n279 drain_right.n278 9.3005
R1570 drain_right.n144 drain_right.n143 9.3005
R1571 drain_right.n273 drain_right.n272 9.3005
R1572 drain_right.n271 drain_right.n270 9.3005
R1573 drain_right.n148 drain_right.n147 9.3005
R1574 drain_right.n265 drain_right.n264 9.3005
R1575 drain_right.n263 drain_right.n262 9.3005
R1576 drain_right.n152 drain_right.n151 9.3005
R1577 drain_right.n165 drain_right.n164 9.3005
R1578 drain_right.n232 drain_right.n231 9.3005
R1579 drain_right.n230 drain_right.n229 9.3005
R1580 drain_right.n169 drain_right.n168 9.3005
R1581 drain_right.n224 drain_right.n223 9.3005
R1582 drain_right.n222 drain_right.n221 9.3005
R1583 drain_right.n173 drain_right.n172 9.3005
R1584 drain_right.n216 drain_right.n215 9.3005
R1585 drain_right.n214 drain_right.n213 9.3005
R1586 drain_right.n52 drain_right.n51 8.92171
R1587 drain_right.n85 drain_right.n26 8.92171
R1588 drain_right.n98 drain_right.n18 8.92171
R1589 drain_right.n132 drain_right.n131 8.92171
R1590 drain_right.n274 drain_right.n273 8.92171
R1591 drain_right.n241 drain_right.n161 8.92171
R1592 drain_right.n228 drain_right.n169 8.92171
R1593 drain_right.n196 drain_right.n195 8.92171
R1594 drain_right.n48 drain_right.n42 8.14595
R1595 drain_right.n86 drain_right.n24 8.14595
R1596 drain_right.n97 drain_right.n20 8.14595
R1597 drain_right.n135 drain_right.n2 8.14595
R1598 drain_right.n277 drain_right.n144 8.14595
R1599 drain_right.n240 drain_right.n163 8.14595
R1600 drain_right.n229 drain_right.n167 8.14595
R1601 drain_right.n192 drain_right.n186 8.14595
R1602 drain_right.n47 drain_right.n44 7.3702
R1603 drain_right.n90 drain_right.n89 7.3702
R1604 drain_right.n94 drain_right.n93 7.3702
R1605 drain_right.n136 drain_right.n0 7.3702
R1606 drain_right.n278 drain_right.n142 7.3702
R1607 drain_right.n237 drain_right.n236 7.3702
R1608 drain_right.n233 drain_right.n232 7.3702
R1609 drain_right.n191 drain_right.n188 7.3702
R1610 drain_right.n90 drain_right.n22 6.59444
R1611 drain_right.n93 drain_right.n22 6.59444
R1612 drain_right.n138 drain_right.n0 6.59444
R1613 drain_right.n280 drain_right.n142 6.59444
R1614 drain_right.n236 drain_right.n165 6.59444
R1615 drain_right.n233 drain_right.n165 6.59444
R1616 drain_right drain_right.n281 5.90322
R1617 drain_right.n48 drain_right.n47 5.81868
R1618 drain_right.n89 drain_right.n24 5.81868
R1619 drain_right.n94 drain_right.n20 5.81868
R1620 drain_right.n136 drain_right.n135 5.81868
R1621 drain_right.n278 drain_right.n277 5.81868
R1622 drain_right.n237 drain_right.n163 5.81868
R1623 drain_right.n232 drain_right.n167 5.81868
R1624 drain_right.n192 drain_right.n191 5.81868
R1625 drain_right.n51 drain_right.n42 5.04292
R1626 drain_right.n86 drain_right.n85 5.04292
R1627 drain_right.n98 drain_right.n97 5.04292
R1628 drain_right.n132 drain_right.n2 5.04292
R1629 drain_right.n274 drain_right.n144 5.04292
R1630 drain_right.n241 drain_right.n240 5.04292
R1631 drain_right.n229 drain_right.n228 5.04292
R1632 drain_right.n195 drain_right.n186 5.04292
R1633 drain_right.n52 drain_right.n40 4.26717
R1634 drain_right.n82 drain_right.n26 4.26717
R1635 drain_right.n101 drain_right.n18 4.26717
R1636 drain_right.n131 drain_right.n4 4.26717
R1637 drain_right.n273 drain_right.n146 4.26717
R1638 drain_right.n244 drain_right.n161 4.26717
R1639 drain_right.n225 drain_right.n169 4.26717
R1640 drain_right.n196 drain_right.n184 4.26717
R1641 drain_right.n56 drain_right.n55 3.49141
R1642 drain_right.n81 drain_right.n28 3.49141
R1643 drain_right.n102 drain_right.n16 3.49141
R1644 drain_right.n128 drain_right.n127 3.49141
R1645 drain_right.n270 drain_right.n269 3.49141
R1646 drain_right.n245 drain_right.n159 3.49141
R1647 drain_right.n224 drain_right.n171 3.49141
R1648 drain_right.n200 drain_right.n199 3.49141
R1649 drain_right.n190 drain_right.n189 2.84303
R1650 drain_right.n46 drain_right.n45 2.84303
R1651 drain_right.n59 drain_right.n38 2.71565
R1652 drain_right.n78 drain_right.n77 2.71565
R1653 drain_right.n106 drain_right.n105 2.71565
R1654 drain_right.n124 drain_right.n6 2.71565
R1655 drain_right.n266 drain_right.n148 2.71565
R1656 drain_right.n249 drain_right.n248 2.71565
R1657 drain_right.n221 drain_right.n220 2.71565
R1658 drain_right.n203 drain_right.n182 2.71565
R1659 drain_right.n60 drain_right.n36 1.93989
R1660 drain_right.n74 drain_right.n30 1.93989
R1661 drain_right.n110 drain_right.n14 1.93989
R1662 drain_right.n123 drain_right.n8 1.93989
R1663 drain_right.n265 drain_right.n150 1.93989
R1664 drain_right.n252 drain_right.n156 1.93989
R1665 drain_right.n217 drain_right.n173 1.93989
R1666 drain_right.n204 drain_right.n180 1.93989
R1667 drain_right.n65 drain_right.n63 1.16414
R1668 drain_right.n73 drain_right.n32 1.16414
R1669 drain_right.n111 drain_right.n12 1.16414
R1670 drain_right.n120 drain_right.n119 1.16414
R1671 drain_right.n262 drain_right.n261 1.16414
R1672 drain_right.n253 drain_right.n154 1.16414
R1673 drain_right.n216 drain_right.n175 1.16414
R1674 drain_right.n208 drain_right.n207 1.16414
R1675 drain_right.n139 drain_right.t3 0.7925
R1676 drain_right.n139 drain_right.t0 0.7925
R1677 drain_right.n141 drain_right.t4 0.7925
R1678 drain_right.n141 drain_right.t1 0.7925
R1679 drain_right.n64 drain_right.n34 0.388379
R1680 drain_right.n70 drain_right.n69 0.388379
R1681 drain_right.n115 drain_right.n114 0.388379
R1682 drain_right.n116 drain_right.n10 0.388379
R1683 drain_right.n258 drain_right.n152 0.388379
R1684 drain_right.n257 drain_right.n256 0.388379
R1685 drain_right.n213 drain_right.n212 0.388379
R1686 drain_right.n179 drain_right.n177 0.388379
R1687 drain_right.n46 drain_right.n41 0.155672
R1688 drain_right.n53 drain_right.n41 0.155672
R1689 drain_right.n54 drain_right.n53 0.155672
R1690 drain_right.n54 drain_right.n37 0.155672
R1691 drain_right.n61 drain_right.n37 0.155672
R1692 drain_right.n62 drain_right.n61 0.155672
R1693 drain_right.n62 drain_right.n33 0.155672
R1694 drain_right.n71 drain_right.n33 0.155672
R1695 drain_right.n72 drain_right.n71 0.155672
R1696 drain_right.n72 drain_right.n29 0.155672
R1697 drain_right.n79 drain_right.n29 0.155672
R1698 drain_right.n80 drain_right.n79 0.155672
R1699 drain_right.n80 drain_right.n25 0.155672
R1700 drain_right.n87 drain_right.n25 0.155672
R1701 drain_right.n88 drain_right.n87 0.155672
R1702 drain_right.n88 drain_right.n21 0.155672
R1703 drain_right.n95 drain_right.n21 0.155672
R1704 drain_right.n96 drain_right.n95 0.155672
R1705 drain_right.n96 drain_right.n17 0.155672
R1706 drain_right.n103 drain_right.n17 0.155672
R1707 drain_right.n104 drain_right.n103 0.155672
R1708 drain_right.n104 drain_right.n13 0.155672
R1709 drain_right.n112 drain_right.n13 0.155672
R1710 drain_right.n113 drain_right.n112 0.155672
R1711 drain_right.n113 drain_right.n9 0.155672
R1712 drain_right.n121 drain_right.n9 0.155672
R1713 drain_right.n122 drain_right.n121 0.155672
R1714 drain_right.n122 drain_right.n5 0.155672
R1715 drain_right.n129 drain_right.n5 0.155672
R1716 drain_right.n130 drain_right.n129 0.155672
R1717 drain_right.n130 drain_right.n1 0.155672
R1718 drain_right.n137 drain_right.n1 0.155672
R1719 drain_right.n279 drain_right.n143 0.155672
R1720 drain_right.n272 drain_right.n143 0.155672
R1721 drain_right.n272 drain_right.n271 0.155672
R1722 drain_right.n271 drain_right.n147 0.155672
R1723 drain_right.n264 drain_right.n147 0.155672
R1724 drain_right.n264 drain_right.n263 0.155672
R1725 drain_right.n263 drain_right.n151 0.155672
R1726 drain_right.n255 drain_right.n151 0.155672
R1727 drain_right.n255 drain_right.n254 0.155672
R1728 drain_right.n254 drain_right.n155 0.155672
R1729 drain_right.n247 drain_right.n155 0.155672
R1730 drain_right.n247 drain_right.n246 0.155672
R1731 drain_right.n246 drain_right.n160 0.155672
R1732 drain_right.n239 drain_right.n160 0.155672
R1733 drain_right.n239 drain_right.n238 0.155672
R1734 drain_right.n238 drain_right.n164 0.155672
R1735 drain_right.n231 drain_right.n164 0.155672
R1736 drain_right.n231 drain_right.n230 0.155672
R1737 drain_right.n230 drain_right.n168 0.155672
R1738 drain_right.n223 drain_right.n168 0.155672
R1739 drain_right.n223 drain_right.n222 0.155672
R1740 drain_right.n222 drain_right.n172 0.155672
R1741 drain_right.n215 drain_right.n172 0.155672
R1742 drain_right.n215 drain_right.n214 0.155672
R1743 drain_right.n214 drain_right.n176 0.155672
R1744 drain_right.n206 drain_right.n176 0.155672
R1745 drain_right.n206 drain_right.n205 0.155672
R1746 drain_right.n205 drain_right.n181 0.155672
R1747 drain_right.n198 drain_right.n181 0.155672
R1748 drain_right.n198 drain_right.n197 0.155672
R1749 drain_right.n197 drain_right.n185 0.155672
R1750 drain_right.n190 drain_right.n185 0.155672
C0 minus drain_left 0.170597f
C1 plus drain_left 4.90024f
C2 source drain_left 29.721f
C3 minus drain_right 4.79626f
C4 plus drain_right 0.267908f
C5 source drain_right 29.697802f
C6 minus plus 7.02963f
C7 minus source 3.70961f
C8 plus source 3.72506f
C9 drain_left drain_right 0.557321f
C10 drain_right a_n1180_n5888# 10.241481f
C11 drain_left a_n1180_n5888# 10.425929f
C12 source a_n1180_n5888# 10.659655f
C13 minus a_n1180_n5888# 5.393314f
C14 plus a_n1180_n5888# 8.519679f
C15 drain_right.n0 a_n1180_n5888# 0.040373f
C16 drain_right.n1 a_n1180_n5888# 0.029285f
C17 drain_right.n2 a_n1180_n5888# 0.015737f
C18 drain_right.n3 a_n1180_n5888# 0.037196f
C19 drain_right.n4 a_n1180_n5888# 0.016662f
C20 drain_right.n5 a_n1180_n5888# 0.029285f
C21 drain_right.n6 a_n1180_n5888# 0.015737f
C22 drain_right.n7 a_n1180_n5888# 0.037196f
C23 drain_right.n8 a_n1180_n5888# 0.016662f
C24 drain_right.n9 a_n1180_n5888# 0.029285f
C25 drain_right.n10 a_n1180_n5888# 0.015737f
C26 drain_right.n11 a_n1180_n5888# 0.037196f
C27 drain_right.n12 a_n1180_n5888# 0.016662f
C28 drain_right.n13 a_n1180_n5888# 0.029285f
C29 drain_right.n14 a_n1180_n5888# 0.015737f
C30 drain_right.n15 a_n1180_n5888# 0.037196f
C31 drain_right.n16 a_n1180_n5888# 0.016662f
C32 drain_right.n17 a_n1180_n5888# 0.029285f
C33 drain_right.n18 a_n1180_n5888# 0.015737f
C34 drain_right.n19 a_n1180_n5888# 0.037196f
C35 drain_right.n20 a_n1180_n5888# 0.016662f
C36 drain_right.n21 a_n1180_n5888# 0.029285f
C37 drain_right.n22 a_n1180_n5888# 0.015737f
C38 drain_right.n23 a_n1180_n5888# 0.037196f
C39 drain_right.n24 a_n1180_n5888# 0.016662f
C40 drain_right.n25 a_n1180_n5888# 0.029285f
C41 drain_right.n26 a_n1180_n5888# 0.015737f
C42 drain_right.n27 a_n1180_n5888# 0.037196f
C43 drain_right.n28 a_n1180_n5888# 0.016662f
C44 drain_right.n29 a_n1180_n5888# 0.029285f
C45 drain_right.n30 a_n1180_n5888# 0.015737f
C46 drain_right.n31 a_n1180_n5888# 0.037196f
C47 drain_right.n32 a_n1180_n5888# 0.016662f
C48 drain_right.n33 a_n1180_n5888# 0.029285f
C49 drain_right.n34 a_n1180_n5888# 0.016199f
C50 drain_right.n35 a_n1180_n5888# 0.037196f
C51 drain_right.n36 a_n1180_n5888# 0.016662f
C52 drain_right.n37 a_n1180_n5888# 0.029285f
C53 drain_right.n38 a_n1180_n5888# 0.015737f
C54 drain_right.n39 a_n1180_n5888# 0.037196f
C55 drain_right.n40 a_n1180_n5888# 0.016662f
C56 drain_right.n41 a_n1180_n5888# 0.029285f
C57 drain_right.n42 a_n1180_n5888# 0.015737f
C58 drain_right.n43 a_n1180_n5888# 0.027897f
C59 drain_right.n44 a_n1180_n5888# 0.026294f
C60 drain_right.t5 a_n1180_n5888# 0.064871f
C61 drain_right.n45 a_n1180_n5888# 0.357305f
C62 drain_right.n46 a_n1180_n5888# 3.17073f
C63 drain_right.n47 a_n1180_n5888# 0.015737f
C64 drain_right.n48 a_n1180_n5888# 0.016662f
C65 drain_right.n49 a_n1180_n5888# 0.037196f
C66 drain_right.n50 a_n1180_n5888# 0.037196f
C67 drain_right.n51 a_n1180_n5888# 0.016662f
C68 drain_right.n52 a_n1180_n5888# 0.015737f
C69 drain_right.n53 a_n1180_n5888# 0.029285f
C70 drain_right.n54 a_n1180_n5888# 0.029285f
C71 drain_right.n55 a_n1180_n5888# 0.015737f
C72 drain_right.n56 a_n1180_n5888# 0.016662f
C73 drain_right.n57 a_n1180_n5888# 0.037196f
C74 drain_right.n58 a_n1180_n5888# 0.037196f
C75 drain_right.n59 a_n1180_n5888# 0.016662f
C76 drain_right.n60 a_n1180_n5888# 0.015737f
C77 drain_right.n61 a_n1180_n5888# 0.029285f
C78 drain_right.n62 a_n1180_n5888# 0.029285f
C79 drain_right.n63 a_n1180_n5888# 0.015737f
C80 drain_right.n64 a_n1180_n5888# 0.015737f
C81 drain_right.n65 a_n1180_n5888# 0.016662f
C82 drain_right.n66 a_n1180_n5888# 0.037196f
C83 drain_right.n67 a_n1180_n5888# 0.037196f
C84 drain_right.n68 a_n1180_n5888# 0.037196f
C85 drain_right.n69 a_n1180_n5888# 0.016199f
C86 drain_right.n70 a_n1180_n5888# 0.015737f
C87 drain_right.n71 a_n1180_n5888# 0.029285f
C88 drain_right.n72 a_n1180_n5888# 0.029285f
C89 drain_right.n73 a_n1180_n5888# 0.015737f
C90 drain_right.n74 a_n1180_n5888# 0.016662f
C91 drain_right.n75 a_n1180_n5888# 0.037196f
C92 drain_right.n76 a_n1180_n5888# 0.037196f
C93 drain_right.n77 a_n1180_n5888# 0.016662f
C94 drain_right.n78 a_n1180_n5888# 0.015737f
C95 drain_right.n79 a_n1180_n5888# 0.029285f
C96 drain_right.n80 a_n1180_n5888# 0.029285f
C97 drain_right.n81 a_n1180_n5888# 0.015737f
C98 drain_right.n82 a_n1180_n5888# 0.016662f
C99 drain_right.n83 a_n1180_n5888# 0.037196f
C100 drain_right.n84 a_n1180_n5888# 0.037196f
C101 drain_right.n85 a_n1180_n5888# 0.016662f
C102 drain_right.n86 a_n1180_n5888# 0.015737f
C103 drain_right.n87 a_n1180_n5888# 0.029285f
C104 drain_right.n88 a_n1180_n5888# 0.029285f
C105 drain_right.n89 a_n1180_n5888# 0.015737f
C106 drain_right.n90 a_n1180_n5888# 0.016662f
C107 drain_right.n91 a_n1180_n5888# 0.037196f
C108 drain_right.n92 a_n1180_n5888# 0.037196f
C109 drain_right.n93 a_n1180_n5888# 0.016662f
C110 drain_right.n94 a_n1180_n5888# 0.015737f
C111 drain_right.n95 a_n1180_n5888# 0.029285f
C112 drain_right.n96 a_n1180_n5888# 0.029285f
C113 drain_right.n97 a_n1180_n5888# 0.015737f
C114 drain_right.n98 a_n1180_n5888# 0.016662f
C115 drain_right.n99 a_n1180_n5888# 0.037196f
C116 drain_right.n100 a_n1180_n5888# 0.037196f
C117 drain_right.n101 a_n1180_n5888# 0.016662f
C118 drain_right.n102 a_n1180_n5888# 0.015737f
C119 drain_right.n103 a_n1180_n5888# 0.029285f
C120 drain_right.n104 a_n1180_n5888# 0.029285f
C121 drain_right.n105 a_n1180_n5888# 0.015737f
C122 drain_right.n106 a_n1180_n5888# 0.016662f
C123 drain_right.n107 a_n1180_n5888# 0.037196f
C124 drain_right.n108 a_n1180_n5888# 0.037196f
C125 drain_right.n109 a_n1180_n5888# 0.037196f
C126 drain_right.n110 a_n1180_n5888# 0.016662f
C127 drain_right.n111 a_n1180_n5888# 0.015737f
C128 drain_right.n112 a_n1180_n5888# 0.029285f
C129 drain_right.n113 a_n1180_n5888# 0.029285f
C130 drain_right.n114 a_n1180_n5888# 0.015737f
C131 drain_right.n115 a_n1180_n5888# 0.016199f
C132 drain_right.n116 a_n1180_n5888# 0.016199f
C133 drain_right.n117 a_n1180_n5888# 0.037196f
C134 drain_right.n118 a_n1180_n5888# 0.037196f
C135 drain_right.n119 a_n1180_n5888# 0.016662f
C136 drain_right.n120 a_n1180_n5888# 0.015737f
C137 drain_right.n121 a_n1180_n5888# 0.029285f
C138 drain_right.n122 a_n1180_n5888# 0.029285f
C139 drain_right.n123 a_n1180_n5888# 0.015737f
C140 drain_right.n124 a_n1180_n5888# 0.016662f
C141 drain_right.n125 a_n1180_n5888# 0.037196f
C142 drain_right.n126 a_n1180_n5888# 0.037196f
C143 drain_right.n127 a_n1180_n5888# 0.016662f
C144 drain_right.n128 a_n1180_n5888# 0.015737f
C145 drain_right.n129 a_n1180_n5888# 0.029285f
C146 drain_right.n130 a_n1180_n5888# 0.029285f
C147 drain_right.n131 a_n1180_n5888# 0.015737f
C148 drain_right.n132 a_n1180_n5888# 0.016662f
C149 drain_right.n133 a_n1180_n5888# 0.037196f
C150 drain_right.n134 a_n1180_n5888# 0.079125f
C151 drain_right.n135 a_n1180_n5888# 0.016662f
C152 drain_right.n136 a_n1180_n5888# 0.015737f
C153 drain_right.n137 a_n1180_n5888# 0.064491f
C154 drain_right.n138 a_n1180_n5888# 0.06486f
C155 drain_right.t3 a_n1180_n5888# 0.578553f
C156 drain_right.t0 a_n1180_n5888# 0.578553f
C157 drain_right.n139 a_n1180_n5888# 5.33237f
C158 drain_right.n140 a_n1180_n5888# 2.53214f
C159 drain_right.t4 a_n1180_n5888# 0.578553f
C160 drain_right.t1 a_n1180_n5888# 0.578553f
C161 drain_right.n141 a_n1180_n5888# 5.33496f
C162 drain_right.n142 a_n1180_n5888# 0.040373f
C163 drain_right.n143 a_n1180_n5888# 0.029285f
C164 drain_right.n144 a_n1180_n5888# 0.015737f
C165 drain_right.n145 a_n1180_n5888# 0.037196f
C166 drain_right.n146 a_n1180_n5888# 0.016662f
C167 drain_right.n147 a_n1180_n5888# 0.029285f
C168 drain_right.n148 a_n1180_n5888# 0.015737f
C169 drain_right.n149 a_n1180_n5888# 0.037196f
C170 drain_right.n150 a_n1180_n5888# 0.016662f
C171 drain_right.n151 a_n1180_n5888# 0.029285f
C172 drain_right.n152 a_n1180_n5888# 0.015737f
C173 drain_right.n153 a_n1180_n5888# 0.037196f
C174 drain_right.n154 a_n1180_n5888# 0.016662f
C175 drain_right.n155 a_n1180_n5888# 0.029285f
C176 drain_right.n156 a_n1180_n5888# 0.015737f
C177 drain_right.n157 a_n1180_n5888# 0.037196f
C178 drain_right.n158 a_n1180_n5888# 0.037196f
C179 drain_right.n159 a_n1180_n5888# 0.016662f
C180 drain_right.n160 a_n1180_n5888# 0.029285f
C181 drain_right.n161 a_n1180_n5888# 0.015737f
C182 drain_right.n162 a_n1180_n5888# 0.037196f
C183 drain_right.n163 a_n1180_n5888# 0.016662f
C184 drain_right.n164 a_n1180_n5888# 0.029285f
C185 drain_right.n165 a_n1180_n5888# 0.015737f
C186 drain_right.n166 a_n1180_n5888# 0.037196f
C187 drain_right.n167 a_n1180_n5888# 0.016662f
C188 drain_right.n168 a_n1180_n5888# 0.029285f
C189 drain_right.n169 a_n1180_n5888# 0.015737f
C190 drain_right.n170 a_n1180_n5888# 0.037196f
C191 drain_right.n171 a_n1180_n5888# 0.016662f
C192 drain_right.n172 a_n1180_n5888# 0.029285f
C193 drain_right.n173 a_n1180_n5888# 0.015737f
C194 drain_right.n174 a_n1180_n5888# 0.037196f
C195 drain_right.n175 a_n1180_n5888# 0.016662f
C196 drain_right.n176 a_n1180_n5888# 0.029285f
C197 drain_right.n177 a_n1180_n5888# 0.016199f
C198 drain_right.n178 a_n1180_n5888# 0.037196f
C199 drain_right.n179 a_n1180_n5888# 0.015737f
C200 drain_right.n180 a_n1180_n5888# 0.016662f
C201 drain_right.n181 a_n1180_n5888# 0.029285f
C202 drain_right.n182 a_n1180_n5888# 0.015737f
C203 drain_right.n183 a_n1180_n5888# 0.037196f
C204 drain_right.n184 a_n1180_n5888# 0.016662f
C205 drain_right.n185 a_n1180_n5888# 0.029285f
C206 drain_right.n186 a_n1180_n5888# 0.015737f
C207 drain_right.n187 a_n1180_n5888# 0.027897f
C208 drain_right.n188 a_n1180_n5888# 0.026294f
C209 drain_right.t2 a_n1180_n5888# 0.064871f
C210 drain_right.n189 a_n1180_n5888# 0.357305f
C211 drain_right.n190 a_n1180_n5888# 3.17073f
C212 drain_right.n191 a_n1180_n5888# 0.015737f
C213 drain_right.n192 a_n1180_n5888# 0.016662f
C214 drain_right.n193 a_n1180_n5888# 0.037196f
C215 drain_right.n194 a_n1180_n5888# 0.037196f
C216 drain_right.n195 a_n1180_n5888# 0.016662f
C217 drain_right.n196 a_n1180_n5888# 0.015737f
C218 drain_right.n197 a_n1180_n5888# 0.029285f
C219 drain_right.n198 a_n1180_n5888# 0.029285f
C220 drain_right.n199 a_n1180_n5888# 0.015737f
C221 drain_right.n200 a_n1180_n5888# 0.016662f
C222 drain_right.n201 a_n1180_n5888# 0.037196f
C223 drain_right.n202 a_n1180_n5888# 0.037196f
C224 drain_right.n203 a_n1180_n5888# 0.016662f
C225 drain_right.n204 a_n1180_n5888# 0.015737f
C226 drain_right.n205 a_n1180_n5888# 0.029285f
C227 drain_right.n206 a_n1180_n5888# 0.029285f
C228 drain_right.n207 a_n1180_n5888# 0.015737f
C229 drain_right.n208 a_n1180_n5888# 0.016662f
C230 drain_right.n209 a_n1180_n5888# 0.037196f
C231 drain_right.n210 a_n1180_n5888# 0.037196f
C232 drain_right.n211 a_n1180_n5888# 0.037196f
C233 drain_right.n212 a_n1180_n5888# 0.016199f
C234 drain_right.n213 a_n1180_n5888# 0.015737f
C235 drain_right.n214 a_n1180_n5888# 0.029285f
C236 drain_right.n215 a_n1180_n5888# 0.029285f
C237 drain_right.n216 a_n1180_n5888# 0.015737f
C238 drain_right.n217 a_n1180_n5888# 0.016662f
C239 drain_right.n218 a_n1180_n5888# 0.037196f
C240 drain_right.n219 a_n1180_n5888# 0.037196f
C241 drain_right.n220 a_n1180_n5888# 0.016662f
C242 drain_right.n221 a_n1180_n5888# 0.015737f
C243 drain_right.n222 a_n1180_n5888# 0.029285f
C244 drain_right.n223 a_n1180_n5888# 0.029285f
C245 drain_right.n224 a_n1180_n5888# 0.015737f
C246 drain_right.n225 a_n1180_n5888# 0.016662f
C247 drain_right.n226 a_n1180_n5888# 0.037196f
C248 drain_right.n227 a_n1180_n5888# 0.037196f
C249 drain_right.n228 a_n1180_n5888# 0.016662f
C250 drain_right.n229 a_n1180_n5888# 0.015737f
C251 drain_right.n230 a_n1180_n5888# 0.029285f
C252 drain_right.n231 a_n1180_n5888# 0.029285f
C253 drain_right.n232 a_n1180_n5888# 0.015737f
C254 drain_right.n233 a_n1180_n5888# 0.016662f
C255 drain_right.n234 a_n1180_n5888# 0.037196f
C256 drain_right.n235 a_n1180_n5888# 0.037196f
C257 drain_right.n236 a_n1180_n5888# 0.016662f
C258 drain_right.n237 a_n1180_n5888# 0.015737f
C259 drain_right.n238 a_n1180_n5888# 0.029285f
C260 drain_right.n239 a_n1180_n5888# 0.029285f
C261 drain_right.n240 a_n1180_n5888# 0.015737f
C262 drain_right.n241 a_n1180_n5888# 0.016662f
C263 drain_right.n242 a_n1180_n5888# 0.037196f
C264 drain_right.n243 a_n1180_n5888# 0.037196f
C265 drain_right.n244 a_n1180_n5888# 0.016662f
C266 drain_right.n245 a_n1180_n5888# 0.015737f
C267 drain_right.n246 a_n1180_n5888# 0.029285f
C268 drain_right.n247 a_n1180_n5888# 0.029285f
C269 drain_right.n248 a_n1180_n5888# 0.015737f
C270 drain_right.n249 a_n1180_n5888# 0.016662f
C271 drain_right.n250 a_n1180_n5888# 0.037196f
C272 drain_right.n251 a_n1180_n5888# 0.037196f
C273 drain_right.n252 a_n1180_n5888# 0.016662f
C274 drain_right.n253 a_n1180_n5888# 0.015737f
C275 drain_right.n254 a_n1180_n5888# 0.029285f
C276 drain_right.n255 a_n1180_n5888# 0.029285f
C277 drain_right.n256 a_n1180_n5888# 0.015737f
C278 drain_right.n257 a_n1180_n5888# 0.016199f
C279 drain_right.n258 a_n1180_n5888# 0.016199f
C280 drain_right.n259 a_n1180_n5888# 0.037196f
C281 drain_right.n260 a_n1180_n5888# 0.037196f
C282 drain_right.n261 a_n1180_n5888# 0.016662f
C283 drain_right.n262 a_n1180_n5888# 0.015737f
C284 drain_right.n263 a_n1180_n5888# 0.029285f
C285 drain_right.n264 a_n1180_n5888# 0.029285f
C286 drain_right.n265 a_n1180_n5888# 0.015737f
C287 drain_right.n266 a_n1180_n5888# 0.016662f
C288 drain_right.n267 a_n1180_n5888# 0.037196f
C289 drain_right.n268 a_n1180_n5888# 0.037196f
C290 drain_right.n269 a_n1180_n5888# 0.016662f
C291 drain_right.n270 a_n1180_n5888# 0.015737f
C292 drain_right.n271 a_n1180_n5888# 0.029285f
C293 drain_right.n272 a_n1180_n5888# 0.029285f
C294 drain_right.n273 a_n1180_n5888# 0.015737f
C295 drain_right.n274 a_n1180_n5888# 0.016662f
C296 drain_right.n275 a_n1180_n5888# 0.037196f
C297 drain_right.n276 a_n1180_n5888# 0.079125f
C298 drain_right.n277 a_n1180_n5888# 0.016662f
C299 drain_right.n278 a_n1180_n5888# 0.015737f
C300 drain_right.n279 a_n1180_n5888# 0.064491f
C301 drain_right.n280 a_n1180_n5888# 0.064277f
C302 drain_right.n281 a_n1180_n5888# 0.693643f
C303 minus.t4 a_n1180_n5888# 1.06626f
C304 minus.n0 a_n1180_n5888# 0.407129f
C305 minus.t3 a_n1180_n5888# 1.06626f
C306 minus.t1 a_n1180_n5888# 1.05896f
C307 minus.n1 a_n1180_n5888# 0.388426f
C308 minus.n2 a_n1180_n5888# 0.407041f
C309 minus.n3 a_n1180_n5888# 2.87505f
C310 minus.t0 a_n1180_n5888# 1.06626f
C311 minus.n4 a_n1180_n5888# 0.407129f
C312 minus.t2 a_n1180_n5888# 1.05896f
C313 minus.n5 a_n1180_n5888# 0.388426f
C314 minus.t5 a_n1180_n5888# 1.06626f
C315 minus.n6 a_n1180_n5888# 0.407041f
C316 minus.n7 a_n1180_n5888# 0.466961f
C317 minus.n8 a_n1180_n5888# 3.33028f
C318 source.n0 a_n1180_n5888# 0.040174f
C319 source.n1 a_n1180_n5888# 0.029141f
C320 source.n2 a_n1180_n5888# 0.015659f
C321 source.n3 a_n1180_n5888# 0.037012f
C322 source.n4 a_n1180_n5888# 0.01658f
C323 source.n5 a_n1180_n5888# 0.029141f
C324 source.n6 a_n1180_n5888# 0.015659f
C325 source.n7 a_n1180_n5888# 0.037012f
C326 source.n8 a_n1180_n5888# 0.01658f
C327 source.n9 a_n1180_n5888# 0.029141f
C328 source.n10 a_n1180_n5888# 0.015659f
C329 source.n11 a_n1180_n5888# 0.037012f
C330 source.n12 a_n1180_n5888# 0.01658f
C331 source.n13 a_n1180_n5888# 0.029141f
C332 source.n14 a_n1180_n5888# 0.015659f
C333 source.n15 a_n1180_n5888# 0.037012f
C334 source.n16 a_n1180_n5888# 0.037012f
C335 source.n17 a_n1180_n5888# 0.01658f
C336 source.n18 a_n1180_n5888# 0.029141f
C337 source.n19 a_n1180_n5888# 0.015659f
C338 source.n20 a_n1180_n5888# 0.037012f
C339 source.n21 a_n1180_n5888# 0.01658f
C340 source.n22 a_n1180_n5888# 0.029141f
C341 source.n23 a_n1180_n5888# 0.015659f
C342 source.n24 a_n1180_n5888# 0.037012f
C343 source.n25 a_n1180_n5888# 0.01658f
C344 source.n26 a_n1180_n5888# 0.029141f
C345 source.n27 a_n1180_n5888# 0.015659f
C346 source.n28 a_n1180_n5888# 0.037012f
C347 source.n29 a_n1180_n5888# 0.01658f
C348 source.n30 a_n1180_n5888# 0.029141f
C349 source.n31 a_n1180_n5888# 0.015659f
C350 source.n32 a_n1180_n5888# 0.037012f
C351 source.n33 a_n1180_n5888# 0.01658f
C352 source.n34 a_n1180_n5888# 0.029141f
C353 source.n35 a_n1180_n5888# 0.01612f
C354 source.n36 a_n1180_n5888# 0.037012f
C355 source.n37 a_n1180_n5888# 0.015659f
C356 source.n38 a_n1180_n5888# 0.01658f
C357 source.n39 a_n1180_n5888# 0.029141f
C358 source.n40 a_n1180_n5888# 0.015659f
C359 source.n41 a_n1180_n5888# 0.037012f
C360 source.n42 a_n1180_n5888# 0.01658f
C361 source.n43 a_n1180_n5888# 0.029141f
C362 source.n44 a_n1180_n5888# 0.015659f
C363 source.n45 a_n1180_n5888# 0.027759f
C364 source.n46 a_n1180_n5888# 0.026165f
C365 source.t9 a_n1180_n5888# 0.064552f
C366 source.n47 a_n1180_n5888# 0.355545f
C367 source.n48 a_n1180_n5888# 3.15511f
C368 source.n49 a_n1180_n5888# 0.015659f
C369 source.n50 a_n1180_n5888# 0.01658f
C370 source.n51 a_n1180_n5888# 0.037012f
C371 source.n52 a_n1180_n5888# 0.037012f
C372 source.n53 a_n1180_n5888# 0.01658f
C373 source.n54 a_n1180_n5888# 0.015659f
C374 source.n55 a_n1180_n5888# 0.029141f
C375 source.n56 a_n1180_n5888# 0.029141f
C376 source.n57 a_n1180_n5888# 0.015659f
C377 source.n58 a_n1180_n5888# 0.01658f
C378 source.n59 a_n1180_n5888# 0.037012f
C379 source.n60 a_n1180_n5888# 0.037012f
C380 source.n61 a_n1180_n5888# 0.01658f
C381 source.n62 a_n1180_n5888# 0.015659f
C382 source.n63 a_n1180_n5888# 0.029141f
C383 source.n64 a_n1180_n5888# 0.029141f
C384 source.n65 a_n1180_n5888# 0.015659f
C385 source.n66 a_n1180_n5888# 0.01658f
C386 source.n67 a_n1180_n5888# 0.037012f
C387 source.n68 a_n1180_n5888# 0.037012f
C388 source.n69 a_n1180_n5888# 0.037012f
C389 source.n70 a_n1180_n5888# 0.01612f
C390 source.n71 a_n1180_n5888# 0.015659f
C391 source.n72 a_n1180_n5888# 0.029141f
C392 source.n73 a_n1180_n5888# 0.029141f
C393 source.n74 a_n1180_n5888# 0.015659f
C394 source.n75 a_n1180_n5888# 0.01658f
C395 source.n76 a_n1180_n5888# 0.037012f
C396 source.n77 a_n1180_n5888# 0.037012f
C397 source.n78 a_n1180_n5888# 0.01658f
C398 source.n79 a_n1180_n5888# 0.015659f
C399 source.n80 a_n1180_n5888# 0.029141f
C400 source.n81 a_n1180_n5888# 0.029141f
C401 source.n82 a_n1180_n5888# 0.015659f
C402 source.n83 a_n1180_n5888# 0.01658f
C403 source.n84 a_n1180_n5888# 0.037012f
C404 source.n85 a_n1180_n5888# 0.037012f
C405 source.n86 a_n1180_n5888# 0.01658f
C406 source.n87 a_n1180_n5888# 0.015659f
C407 source.n88 a_n1180_n5888# 0.029141f
C408 source.n89 a_n1180_n5888# 0.029141f
C409 source.n90 a_n1180_n5888# 0.015659f
C410 source.n91 a_n1180_n5888# 0.01658f
C411 source.n92 a_n1180_n5888# 0.037012f
C412 source.n93 a_n1180_n5888# 0.037012f
C413 source.n94 a_n1180_n5888# 0.01658f
C414 source.n95 a_n1180_n5888# 0.015659f
C415 source.n96 a_n1180_n5888# 0.029141f
C416 source.n97 a_n1180_n5888# 0.029141f
C417 source.n98 a_n1180_n5888# 0.015659f
C418 source.n99 a_n1180_n5888# 0.01658f
C419 source.n100 a_n1180_n5888# 0.037012f
C420 source.n101 a_n1180_n5888# 0.037012f
C421 source.n102 a_n1180_n5888# 0.01658f
C422 source.n103 a_n1180_n5888# 0.015659f
C423 source.n104 a_n1180_n5888# 0.029141f
C424 source.n105 a_n1180_n5888# 0.029141f
C425 source.n106 a_n1180_n5888# 0.015659f
C426 source.n107 a_n1180_n5888# 0.01658f
C427 source.n108 a_n1180_n5888# 0.037012f
C428 source.n109 a_n1180_n5888# 0.037012f
C429 source.n110 a_n1180_n5888# 0.01658f
C430 source.n111 a_n1180_n5888# 0.015659f
C431 source.n112 a_n1180_n5888# 0.029141f
C432 source.n113 a_n1180_n5888# 0.029141f
C433 source.n114 a_n1180_n5888# 0.015659f
C434 source.n115 a_n1180_n5888# 0.01612f
C435 source.n116 a_n1180_n5888# 0.01612f
C436 source.n117 a_n1180_n5888# 0.037012f
C437 source.n118 a_n1180_n5888# 0.037012f
C438 source.n119 a_n1180_n5888# 0.01658f
C439 source.n120 a_n1180_n5888# 0.015659f
C440 source.n121 a_n1180_n5888# 0.029141f
C441 source.n122 a_n1180_n5888# 0.029141f
C442 source.n123 a_n1180_n5888# 0.015659f
C443 source.n124 a_n1180_n5888# 0.01658f
C444 source.n125 a_n1180_n5888# 0.037012f
C445 source.n126 a_n1180_n5888# 0.037012f
C446 source.n127 a_n1180_n5888# 0.01658f
C447 source.n128 a_n1180_n5888# 0.015659f
C448 source.n129 a_n1180_n5888# 0.029141f
C449 source.n130 a_n1180_n5888# 0.029141f
C450 source.n131 a_n1180_n5888# 0.015659f
C451 source.n132 a_n1180_n5888# 0.01658f
C452 source.n133 a_n1180_n5888# 0.037012f
C453 source.n134 a_n1180_n5888# 0.078735f
C454 source.n135 a_n1180_n5888# 0.01658f
C455 source.n136 a_n1180_n5888# 0.015659f
C456 source.n137 a_n1180_n5888# 0.064173f
C457 source.n138 a_n1180_n5888# 0.043812f
C458 source.n139 a_n1180_n5888# 2.28399f
C459 source.t10 a_n1180_n5888# 0.575702f
C460 source.t11 a_n1180_n5888# 0.575702f
C461 source.n140 a_n1180_n5888# 5.21019f
C462 source.n141 a_n1180_n5888# 0.41679f
C463 source.n142 a_n1180_n5888# 0.040174f
C464 source.n143 a_n1180_n5888# 0.029141f
C465 source.n144 a_n1180_n5888# 0.015659f
C466 source.n145 a_n1180_n5888# 0.037012f
C467 source.n146 a_n1180_n5888# 0.01658f
C468 source.n147 a_n1180_n5888# 0.029141f
C469 source.n148 a_n1180_n5888# 0.015659f
C470 source.n149 a_n1180_n5888# 0.037012f
C471 source.n150 a_n1180_n5888# 0.01658f
C472 source.n151 a_n1180_n5888# 0.029141f
C473 source.n152 a_n1180_n5888# 0.015659f
C474 source.n153 a_n1180_n5888# 0.037012f
C475 source.n154 a_n1180_n5888# 0.01658f
C476 source.n155 a_n1180_n5888# 0.029141f
C477 source.n156 a_n1180_n5888# 0.015659f
C478 source.n157 a_n1180_n5888# 0.037012f
C479 source.n158 a_n1180_n5888# 0.037012f
C480 source.n159 a_n1180_n5888# 0.01658f
C481 source.n160 a_n1180_n5888# 0.029141f
C482 source.n161 a_n1180_n5888# 0.015659f
C483 source.n162 a_n1180_n5888# 0.037012f
C484 source.n163 a_n1180_n5888# 0.01658f
C485 source.n164 a_n1180_n5888# 0.029141f
C486 source.n165 a_n1180_n5888# 0.015659f
C487 source.n166 a_n1180_n5888# 0.037012f
C488 source.n167 a_n1180_n5888# 0.01658f
C489 source.n168 a_n1180_n5888# 0.029141f
C490 source.n169 a_n1180_n5888# 0.015659f
C491 source.n170 a_n1180_n5888# 0.037012f
C492 source.n171 a_n1180_n5888# 0.01658f
C493 source.n172 a_n1180_n5888# 0.029141f
C494 source.n173 a_n1180_n5888# 0.015659f
C495 source.n174 a_n1180_n5888# 0.037012f
C496 source.n175 a_n1180_n5888# 0.01658f
C497 source.n176 a_n1180_n5888# 0.029141f
C498 source.n177 a_n1180_n5888# 0.01612f
C499 source.n178 a_n1180_n5888# 0.037012f
C500 source.n179 a_n1180_n5888# 0.015659f
C501 source.n180 a_n1180_n5888# 0.01658f
C502 source.n181 a_n1180_n5888# 0.029141f
C503 source.n182 a_n1180_n5888# 0.015659f
C504 source.n183 a_n1180_n5888# 0.037012f
C505 source.n184 a_n1180_n5888# 0.01658f
C506 source.n185 a_n1180_n5888# 0.029141f
C507 source.n186 a_n1180_n5888# 0.015659f
C508 source.n187 a_n1180_n5888# 0.027759f
C509 source.n188 a_n1180_n5888# 0.026165f
C510 source.t5 a_n1180_n5888# 0.064552f
C511 source.n189 a_n1180_n5888# 0.355545f
C512 source.n190 a_n1180_n5888# 3.15511f
C513 source.n191 a_n1180_n5888# 0.015659f
C514 source.n192 a_n1180_n5888# 0.01658f
C515 source.n193 a_n1180_n5888# 0.037012f
C516 source.n194 a_n1180_n5888# 0.037012f
C517 source.n195 a_n1180_n5888# 0.01658f
C518 source.n196 a_n1180_n5888# 0.015659f
C519 source.n197 a_n1180_n5888# 0.029141f
C520 source.n198 a_n1180_n5888# 0.029141f
C521 source.n199 a_n1180_n5888# 0.015659f
C522 source.n200 a_n1180_n5888# 0.01658f
C523 source.n201 a_n1180_n5888# 0.037012f
C524 source.n202 a_n1180_n5888# 0.037012f
C525 source.n203 a_n1180_n5888# 0.01658f
C526 source.n204 a_n1180_n5888# 0.015659f
C527 source.n205 a_n1180_n5888# 0.029141f
C528 source.n206 a_n1180_n5888# 0.029141f
C529 source.n207 a_n1180_n5888# 0.015659f
C530 source.n208 a_n1180_n5888# 0.01658f
C531 source.n209 a_n1180_n5888# 0.037012f
C532 source.n210 a_n1180_n5888# 0.037012f
C533 source.n211 a_n1180_n5888# 0.037012f
C534 source.n212 a_n1180_n5888# 0.01612f
C535 source.n213 a_n1180_n5888# 0.015659f
C536 source.n214 a_n1180_n5888# 0.029141f
C537 source.n215 a_n1180_n5888# 0.029141f
C538 source.n216 a_n1180_n5888# 0.015659f
C539 source.n217 a_n1180_n5888# 0.01658f
C540 source.n218 a_n1180_n5888# 0.037012f
C541 source.n219 a_n1180_n5888# 0.037012f
C542 source.n220 a_n1180_n5888# 0.01658f
C543 source.n221 a_n1180_n5888# 0.015659f
C544 source.n222 a_n1180_n5888# 0.029141f
C545 source.n223 a_n1180_n5888# 0.029141f
C546 source.n224 a_n1180_n5888# 0.015659f
C547 source.n225 a_n1180_n5888# 0.01658f
C548 source.n226 a_n1180_n5888# 0.037012f
C549 source.n227 a_n1180_n5888# 0.037012f
C550 source.n228 a_n1180_n5888# 0.01658f
C551 source.n229 a_n1180_n5888# 0.015659f
C552 source.n230 a_n1180_n5888# 0.029141f
C553 source.n231 a_n1180_n5888# 0.029141f
C554 source.n232 a_n1180_n5888# 0.015659f
C555 source.n233 a_n1180_n5888# 0.01658f
C556 source.n234 a_n1180_n5888# 0.037012f
C557 source.n235 a_n1180_n5888# 0.037012f
C558 source.n236 a_n1180_n5888# 0.01658f
C559 source.n237 a_n1180_n5888# 0.015659f
C560 source.n238 a_n1180_n5888# 0.029141f
C561 source.n239 a_n1180_n5888# 0.029141f
C562 source.n240 a_n1180_n5888# 0.015659f
C563 source.n241 a_n1180_n5888# 0.01658f
C564 source.n242 a_n1180_n5888# 0.037012f
C565 source.n243 a_n1180_n5888# 0.037012f
C566 source.n244 a_n1180_n5888# 0.01658f
C567 source.n245 a_n1180_n5888# 0.015659f
C568 source.n246 a_n1180_n5888# 0.029141f
C569 source.n247 a_n1180_n5888# 0.029141f
C570 source.n248 a_n1180_n5888# 0.015659f
C571 source.n249 a_n1180_n5888# 0.01658f
C572 source.n250 a_n1180_n5888# 0.037012f
C573 source.n251 a_n1180_n5888# 0.037012f
C574 source.n252 a_n1180_n5888# 0.01658f
C575 source.n253 a_n1180_n5888# 0.015659f
C576 source.n254 a_n1180_n5888# 0.029141f
C577 source.n255 a_n1180_n5888# 0.029141f
C578 source.n256 a_n1180_n5888# 0.015659f
C579 source.n257 a_n1180_n5888# 0.01612f
C580 source.n258 a_n1180_n5888# 0.01612f
C581 source.n259 a_n1180_n5888# 0.037012f
C582 source.n260 a_n1180_n5888# 0.037012f
C583 source.n261 a_n1180_n5888# 0.01658f
C584 source.n262 a_n1180_n5888# 0.015659f
C585 source.n263 a_n1180_n5888# 0.029141f
C586 source.n264 a_n1180_n5888# 0.029141f
C587 source.n265 a_n1180_n5888# 0.015659f
C588 source.n266 a_n1180_n5888# 0.01658f
C589 source.n267 a_n1180_n5888# 0.037012f
C590 source.n268 a_n1180_n5888# 0.037012f
C591 source.n269 a_n1180_n5888# 0.01658f
C592 source.n270 a_n1180_n5888# 0.015659f
C593 source.n271 a_n1180_n5888# 0.029141f
C594 source.n272 a_n1180_n5888# 0.029141f
C595 source.n273 a_n1180_n5888# 0.015659f
C596 source.n274 a_n1180_n5888# 0.01658f
C597 source.n275 a_n1180_n5888# 0.037012f
C598 source.n276 a_n1180_n5888# 0.078735f
C599 source.n277 a_n1180_n5888# 0.01658f
C600 source.n278 a_n1180_n5888# 0.015659f
C601 source.n279 a_n1180_n5888# 0.064173f
C602 source.n280 a_n1180_n5888# 0.043812f
C603 source.n281 a_n1180_n5888# 0.137634f
C604 source.t0 a_n1180_n5888# 0.575702f
C605 source.t3 a_n1180_n5888# 0.575702f
C606 source.n282 a_n1180_n5888# 5.21019f
C607 source.n283 a_n1180_n5888# 3.14736f
C608 source.t8 a_n1180_n5888# 0.575702f
C609 source.t7 a_n1180_n5888# 0.575702f
C610 source.n284 a_n1180_n5888# 5.21019f
C611 source.n285 a_n1180_n5888# 3.14737f
C612 source.n286 a_n1180_n5888# 0.040174f
C613 source.n287 a_n1180_n5888# 0.029141f
C614 source.n288 a_n1180_n5888# 0.015659f
C615 source.n289 a_n1180_n5888# 0.037012f
C616 source.n290 a_n1180_n5888# 0.01658f
C617 source.n291 a_n1180_n5888# 0.029141f
C618 source.n292 a_n1180_n5888# 0.015659f
C619 source.n293 a_n1180_n5888# 0.037012f
C620 source.n294 a_n1180_n5888# 0.01658f
C621 source.n295 a_n1180_n5888# 0.029141f
C622 source.n296 a_n1180_n5888# 0.015659f
C623 source.n297 a_n1180_n5888# 0.037012f
C624 source.n298 a_n1180_n5888# 0.01658f
C625 source.n299 a_n1180_n5888# 0.029141f
C626 source.n300 a_n1180_n5888# 0.015659f
C627 source.n301 a_n1180_n5888# 0.037012f
C628 source.n302 a_n1180_n5888# 0.01658f
C629 source.n303 a_n1180_n5888# 0.029141f
C630 source.n304 a_n1180_n5888# 0.015659f
C631 source.n305 a_n1180_n5888# 0.037012f
C632 source.n306 a_n1180_n5888# 0.01658f
C633 source.n307 a_n1180_n5888# 0.029141f
C634 source.n308 a_n1180_n5888# 0.015659f
C635 source.n309 a_n1180_n5888# 0.037012f
C636 source.n310 a_n1180_n5888# 0.01658f
C637 source.n311 a_n1180_n5888# 0.029141f
C638 source.n312 a_n1180_n5888# 0.015659f
C639 source.n313 a_n1180_n5888# 0.037012f
C640 source.n314 a_n1180_n5888# 0.01658f
C641 source.n315 a_n1180_n5888# 0.029141f
C642 source.n316 a_n1180_n5888# 0.015659f
C643 source.n317 a_n1180_n5888# 0.037012f
C644 source.n318 a_n1180_n5888# 0.01658f
C645 source.n319 a_n1180_n5888# 0.029141f
C646 source.n320 a_n1180_n5888# 0.01612f
C647 source.n321 a_n1180_n5888# 0.037012f
C648 source.n322 a_n1180_n5888# 0.01658f
C649 source.n323 a_n1180_n5888# 0.029141f
C650 source.n324 a_n1180_n5888# 0.015659f
C651 source.n325 a_n1180_n5888# 0.037012f
C652 source.n326 a_n1180_n5888# 0.01658f
C653 source.n327 a_n1180_n5888# 0.029141f
C654 source.n328 a_n1180_n5888# 0.015659f
C655 source.n329 a_n1180_n5888# 0.027759f
C656 source.n330 a_n1180_n5888# 0.026165f
C657 source.t6 a_n1180_n5888# 0.064552f
C658 source.n331 a_n1180_n5888# 0.355545f
C659 source.n332 a_n1180_n5888# 3.15511f
C660 source.n333 a_n1180_n5888# 0.015659f
C661 source.n334 a_n1180_n5888# 0.01658f
C662 source.n335 a_n1180_n5888# 0.037012f
C663 source.n336 a_n1180_n5888# 0.037012f
C664 source.n337 a_n1180_n5888# 0.01658f
C665 source.n338 a_n1180_n5888# 0.015659f
C666 source.n339 a_n1180_n5888# 0.029141f
C667 source.n340 a_n1180_n5888# 0.029141f
C668 source.n341 a_n1180_n5888# 0.015659f
C669 source.n342 a_n1180_n5888# 0.01658f
C670 source.n343 a_n1180_n5888# 0.037012f
C671 source.n344 a_n1180_n5888# 0.037012f
C672 source.n345 a_n1180_n5888# 0.01658f
C673 source.n346 a_n1180_n5888# 0.015659f
C674 source.n347 a_n1180_n5888# 0.029141f
C675 source.n348 a_n1180_n5888# 0.029141f
C676 source.n349 a_n1180_n5888# 0.015659f
C677 source.n350 a_n1180_n5888# 0.015659f
C678 source.n351 a_n1180_n5888# 0.01658f
C679 source.n352 a_n1180_n5888# 0.037012f
C680 source.n353 a_n1180_n5888# 0.037012f
C681 source.n354 a_n1180_n5888# 0.037012f
C682 source.n355 a_n1180_n5888# 0.01612f
C683 source.n356 a_n1180_n5888# 0.015659f
C684 source.n357 a_n1180_n5888# 0.029141f
C685 source.n358 a_n1180_n5888# 0.029141f
C686 source.n359 a_n1180_n5888# 0.015659f
C687 source.n360 a_n1180_n5888# 0.01658f
C688 source.n361 a_n1180_n5888# 0.037012f
C689 source.n362 a_n1180_n5888# 0.037012f
C690 source.n363 a_n1180_n5888# 0.01658f
C691 source.n364 a_n1180_n5888# 0.015659f
C692 source.n365 a_n1180_n5888# 0.029141f
C693 source.n366 a_n1180_n5888# 0.029141f
C694 source.n367 a_n1180_n5888# 0.015659f
C695 source.n368 a_n1180_n5888# 0.01658f
C696 source.n369 a_n1180_n5888# 0.037012f
C697 source.n370 a_n1180_n5888# 0.037012f
C698 source.n371 a_n1180_n5888# 0.01658f
C699 source.n372 a_n1180_n5888# 0.015659f
C700 source.n373 a_n1180_n5888# 0.029141f
C701 source.n374 a_n1180_n5888# 0.029141f
C702 source.n375 a_n1180_n5888# 0.015659f
C703 source.n376 a_n1180_n5888# 0.01658f
C704 source.n377 a_n1180_n5888# 0.037012f
C705 source.n378 a_n1180_n5888# 0.037012f
C706 source.n379 a_n1180_n5888# 0.01658f
C707 source.n380 a_n1180_n5888# 0.015659f
C708 source.n381 a_n1180_n5888# 0.029141f
C709 source.n382 a_n1180_n5888# 0.029141f
C710 source.n383 a_n1180_n5888# 0.015659f
C711 source.n384 a_n1180_n5888# 0.01658f
C712 source.n385 a_n1180_n5888# 0.037012f
C713 source.n386 a_n1180_n5888# 0.037012f
C714 source.n387 a_n1180_n5888# 0.01658f
C715 source.n388 a_n1180_n5888# 0.015659f
C716 source.n389 a_n1180_n5888# 0.029141f
C717 source.n390 a_n1180_n5888# 0.029141f
C718 source.n391 a_n1180_n5888# 0.015659f
C719 source.n392 a_n1180_n5888# 0.01658f
C720 source.n393 a_n1180_n5888# 0.037012f
C721 source.n394 a_n1180_n5888# 0.037012f
C722 source.n395 a_n1180_n5888# 0.037012f
C723 source.n396 a_n1180_n5888# 0.01658f
C724 source.n397 a_n1180_n5888# 0.015659f
C725 source.n398 a_n1180_n5888# 0.029141f
C726 source.n399 a_n1180_n5888# 0.029141f
C727 source.n400 a_n1180_n5888# 0.015659f
C728 source.n401 a_n1180_n5888# 0.01612f
C729 source.n402 a_n1180_n5888# 0.01612f
C730 source.n403 a_n1180_n5888# 0.037012f
C731 source.n404 a_n1180_n5888# 0.037012f
C732 source.n405 a_n1180_n5888# 0.01658f
C733 source.n406 a_n1180_n5888# 0.015659f
C734 source.n407 a_n1180_n5888# 0.029141f
C735 source.n408 a_n1180_n5888# 0.029141f
C736 source.n409 a_n1180_n5888# 0.015659f
C737 source.n410 a_n1180_n5888# 0.01658f
C738 source.n411 a_n1180_n5888# 0.037012f
C739 source.n412 a_n1180_n5888# 0.037012f
C740 source.n413 a_n1180_n5888# 0.01658f
C741 source.n414 a_n1180_n5888# 0.015659f
C742 source.n415 a_n1180_n5888# 0.029141f
C743 source.n416 a_n1180_n5888# 0.029141f
C744 source.n417 a_n1180_n5888# 0.015659f
C745 source.n418 a_n1180_n5888# 0.01658f
C746 source.n419 a_n1180_n5888# 0.037012f
C747 source.n420 a_n1180_n5888# 0.078735f
C748 source.n421 a_n1180_n5888# 0.01658f
C749 source.n422 a_n1180_n5888# 0.015659f
C750 source.n423 a_n1180_n5888# 0.064173f
C751 source.n424 a_n1180_n5888# 0.043812f
C752 source.n425 a_n1180_n5888# 0.137634f
C753 source.t2 a_n1180_n5888# 0.575702f
C754 source.t1 a_n1180_n5888# 0.575702f
C755 source.n426 a_n1180_n5888# 5.21019f
C756 source.n427 a_n1180_n5888# 0.416792f
C757 source.n428 a_n1180_n5888# 0.040174f
C758 source.n429 a_n1180_n5888# 0.029141f
C759 source.n430 a_n1180_n5888# 0.015659f
C760 source.n431 a_n1180_n5888# 0.037012f
C761 source.n432 a_n1180_n5888# 0.01658f
C762 source.n433 a_n1180_n5888# 0.029141f
C763 source.n434 a_n1180_n5888# 0.015659f
C764 source.n435 a_n1180_n5888# 0.037012f
C765 source.n436 a_n1180_n5888# 0.01658f
C766 source.n437 a_n1180_n5888# 0.029141f
C767 source.n438 a_n1180_n5888# 0.015659f
C768 source.n439 a_n1180_n5888# 0.037012f
C769 source.n440 a_n1180_n5888# 0.01658f
C770 source.n441 a_n1180_n5888# 0.029141f
C771 source.n442 a_n1180_n5888# 0.015659f
C772 source.n443 a_n1180_n5888# 0.037012f
C773 source.n444 a_n1180_n5888# 0.01658f
C774 source.n445 a_n1180_n5888# 0.029141f
C775 source.n446 a_n1180_n5888# 0.015659f
C776 source.n447 a_n1180_n5888# 0.037012f
C777 source.n448 a_n1180_n5888# 0.01658f
C778 source.n449 a_n1180_n5888# 0.029141f
C779 source.n450 a_n1180_n5888# 0.015659f
C780 source.n451 a_n1180_n5888# 0.037012f
C781 source.n452 a_n1180_n5888# 0.01658f
C782 source.n453 a_n1180_n5888# 0.029141f
C783 source.n454 a_n1180_n5888# 0.015659f
C784 source.n455 a_n1180_n5888# 0.037012f
C785 source.n456 a_n1180_n5888# 0.01658f
C786 source.n457 a_n1180_n5888# 0.029141f
C787 source.n458 a_n1180_n5888# 0.015659f
C788 source.n459 a_n1180_n5888# 0.037012f
C789 source.n460 a_n1180_n5888# 0.01658f
C790 source.n461 a_n1180_n5888# 0.029141f
C791 source.n462 a_n1180_n5888# 0.01612f
C792 source.n463 a_n1180_n5888# 0.037012f
C793 source.n464 a_n1180_n5888# 0.01658f
C794 source.n465 a_n1180_n5888# 0.029141f
C795 source.n466 a_n1180_n5888# 0.015659f
C796 source.n467 a_n1180_n5888# 0.037012f
C797 source.n468 a_n1180_n5888# 0.01658f
C798 source.n469 a_n1180_n5888# 0.029141f
C799 source.n470 a_n1180_n5888# 0.015659f
C800 source.n471 a_n1180_n5888# 0.027759f
C801 source.n472 a_n1180_n5888# 0.026165f
C802 source.t4 a_n1180_n5888# 0.064552f
C803 source.n473 a_n1180_n5888# 0.355545f
C804 source.n474 a_n1180_n5888# 3.15511f
C805 source.n475 a_n1180_n5888# 0.015659f
C806 source.n476 a_n1180_n5888# 0.01658f
C807 source.n477 a_n1180_n5888# 0.037012f
C808 source.n478 a_n1180_n5888# 0.037012f
C809 source.n479 a_n1180_n5888# 0.01658f
C810 source.n480 a_n1180_n5888# 0.015659f
C811 source.n481 a_n1180_n5888# 0.029141f
C812 source.n482 a_n1180_n5888# 0.029141f
C813 source.n483 a_n1180_n5888# 0.015659f
C814 source.n484 a_n1180_n5888# 0.01658f
C815 source.n485 a_n1180_n5888# 0.037012f
C816 source.n486 a_n1180_n5888# 0.037012f
C817 source.n487 a_n1180_n5888# 0.01658f
C818 source.n488 a_n1180_n5888# 0.015659f
C819 source.n489 a_n1180_n5888# 0.029141f
C820 source.n490 a_n1180_n5888# 0.029141f
C821 source.n491 a_n1180_n5888# 0.015659f
C822 source.n492 a_n1180_n5888# 0.015659f
C823 source.n493 a_n1180_n5888# 0.01658f
C824 source.n494 a_n1180_n5888# 0.037012f
C825 source.n495 a_n1180_n5888# 0.037012f
C826 source.n496 a_n1180_n5888# 0.037012f
C827 source.n497 a_n1180_n5888# 0.01612f
C828 source.n498 a_n1180_n5888# 0.015659f
C829 source.n499 a_n1180_n5888# 0.029141f
C830 source.n500 a_n1180_n5888# 0.029141f
C831 source.n501 a_n1180_n5888# 0.015659f
C832 source.n502 a_n1180_n5888# 0.01658f
C833 source.n503 a_n1180_n5888# 0.037012f
C834 source.n504 a_n1180_n5888# 0.037012f
C835 source.n505 a_n1180_n5888# 0.01658f
C836 source.n506 a_n1180_n5888# 0.015659f
C837 source.n507 a_n1180_n5888# 0.029141f
C838 source.n508 a_n1180_n5888# 0.029141f
C839 source.n509 a_n1180_n5888# 0.015659f
C840 source.n510 a_n1180_n5888# 0.01658f
C841 source.n511 a_n1180_n5888# 0.037012f
C842 source.n512 a_n1180_n5888# 0.037012f
C843 source.n513 a_n1180_n5888# 0.01658f
C844 source.n514 a_n1180_n5888# 0.015659f
C845 source.n515 a_n1180_n5888# 0.029141f
C846 source.n516 a_n1180_n5888# 0.029141f
C847 source.n517 a_n1180_n5888# 0.015659f
C848 source.n518 a_n1180_n5888# 0.01658f
C849 source.n519 a_n1180_n5888# 0.037012f
C850 source.n520 a_n1180_n5888# 0.037012f
C851 source.n521 a_n1180_n5888# 0.01658f
C852 source.n522 a_n1180_n5888# 0.015659f
C853 source.n523 a_n1180_n5888# 0.029141f
C854 source.n524 a_n1180_n5888# 0.029141f
C855 source.n525 a_n1180_n5888# 0.015659f
C856 source.n526 a_n1180_n5888# 0.01658f
C857 source.n527 a_n1180_n5888# 0.037012f
C858 source.n528 a_n1180_n5888# 0.037012f
C859 source.n529 a_n1180_n5888# 0.01658f
C860 source.n530 a_n1180_n5888# 0.015659f
C861 source.n531 a_n1180_n5888# 0.029141f
C862 source.n532 a_n1180_n5888# 0.029141f
C863 source.n533 a_n1180_n5888# 0.015659f
C864 source.n534 a_n1180_n5888# 0.01658f
C865 source.n535 a_n1180_n5888# 0.037012f
C866 source.n536 a_n1180_n5888# 0.037012f
C867 source.n537 a_n1180_n5888# 0.037012f
C868 source.n538 a_n1180_n5888# 0.01658f
C869 source.n539 a_n1180_n5888# 0.015659f
C870 source.n540 a_n1180_n5888# 0.029141f
C871 source.n541 a_n1180_n5888# 0.029141f
C872 source.n542 a_n1180_n5888# 0.015659f
C873 source.n543 a_n1180_n5888# 0.01612f
C874 source.n544 a_n1180_n5888# 0.01612f
C875 source.n545 a_n1180_n5888# 0.037012f
C876 source.n546 a_n1180_n5888# 0.037012f
C877 source.n547 a_n1180_n5888# 0.01658f
C878 source.n548 a_n1180_n5888# 0.015659f
C879 source.n549 a_n1180_n5888# 0.029141f
C880 source.n550 a_n1180_n5888# 0.029141f
C881 source.n551 a_n1180_n5888# 0.015659f
C882 source.n552 a_n1180_n5888# 0.01658f
C883 source.n553 a_n1180_n5888# 0.037012f
C884 source.n554 a_n1180_n5888# 0.037012f
C885 source.n555 a_n1180_n5888# 0.01658f
C886 source.n556 a_n1180_n5888# 0.015659f
C887 source.n557 a_n1180_n5888# 0.029141f
C888 source.n558 a_n1180_n5888# 0.029141f
C889 source.n559 a_n1180_n5888# 0.015659f
C890 source.n560 a_n1180_n5888# 0.01658f
C891 source.n561 a_n1180_n5888# 0.037012f
C892 source.n562 a_n1180_n5888# 0.078735f
C893 source.n563 a_n1180_n5888# 0.01658f
C894 source.n564 a_n1180_n5888# 0.015659f
C895 source.n565 a_n1180_n5888# 0.064173f
C896 source.n566 a_n1180_n5888# 0.043812f
C897 source.n567 a_n1180_n5888# 0.27542f
C898 source.n568 a_n1180_n5888# 3.10384f
C899 drain_left.n0 a_n1180_n5888# 0.040356f
C900 drain_left.n1 a_n1180_n5888# 0.029273f
C901 drain_left.n2 a_n1180_n5888# 0.01573f
C902 drain_left.n3 a_n1180_n5888# 0.03718f
C903 drain_left.n4 a_n1180_n5888# 0.016655f
C904 drain_left.n5 a_n1180_n5888# 0.029273f
C905 drain_left.n6 a_n1180_n5888# 0.01573f
C906 drain_left.n7 a_n1180_n5888# 0.03718f
C907 drain_left.n8 a_n1180_n5888# 0.016655f
C908 drain_left.n9 a_n1180_n5888# 0.029273f
C909 drain_left.n10 a_n1180_n5888# 0.01573f
C910 drain_left.n11 a_n1180_n5888# 0.03718f
C911 drain_left.n12 a_n1180_n5888# 0.016655f
C912 drain_left.n13 a_n1180_n5888# 0.029273f
C913 drain_left.n14 a_n1180_n5888# 0.01573f
C914 drain_left.n15 a_n1180_n5888# 0.03718f
C915 drain_left.n16 a_n1180_n5888# 0.016655f
C916 drain_left.n17 a_n1180_n5888# 0.029273f
C917 drain_left.n18 a_n1180_n5888# 0.01573f
C918 drain_left.n19 a_n1180_n5888# 0.03718f
C919 drain_left.n20 a_n1180_n5888# 0.016655f
C920 drain_left.n21 a_n1180_n5888# 0.029273f
C921 drain_left.n22 a_n1180_n5888# 0.01573f
C922 drain_left.n23 a_n1180_n5888# 0.03718f
C923 drain_left.n24 a_n1180_n5888# 0.016655f
C924 drain_left.n25 a_n1180_n5888# 0.029273f
C925 drain_left.n26 a_n1180_n5888# 0.01573f
C926 drain_left.n27 a_n1180_n5888# 0.03718f
C927 drain_left.n28 a_n1180_n5888# 0.016655f
C928 drain_left.n29 a_n1180_n5888# 0.029273f
C929 drain_left.n30 a_n1180_n5888# 0.01573f
C930 drain_left.n31 a_n1180_n5888# 0.03718f
C931 drain_left.n32 a_n1180_n5888# 0.016655f
C932 drain_left.n33 a_n1180_n5888# 0.029273f
C933 drain_left.n34 a_n1180_n5888# 0.016193f
C934 drain_left.n35 a_n1180_n5888# 0.03718f
C935 drain_left.n36 a_n1180_n5888# 0.016655f
C936 drain_left.n37 a_n1180_n5888# 0.029273f
C937 drain_left.n38 a_n1180_n5888# 0.01573f
C938 drain_left.n39 a_n1180_n5888# 0.03718f
C939 drain_left.n40 a_n1180_n5888# 0.016655f
C940 drain_left.n41 a_n1180_n5888# 0.029273f
C941 drain_left.n42 a_n1180_n5888# 0.01573f
C942 drain_left.n43 a_n1180_n5888# 0.027885f
C943 drain_left.n44 a_n1180_n5888# 0.026283f
C944 drain_left.t1 a_n1180_n5888# 0.064844f
C945 drain_left.n45 a_n1180_n5888# 0.357155f
C946 drain_left.n46 a_n1180_n5888# 3.1694f
C947 drain_left.n47 a_n1180_n5888# 0.01573f
C948 drain_left.n48 a_n1180_n5888# 0.016655f
C949 drain_left.n49 a_n1180_n5888# 0.03718f
C950 drain_left.n50 a_n1180_n5888# 0.03718f
C951 drain_left.n51 a_n1180_n5888# 0.016655f
C952 drain_left.n52 a_n1180_n5888# 0.01573f
C953 drain_left.n53 a_n1180_n5888# 0.029273f
C954 drain_left.n54 a_n1180_n5888# 0.029273f
C955 drain_left.n55 a_n1180_n5888# 0.01573f
C956 drain_left.n56 a_n1180_n5888# 0.016655f
C957 drain_left.n57 a_n1180_n5888# 0.03718f
C958 drain_left.n58 a_n1180_n5888# 0.03718f
C959 drain_left.n59 a_n1180_n5888# 0.016655f
C960 drain_left.n60 a_n1180_n5888# 0.01573f
C961 drain_left.n61 a_n1180_n5888# 0.029273f
C962 drain_left.n62 a_n1180_n5888# 0.029273f
C963 drain_left.n63 a_n1180_n5888# 0.01573f
C964 drain_left.n64 a_n1180_n5888# 0.01573f
C965 drain_left.n65 a_n1180_n5888# 0.016655f
C966 drain_left.n66 a_n1180_n5888# 0.03718f
C967 drain_left.n67 a_n1180_n5888# 0.03718f
C968 drain_left.n68 a_n1180_n5888# 0.03718f
C969 drain_left.n69 a_n1180_n5888# 0.016193f
C970 drain_left.n70 a_n1180_n5888# 0.01573f
C971 drain_left.n71 a_n1180_n5888# 0.029273f
C972 drain_left.n72 a_n1180_n5888# 0.029273f
C973 drain_left.n73 a_n1180_n5888# 0.01573f
C974 drain_left.n74 a_n1180_n5888# 0.016655f
C975 drain_left.n75 a_n1180_n5888# 0.03718f
C976 drain_left.n76 a_n1180_n5888# 0.03718f
C977 drain_left.n77 a_n1180_n5888# 0.016655f
C978 drain_left.n78 a_n1180_n5888# 0.01573f
C979 drain_left.n79 a_n1180_n5888# 0.029273f
C980 drain_left.n80 a_n1180_n5888# 0.029273f
C981 drain_left.n81 a_n1180_n5888# 0.01573f
C982 drain_left.n82 a_n1180_n5888# 0.016655f
C983 drain_left.n83 a_n1180_n5888# 0.03718f
C984 drain_left.n84 a_n1180_n5888# 0.03718f
C985 drain_left.n85 a_n1180_n5888# 0.016655f
C986 drain_left.n86 a_n1180_n5888# 0.01573f
C987 drain_left.n87 a_n1180_n5888# 0.029273f
C988 drain_left.n88 a_n1180_n5888# 0.029273f
C989 drain_left.n89 a_n1180_n5888# 0.01573f
C990 drain_left.n90 a_n1180_n5888# 0.016655f
C991 drain_left.n91 a_n1180_n5888# 0.03718f
C992 drain_left.n92 a_n1180_n5888# 0.03718f
C993 drain_left.n93 a_n1180_n5888# 0.016655f
C994 drain_left.n94 a_n1180_n5888# 0.01573f
C995 drain_left.n95 a_n1180_n5888# 0.029273f
C996 drain_left.n96 a_n1180_n5888# 0.029273f
C997 drain_left.n97 a_n1180_n5888# 0.01573f
C998 drain_left.n98 a_n1180_n5888# 0.016655f
C999 drain_left.n99 a_n1180_n5888# 0.03718f
C1000 drain_left.n100 a_n1180_n5888# 0.03718f
C1001 drain_left.n101 a_n1180_n5888# 0.016655f
C1002 drain_left.n102 a_n1180_n5888# 0.01573f
C1003 drain_left.n103 a_n1180_n5888# 0.029273f
C1004 drain_left.n104 a_n1180_n5888# 0.029273f
C1005 drain_left.n105 a_n1180_n5888# 0.01573f
C1006 drain_left.n106 a_n1180_n5888# 0.016655f
C1007 drain_left.n107 a_n1180_n5888# 0.03718f
C1008 drain_left.n108 a_n1180_n5888# 0.03718f
C1009 drain_left.n109 a_n1180_n5888# 0.03718f
C1010 drain_left.n110 a_n1180_n5888# 0.016655f
C1011 drain_left.n111 a_n1180_n5888# 0.01573f
C1012 drain_left.n112 a_n1180_n5888# 0.029273f
C1013 drain_left.n113 a_n1180_n5888# 0.029273f
C1014 drain_left.n114 a_n1180_n5888# 0.01573f
C1015 drain_left.n115 a_n1180_n5888# 0.016193f
C1016 drain_left.n116 a_n1180_n5888# 0.016193f
C1017 drain_left.n117 a_n1180_n5888# 0.03718f
C1018 drain_left.n118 a_n1180_n5888# 0.03718f
C1019 drain_left.n119 a_n1180_n5888# 0.016655f
C1020 drain_left.n120 a_n1180_n5888# 0.01573f
C1021 drain_left.n121 a_n1180_n5888# 0.029273f
C1022 drain_left.n122 a_n1180_n5888# 0.029273f
C1023 drain_left.n123 a_n1180_n5888# 0.01573f
C1024 drain_left.n124 a_n1180_n5888# 0.016655f
C1025 drain_left.n125 a_n1180_n5888# 0.03718f
C1026 drain_left.n126 a_n1180_n5888# 0.03718f
C1027 drain_left.n127 a_n1180_n5888# 0.016655f
C1028 drain_left.n128 a_n1180_n5888# 0.01573f
C1029 drain_left.n129 a_n1180_n5888# 0.029273f
C1030 drain_left.n130 a_n1180_n5888# 0.029273f
C1031 drain_left.n131 a_n1180_n5888# 0.01573f
C1032 drain_left.n132 a_n1180_n5888# 0.016655f
C1033 drain_left.n133 a_n1180_n5888# 0.03718f
C1034 drain_left.n134 a_n1180_n5888# 0.079091f
C1035 drain_left.n135 a_n1180_n5888# 0.016655f
C1036 drain_left.n136 a_n1180_n5888# 0.01573f
C1037 drain_left.n137 a_n1180_n5888# 0.064464f
C1038 drain_left.n138 a_n1180_n5888# 0.064832f
C1039 drain_left.t5 a_n1180_n5888# 0.578309f
C1040 drain_left.t0 a_n1180_n5888# 0.578309f
C1041 drain_left.n139 a_n1180_n5888# 5.33013f
C1042 drain_left.n140 a_n1180_n5888# 2.59231f
C1043 drain_left.n141 a_n1180_n5888# 0.040356f
C1044 drain_left.n142 a_n1180_n5888# 0.029273f
C1045 drain_left.n143 a_n1180_n5888# 0.01573f
C1046 drain_left.n144 a_n1180_n5888# 0.03718f
C1047 drain_left.n145 a_n1180_n5888# 0.016655f
C1048 drain_left.n146 a_n1180_n5888# 0.029273f
C1049 drain_left.n147 a_n1180_n5888# 0.01573f
C1050 drain_left.n148 a_n1180_n5888# 0.03718f
C1051 drain_left.n149 a_n1180_n5888# 0.016655f
C1052 drain_left.n150 a_n1180_n5888# 0.029273f
C1053 drain_left.n151 a_n1180_n5888# 0.01573f
C1054 drain_left.n152 a_n1180_n5888# 0.03718f
C1055 drain_left.n153 a_n1180_n5888# 0.016655f
C1056 drain_left.n154 a_n1180_n5888# 0.029273f
C1057 drain_left.n155 a_n1180_n5888# 0.01573f
C1058 drain_left.n156 a_n1180_n5888# 0.03718f
C1059 drain_left.n157 a_n1180_n5888# 0.03718f
C1060 drain_left.n158 a_n1180_n5888# 0.016655f
C1061 drain_left.n159 a_n1180_n5888# 0.029273f
C1062 drain_left.n160 a_n1180_n5888# 0.01573f
C1063 drain_left.n161 a_n1180_n5888# 0.03718f
C1064 drain_left.n162 a_n1180_n5888# 0.016655f
C1065 drain_left.n163 a_n1180_n5888# 0.029273f
C1066 drain_left.n164 a_n1180_n5888# 0.01573f
C1067 drain_left.n165 a_n1180_n5888# 0.03718f
C1068 drain_left.n166 a_n1180_n5888# 0.016655f
C1069 drain_left.n167 a_n1180_n5888# 0.029273f
C1070 drain_left.n168 a_n1180_n5888# 0.01573f
C1071 drain_left.n169 a_n1180_n5888# 0.03718f
C1072 drain_left.n170 a_n1180_n5888# 0.016655f
C1073 drain_left.n171 a_n1180_n5888# 0.029273f
C1074 drain_left.n172 a_n1180_n5888# 0.01573f
C1075 drain_left.n173 a_n1180_n5888# 0.03718f
C1076 drain_left.n174 a_n1180_n5888# 0.016655f
C1077 drain_left.n175 a_n1180_n5888# 0.029273f
C1078 drain_left.n176 a_n1180_n5888# 0.016193f
C1079 drain_left.n177 a_n1180_n5888# 0.03718f
C1080 drain_left.n178 a_n1180_n5888# 0.01573f
C1081 drain_left.n179 a_n1180_n5888# 0.016655f
C1082 drain_left.n180 a_n1180_n5888# 0.029273f
C1083 drain_left.n181 a_n1180_n5888# 0.01573f
C1084 drain_left.n182 a_n1180_n5888# 0.03718f
C1085 drain_left.n183 a_n1180_n5888# 0.016655f
C1086 drain_left.n184 a_n1180_n5888# 0.029273f
C1087 drain_left.n185 a_n1180_n5888# 0.01573f
C1088 drain_left.n186 a_n1180_n5888# 0.027885f
C1089 drain_left.n187 a_n1180_n5888# 0.026283f
C1090 drain_left.t3 a_n1180_n5888# 0.064844f
C1091 drain_left.n188 a_n1180_n5888# 0.357155f
C1092 drain_left.n189 a_n1180_n5888# 3.1694f
C1093 drain_left.n190 a_n1180_n5888# 0.01573f
C1094 drain_left.n191 a_n1180_n5888# 0.016655f
C1095 drain_left.n192 a_n1180_n5888# 0.03718f
C1096 drain_left.n193 a_n1180_n5888# 0.03718f
C1097 drain_left.n194 a_n1180_n5888# 0.016655f
C1098 drain_left.n195 a_n1180_n5888# 0.01573f
C1099 drain_left.n196 a_n1180_n5888# 0.029273f
C1100 drain_left.n197 a_n1180_n5888# 0.029273f
C1101 drain_left.n198 a_n1180_n5888# 0.01573f
C1102 drain_left.n199 a_n1180_n5888# 0.016655f
C1103 drain_left.n200 a_n1180_n5888# 0.03718f
C1104 drain_left.n201 a_n1180_n5888# 0.03718f
C1105 drain_left.n202 a_n1180_n5888# 0.016655f
C1106 drain_left.n203 a_n1180_n5888# 0.01573f
C1107 drain_left.n204 a_n1180_n5888# 0.029273f
C1108 drain_left.n205 a_n1180_n5888# 0.029273f
C1109 drain_left.n206 a_n1180_n5888# 0.01573f
C1110 drain_left.n207 a_n1180_n5888# 0.016655f
C1111 drain_left.n208 a_n1180_n5888# 0.03718f
C1112 drain_left.n209 a_n1180_n5888# 0.03718f
C1113 drain_left.n210 a_n1180_n5888# 0.03718f
C1114 drain_left.n211 a_n1180_n5888# 0.016193f
C1115 drain_left.n212 a_n1180_n5888# 0.01573f
C1116 drain_left.n213 a_n1180_n5888# 0.029273f
C1117 drain_left.n214 a_n1180_n5888# 0.029273f
C1118 drain_left.n215 a_n1180_n5888# 0.01573f
C1119 drain_left.n216 a_n1180_n5888# 0.016655f
C1120 drain_left.n217 a_n1180_n5888# 0.03718f
C1121 drain_left.n218 a_n1180_n5888# 0.03718f
C1122 drain_left.n219 a_n1180_n5888# 0.016655f
C1123 drain_left.n220 a_n1180_n5888# 0.01573f
C1124 drain_left.n221 a_n1180_n5888# 0.029273f
C1125 drain_left.n222 a_n1180_n5888# 0.029273f
C1126 drain_left.n223 a_n1180_n5888# 0.01573f
C1127 drain_left.n224 a_n1180_n5888# 0.016655f
C1128 drain_left.n225 a_n1180_n5888# 0.03718f
C1129 drain_left.n226 a_n1180_n5888# 0.03718f
C1130 drain_left.n227 a_n1180_n5888# 0.016655f
C1131 drain_left.n228 a_n1180_n5888# 0.01573f
C1132 drain_left.n229 a_n1180_n5888# 0.029273f
C1133 drain_left.n230 a_n1180_n5888# 0.029273f
C1134 drain_left.n231 a_n1180_n5888# 0.01573f
C1135 drain_left.n232 a_n1180_n5888# 0.016655f
C1136 drain_left.n233 a_n1180_n5888# 0.03718f
C1137 drain_left.n234 a_n1180_n5888# 0.03718f
C1138 drain_left.n235 a_n1180_n5888# 0.016655f
C1139 drain_left.n236 a_n1180_n5888# 0.01573f
C1140 drain_left.n237 a_n1180_n5888# 0.029273f
C1141 drain_left.n238 a_n1180_n5888# 0.029273f
C1142 drain_left.n239 a_n1180_n5888# 0.01573f
C1143 drain_left.n240 a_n1180_n5888# 0.016655f
C1144 drain_left.n241 a_n1180_n5888# 0.03718f
C1145 drain_left.n242 a_n1180_n5888# 0.03718f
C1146 drain_left.n243 a_n1180_n5888# 0.016655f
C1147 drain_left.n244 a_n1180_n5888# 0.01573f
C1148 drain_left.n245 a_n1180_n5888# 0.029273f
C1149 drain_left.n246 a_n1180_n5888# 0.029273f
C1150 drain_left.n247 a_n1180_n5888# 0.01573f
C1151 drain_left.n248 a_n1180_n5888# 0.016655f
C1152 drain_left.n249 a_n1180_n5888# 0.03718f
C1153 drain_left.n250 a_n1180_n5888# 0.03718f
C1154 drain_left.n251 a_n1180_n5888# 0.016655f
C1155 drain_left.n252 a_n1180_n5888# 0.01573f
C1156 drain_left.n253 a_n1180_n5888# 0.029273f
C1157 drain_left.n254 a_n1180_n5888# 0.029273f
C1158 drain_left.n255 a_n1180_n5888# 0.01573f
C1159 drain_left.n256 a_n1180_n5888# 0.016193f
C1160 drain_left.n257 a_n1180_n5888# 0.016193f
C1161 drain_left.n258 a_n1180_n5888# 0.03718f
C1162 drain_left.n259 a_n1180_n5888# 0.03718f
C1163 drain_left.n260 a_n1180_n5888# 0.016655f
C1164 drain_left.n261 a_n1180_n5888# 0.01573f
C1165 drain_left.n262 a_n1180_n5888# 0.029273f
C1166 drain_left.n263 a_n1180_n5888# 0.029273f
C1167 drain_left.n264 a_n1180_n5888# 0.01573f
C1168 drain_left.n265 a_n1180_n5888# 0.016655f
C1169 drain_left.n266 a_n1180_n5888# 0.03718f
C1170 drain_left.n267 a_n1180_n5888# 0.03718f
C1171 drain_left.n268 a_n1180_n5888# 0.016655f
C1172 drain_left.n269 a_n1180_n5888# 0.01573f
C1173 drain_left.n270 a_n1180_n5888# 0.029273f
C1174 drain_left.n271 a_n1180_n5888# 0.029273f
C1175 drain_left.n272 a_n1180_n5888# 0.01573f
C1176 drain_left.n273 a_n1180_n5888# 0.016655f
C1177 drain_left.n274 a_n1180_n5888# 0.03718f
C1178 drain_left.n275 a_n1180_n5888# 0.079091f
C1179 drain_left.n276 a_n1180_n5888# 0.016655f
C1180 drain_left.n277 a_n1180_n5888# 0.01573f
C1181 drain_left.n278 a_n1180_n5888# 0.064464f
C1182 drain_left.n279 a_n1180_n5888# 0.065313f
C1183 drain_left.t2 a_n1180_n5888# 0.578309f
C1184 drain_left.t4 a_n1180_n5888# 0.578309f
C1185 drain_left.n280 a_n1180_n5888# 5.32973f
C1186 drain_left.n281 a_n1180_n5888# 0.684041f
C1187 plus.t1 a_n1180_n5888# 1.08164f
C1188 plus.n0 a_n1180_n5888# 0.413001f
C1189 plus.t0 a_n1180_n5888# 1.07423f
C1190 plus.n1 a_n1180_n5888# 0.394028f
C1191 plus.t2 a_n1180_n5888# 1.08164f
C1192 plus.n2 a_n1180_n5888# 0.412911f
C1193 plus.n3 a_n1180_n5888# 1.16485f
C1194 plus.t5 a_n1180_n5888# 1.08164f
C1195 plus.n4 a_n1180_n5888# 0.413001f
C1196 plus.t3 a_n1180_n5888# 1.08164f
C1197 plus.t4 a_n1180_n5888# 1.07423f
C1198 plus.n5 a_n1180_n5888# 0.394028f
C1199 plus.n6 a_n1180_n5888# 0.412911f
C1200 plus.n7 a_n1180_n5888# 2.22496f
.ends

