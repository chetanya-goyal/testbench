* NGSPICE file created from diffpair596.ext - technology: sky130A

.subckt diffpair596 minus drain_right drain_left source plus
X0 drain_left.t13 plus.t0 source.t16 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X1 drain_left.t12 plus.t1 source.t25 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X2 source.t2 minus.t0 drain_right.t13 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X3 drain_right.t12 minus.t1 source.t6 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X4 a_n1724_n4888# a_n1724_n4888# a_n1724_n4888# a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=62.4 ps=326.24 w=20 l=0.3
X5 drain_right.t11 minus.t2 source.t8 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X6 drain_right.t10 minus.t3 source.t1 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X7 drain_left.t11 plus.t2 source.t17 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X8 drain_right.t9 minus.t4 source.t0 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X9 drain_left.t10 plus.t3 source.t20 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X10 drain_left.t9 plus.t4 source.t22 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=3.3 ps=20.33 w=20 l=0.3
X11 a_n1724_n4888# a_n1724_n4888# a_n1724_n4888# a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X12 drain_left.t8 plus.t5 source.t26 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X13 source.t14 plus.t6 drain_left.t7 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X14 drain_right.t8 minus.t5 source.t11 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X15 drain_right.t7 minus.t6 source.t7 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X16 source.t10 minus.t7 drain_right.t6 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X17 drain_right.t5 minus.t8 source.t4 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X18 source.t18 plus.t7 drain_left.t6 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X19 source.t21 plus.t8 drain_left.t5 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X20 drain_left.t4 plus.t9 source.t24 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X21 source.t19 plus.t10 drain_left.t3 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X22 source.t27 plus.t11 drain_left.t2 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X23 source.t12 minus.t9 drain_right.t4 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X24 source.t13 minus.t10 drain_right.t3 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X25 a_n1724_n4888# a_n1724_n4888# a_n1724_n4888# a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X26 drain_right.t2 minus.t11 source.t3 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X27 a_n1724_n4888# a_n1724_n4888# a_n1724_n4888# a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=7.8 pd=40.78 as=0 ps=0 w=20 l=0.3
X28 source.t9 minus.t12 drain_right.t1 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X29 source.t5 minus.t13 drain_right.t0 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
X30 drain_left.t1 plus.t12 source.t15 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=7.8 ps=40.78 w=20 l=0.3
X31 source.t23 plus.t13 drain_left.t0 a_n1724_n4888# sky130_fd_pr__nfet_01v8 ad=3.3 pd=20.33 as=3.3 ps=20.33 w=20 l=0.3
R0 plus.n3 plus.t2 1768.06
R1 plus.n15 plus.t12 1768.06
R2 plus.n20 plus.t0 1768.06
R3 plus.n32 plus.t4 1768.06
R4 plus.n1 plus.t13 1711.1
R5 plus.n4 plus.t6 1711.1
R6 plus.n6 plus.t9 1711.1
R7 plus.n12 plus.t5 1711.1
R8 plus.n14 plus.t7 1711.1
R9 plus.n18 plus.t10 1711.1
R10 plus.n21 plus.t8 1711.1
R11 plus.n23 plus.t1 1711.1
R12 plus.n29 plus.t3 1711.1
R13 plus.n31 plus.t11 1711.1
R14 plus.n3 plus.n2 161.489
R15 plus.n20 plus.n19 161.489
R16 plus.n5 plus.n2 161.3
R17 plus.n8 plus.n7 161.3
R18 plus.n9 plus.n1 161.3
R19 plus.n11 plus.n10 161.3
R20 plus.n13 plus.n0 161.3
R21 plus.n16 plus.n15 161.3
R22 plus.n22 plus.n19 161.3
R23 plus.n25 plus.n24 161.3
R24 plus.n26 plus.n18 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n17 161.3
R27 plus.n33 plus.n32 161.3
R28 plus.n7 plus.n1 73.0308
R29 plus.n11 plus.n1 73.0308
R30 plus.n28 plus.n18 73.0308
R31 plus.n24 plus.n18 73.0308
R32 plus.n6 plus.n5 54.0429
R33 plus.n13 plus.n12 54.0429
R34 plus.n30 plus.n29 54.0429
R35 plus.n23 plus.n22 54.0429
R36 plus.n5 plus.n4 37.9763
R37 plus.n14 plus.n13 37.9763
R38 plus.n31 plus.n30 37.9763
R39 plus.n22 plus.n21 37.9763
R40 plus.n4 plus.n3 35.055
R41 plus.n15 plus.n14 35.055
R42 plus.n32 plus.n31 35.055
R43 plus.n21 plus.n20 35.055
R44 plus plus.n33 32.5994
R45 plus.n7 plus.n6 18.9884
R46 plus.n12 plus.n11 18.9884
R47 plus.n29 plus.n28 18.9884
R48 plus.n24 plus.n23 18.9884
R49 plus plus.n16 15.2107
R50 plus.n8 plus.n2 0.189894
R51 plus.n9 plus.n8 0.189894
R52 plus.n10 plus.n9 0.189894
R53 plus.n10 plus.n0 0.189894
R54 plus.n16 plus.n0 0.189894
R55 plus.n33 plus.n17 0.189894
R56 plus.n27 plus.n17 0.189894
R57 plus.n27 plus.n26 0.189894
R58 plus.n26 plus.n25 0.189894
R59 plus.n25 plus.n19 0.189894
R60 source.n0 source.t15 44.1297
R61 source.n7 source.t4 44.1296
R62 source.n27 source.t11 44.1295
R63 source.n20 source.t16 44.1295
R64 source.n2 source.n1 43.1397
R65 source.n4 source.n3 43.1397
R66 source.n6 source.n5 43.1397
R67 source.n9 source.n8 43.1397
R68 source.n11 source.n10 43.1397
R69 source.n13 source.n12 43.1397
R70 source.n26 source.n25 43.1396
R71 source.n24 source.n23 43.1396
R72 source.n22 source.n21 43.1396
R73 source.n19 source.n18 43.1396
R74 source.n17 source.n16 43.1396
R75 source.n15 source.n14 43.1396
R76 source.n15 source.n13 28.4345
R77 source.n28 source.n0 22.357
R78 source.n28 source.n27 5.53498
R79 source.n25 source.t7 0.9905
R80 source.n25 source.t5 0.9905
R81 source.n23 source.t8 0.9905
R82 source.n23 source.t12 0.9905
R83 source.n21 source.t1 0.9905
R84 source.n21 source.t13 0.9905
R85 source.n18 source.t25 0.9905
R86 source.n18 source.t21 0.9905
R87 source.n16 source.t20 0.9905
R88 source.n16 source.t19 0.9905
R89 source.n14 source.t22 0.9905
R90 source.n14 source.t27 0.9905
R91 source.n1 source.t26 0.9905
R92 source.n1 source.t18 0.9905
R93 source.n3 source.t24 0.9905
R94 source.n3 source.t23 0.9905
R95 source.n5 source.t17 0.9905
R96 source.n5 source.t14 0.9905
R97 source.n8 source.t6 0.9905
R98 source.n8 source.t9 0.9905
R99 source.n10 source.t3 0.9905
R100 source.n10 source.t10 0.9905
R101 source.n12 source.t0 0.9905
R102 source.n12 source.t2 0.9905
R103 source.n7 source.n6 0.741879
R104 source.n22 source.n20 0.741879
R105 source.n13 source.n11 0.543603
R106 source.n11 source.n9 0.543603
R107 source.n9 source.n7 0.543603
R108 source.n6 source.n4 0.543603
R109 source.n4 source.n2 0.543603
R110 source.n2 source.n0 0.543603
R111 source.n17 source.n15 0.543603
R112 source.n19 source.n17 0.543603
R113 source.n20 source.n19 0.543603
R114 source.n24 source.n22 0.543603
R115 source.n26 source.n24 0.543603
R116 source.n27 source.n26 0.543603
R117 source source.n28 0.188
R118 drain_left.n7 drain_left.t11 61.3515
R119 drain_left.n1 drain_left.t9 61.3514
R120 drain_left.n4 drain_left.n2 60.3615
R121 drain_left.n11 drain_left.n10 59.8185
R122 drain_left.n9 drain_left.n8 59.8185
R123 drain_left.n7 drain_left.n6 59.8185
R124 drain_left.n4 drain_left.n3 59.8184
R125 drain_left.n1 drain_left.n0 59.8184
R126 drain_left drain_left.n5 36.5505
R127 drain_left drain_left.n11 6.19632
R128 drain_left.n2 drain_left.t5 0.9905
R129 drain_left.n2 drain_left.t13 0.9905
R130 drain_left.n3 drain_left.t3 0.9905
R131 drain_left.n3 drain_left.t12 0.9905
R132 drain_left.n0 drain_left.t2 0.9905
R133 drain_left.n0 drain_left.t10 0.9905
R134 drain_left.n10 drain_left.t6 0.9905
R135 drain_left.n10 drain_left.t1 0.9905
R136 drain_left.n8 drain_left.t0 0.9905
R137 drain_left.n8 drain_left.t8 0.9905
R138 drain_left.n6 drain_left.t7 0.9905
R139 drain_left.n6 drain_left.t4 0.9905
R140 drain_left.n9 drain_left.n7 0.543603
R141 drain_left.n11 drain_left.n9 0.543603
R142 drain_left.n5 drain_left.n1 0.352482
R143 drain_left.n5 drain_left.n4 0.0809298
R144 minus.n15 minus.t4 1768.06
R145 minus.n3 minus.t8 1768.06
R146 minus.n32 minus.t5 1768.06
R147 minus.n20 minus.t3 1768.06
R148 minus.n1 minus.t7 1711.1
R149 minus.n14 minus.t0 1711.1
R150 minus.n12 minus.t11 1711.1
R151 minus.n6 minus.t1 1711.1
R152 minus.n4 minus.t12 1711.1
R153 minus.n18 minus.t9 1711.1
R154 minus.n31 minus.t13 1711.1
R155 minus.n29 minus.t6 1711.1
R156 minus.n23 minus.t2 1711.1
R157 minus.n21 minus.t10 1711.1
R158 minus.n3 minus.n2 161.489
R159 minus.n20 minus.n19 161.489
R160 minus.n16 minus.n15 161.3
R161 minus.n13 minus.n0 161.3
R162 minus.n11 minus.n10 161.3
R163 minus.n9 minus.n1 161.3
R164 minus.n8 minus.n7 161.3
R165 minus.n5 minus.n2 161.3
R166 minus.n33 minus.n32 161.3
R167 minus.n30 minus.n17 161.3
R168 minus.n28 minus.n27 161.3
R169 minus.n26 minus.n18 161.3
R170 minus.n25 minus.n24 161.3
R171 minus.n22 minus.n19 161.3
R172 minus.n11 minus.n1 73.0308
R173 minus.n7 minus.n1 73.0308
R174 minus.n24 minus.n18 73.0308
R175 minus.n28 minus.n18 73.0308
R176 minus.n13 minus.n12 54.0429
R177 minus.n6 minus.n5 54.0429
R178 minus.n23 minus.n22 54.0429
R179 minus.n30 minus.n29 54.0429
R180 minus.n34 minus.n16 41.7486
R181 minus.n14 minus.n13 37.9763
R182 minus.n5 minus.n4 37.9763
R183 minus.n22 minus.n21 37.9763
R184 minus.n31 minus.n30 37.9763
R185 minus.n15 minus.n14 35.055
R186 minus.n4 minus.n3 35.055
R187 minus.n21 minus.n20 35.055
R188 minus.n32 minus.n31 35.055
R189 minus.n12 minus.n11 18.9884
R190 minus.n7 minus.n6 18.9884
R191 minus.n24 minus.n23 18.9884
R192 minus.n29 minus.n28 18.9884
R193 minus.n34 minus.n33 6.53648
R194 minus.n16 minus.n0 0.189894
R195 minus.n10 minus.n0 0.189894
R196 minus.n10 minus.n9 0.189894
R197 minus.n9 minus.n8 0.189894
R198 minus.n8 minus.n2 0.189894
R199 minus.n25 minus.n19 0.189894
R200 minus.n26 minus.n25 0.189894
R201 minus.n27 minus.n26 0.189894
R202 minus.n27 minus.n17 0.189894
R203 minus.n33 minus.n17 0.189894
R204 minus minus.n34 0.188
R205 drain_right.n1 drain_right.t10 61.3514
R206 drain_right.n11 drain_right.t9 60.8084
R207 drain_right.n8 drain_right.n6 60.3616
R208 drain_right.n4 drain_right.n2 60.3615
R209 drain_right.n8 drain_right.n7 59.8185
R210 drain_right.n10 drain_right.n9 59.8185
R211 drain_right.n4 drain_right.n3 59.8184
R212 drain_right.n1 drain_right.n0 59.8184
R213 drain_right drain_right.n5 35.9973
R214 drain_right drain_right.n11 5.92477
R215 drain_right.n2 drain_right.t0 0.9905
R216 drain_right.n2 drain_right.t8 0.9905
R217 drain_right.n3 drain_right.t4 0.9905
R218 drain_right.n3 drain_right.t7 0.9905
R219 drain_right.n0 drain_right.t3 0.9905
R220 drain_right.n0 drain_right.t11 0.9905
R221 drain_right.n6 drain_right.t1 0.9905
R222 drain_right.n6 drain_right.t5 0.9905
R223 drain_right.n7 drain_right.t6 0.9905
R224 drain_right.n7 drain_right.t12 0.9905
R225 drain_right.n9 drain_right.t13 0.9905
R226 drain_right.n9 drain_right.t2 0.9905
R227 drain_right.n11 drain_right.n10 0.543603
R228 drain_right.n10 drain_right.n8 0.543603
R229 drain_right.n5 drain_right.n1 0.352482
R230 drain_right.n5 drain_right.n4 0.0809298
C0 plus minus 6.78065f
C1 source plus 7.80588f
C2 drain_left plus 8.63026f
C3 drain_right minus 8.4683f
C4 source drain_right 44.909f
C5 drain_left drain_right 0.886973f
C6 source minus 7.79075f
C7 drain_left minus 0.171678f
C8 source drain_left 44.926003f
C9 drain_right plus 0.324825f
C10 drain_right a_n1724_n4888# 9.77127f
C11 drain_left a_n1724_n4888# 10.044279f
C12 source a_n1724_n4888# 8.954455f
C13 minus a_n1724_n4888# 7.243491f
C14 plus a_n1724_n4888# 9.757781f
C15 drain_right.t10 a_n1724_n4888# 5.73059f
C16 drain_right.t3 a_n1724_n4888# 0.489794f
C17 drain_right.t11 a_n1724_n4888# 0.489794f
C18 drain_right.n0 a_n1724_n4888# 4.47781f
C19 drain_right.n1 a_n1724_n4888# 0.764194f
C20 drain_right.t0 a_n1724_n4888# 0.489794f
C21 drain_right.t8 a_n1724_n4888# 0.489794f
C22 drain_right.n2 a_n1724_n4888# 4.48125f
C23 drain_right.t4 a_n1724_n4888# 0.489794f
C24 drain_right.t7 a_n1724_n4888# 0.489794f
C25 drain_right.n3 a_n1724_n4888# 4.47781f
C26 drain_right.n4 a_n1724_n4888# 0.711739f
C27 drain_right.n5 a_n1724_n4888# 2.01855f
C28 drain_right.t1 a_n1724_n4888# 0.489794f
C29 drain_right.t5 a_n1724_n4888# 0.489794f
C30 drain_right.n6 a_n1724_n4888# 4.48124f
C31 drain_right.t6 a_n1724_n4888# 0.489794f
C32 drain_right.t12 a_n1724_n4888# 0.489794f
C33 drain_right.n7 a_n1724_n4888# 4.4778f
C34 drain_right.n8 a_n1724_n4888# 0.749021f
C35 drain_right.t13 a_n1724_n4888# 0.489794f
C36 drain_right.t2 a_n1724_n4888# 0.489794f
C37 drain_right.n9 a_n1724_n4888# 4.4778f
C38 drain_right.n10 a_n1724_n4888# 0.36999f
C39 drain_right.t9 a_n1724_n4888# 5.72694f
C40 drain_right.n11 a_n1724_n4888# 0.673444f
C41 minus.n0 a_n1724_n4888# 0.051686f
C42 minus.t4 a_n1724_n4888# 0.884091f
C43 minus.t0 a_n1724_n4888# 0.873442f
C44 minus.t11 a_n1724_n4888# 0.873442f
C45 minus.t7 a_n1724_n4888# 0.873442f
C46 minus.n1 a_n1724_n4888# 0.341609f
C47 minus.n2 a_n1724_n4888# 0.121773f
C48 minus.t1 a_n1724_n4888# 0.873442f
C49 minus.t12 a_n1724_n4888# 0.873442f
C50 minus.t8 a_n1724_n4888# 0.884091f
C51 minus.n3 a_n1724_n4888# 0.34124f
C52 minus.n4 a_n1724_n4888# 0.324463f
C53 minus.n5 a_n1724_n4888# 0.021289f
C54 minus.n6 a_n1724_n4888# 0.324463f
C55 minus.n7 a_n1724_n4888# 0.021289f
C56 minus.n8 a_n1724_n4888# 0.051686f
C57 minus.n9 a_n1724_n4888# 0.051686f
C58 minus.n10 a_n1724_n4888# 0.051686f
C59 minus.n11 a_n1724_n4888# 0.021289f
C60 minus.n12 a_n1724_n4888# 0.324463f
C61 minus.n13 a_n1724_n4888# 0.021289f
C62 minus.n14 a_n1724_n4888# 0.324463f
C63 minus.n15 a_n1724_n4888# 0.341158f
C64 minus.n16 a_n1724_n4888# 2.2701f
C65 minus.n17 a_n1724_n4888# 0.051686f
C66 minus.t13 a_n1724_n4888# 0.873442f
C67 minus.t6 a_n1724_n4888# 0.873442f
C68 minus.t9 a_n1724_n4888# 0.873442f
C69 minus.n18 a_n1724_n4888# 0.341609f
C70 minus.n19 a_n1724_n4888# 0.121773f
C71 minus.t2 a_n1724_n4888# 0.873442f
C72 minus.t10 a_n1724_n4888# 0.873442f
C73 minus.t3 a_n1724_n4888# 0.884091f
C74 minus.n20 a_n1724_n4888# 0.34124f
C75 minus.n21 a_n1724_n4888# 0.324463f
C76 minus.n22 a_n1724_n4888# 0.021289f
C77 minus.n23 a_n1724_n4888# 0.324463f
C78 minus.n24 a_n1724_n4888# 0.021289f
C79 minus.n25 a_n1724_n4888# 0.051686f
C80 minus.n26 a_n1724_n4888# 0.051686f
C81 minus.n27 a_n1724_n4888# 0.051686f
C82 minus.n28 a_n1724_n4888# 0.021289f
C83 minus.n29 a_n1724_n4888# 0.324463f
C84 minus.n30 a_n1724_n4888# 0.021289f
C85 minus.n31 a_n1724_n4888# 0.324463f
C86 minus.t5 a_n1724_n4888# 0.884091f
C87 minus.n32 a_n1724_n4888# 0.341158f
C88 minus.n33 a_n1724_n4888# 0.342347f
C89 minus.n34 a_n1724_n4888# 2.71176f
C90 drain_left.t9 a_n1724_n4888# 5.72832f
C91 drain_left.t2 a_n1724_n4888# 0.4896f
C92 drain_left.t10 a_n1724_n4888# 0.4896f
C93 drain_left.n0 a_n1724_n4888# 4.47603f
C94 drain_left.n1 a_n1724_n4888# 0.763891f
C95 drain_left.t5 a_n1724_n4888# 0.4896f
C96 drain_left.t13 a_n1724_n4888# 0.4896f
C97 drain_left.n2 a_n1724_n4888# 4.47947f
C98 drain_left.t3 a_n1724_n4888# 0.4896f
C99 drain_left.t12 a_n1724_n4888# 0.4896f
C100 drain_left.n3 a_n1724_n4888# 4.47603f
C101 drain_left.n4 a_n1724_n4888# 0.711457f
C102 drain_left.n5 a_n1724_n4888# 2.08234f
C103 drain_left.t11 a_n1724_n4888# 5.72834f
C104 drain_left.t7 a_n1724_n4888# 0.4896f
C105 drain_left.t4 a_n1724_n4888# 0.4896f
C106 drain_left.n6 a_n1724_n4888# 4.47603f
C107 drain_left.n7 a_n1724_n4888# 0.780913f
C108 drain_left.t0 a_n1724_n4888# 0.4896f
C109 drain_left.t8 a_n1724_n4888# 0.4896f
C110 drain_left.n8 a_n1724_n4888# 4.47603f
C111 drain_left.n9 a_n1724_n4888# 0.369843f
C112 drain_left.t6 a_n1724_n4888# 0.4896f
C113 drain_left.t1 a_n1724_n4888# 0.4896f
C114 drain_left.n10 a_n1724_n4888# 4.47603f
C115 drain_left.n11 a_n1724_n4888# 0.627695f
C116 source.t15 a_n1724_n4888# 5.6841f
C117 source.n0 a_n1724_n4888# 2.41764f
C118 source.t26 a_n1724_n4888# 0.497367f
C119 source.t18 a_n1724_n4888# 0.497367f
C120 source.n1 a_n1724_n4888# 4.44667f
C121 source.n2 a_n1724_n4888# 0.433295f
C122 source.t24 a_n1724_n4888# 0.497367f
C123 source.t23 a_n1724_n4888# 0.497367f
C124 source.n3 a_n1724_n4888# 4.44667f
C125 source.n4 a_n1724_n4888# 0.433295f
C126 source.t17 a_n1724_n4888# 0.497367f
C127 source.t14 a_n1724_n4888# 0.497367f
C128 source.n5 a_n1724_n4888# 4.44667f
C129 source.n6 a_n1724_n4888# 0.453401f
C130 source.t4 a_n1724_n4888# 5.68411f
C131 source.n7 a_n1724_n4888# 0.572418f
C132 source.t6 a_n1724_n4888# 0.497367f
C133 source.t9 a_n1724_n4888# 0.497367f
C134 source.n8 a_n1724_n4888# 4.44667f
C135 source.n9 a_n1724_n4888# 0.433295f
C136 source.t3 a_n1724_n4888# 0.497367f
C137 source.t10 a_n1724_n4888# 0.497367f
C138 source.n10 a_n1724_n4888# 4.44667f
C139 source.n11 a_n1724_n4888# 0.433295f
C140 source.t0 a_n1724_n4888# 0.497367f
C141 source.t2 a_n1724_n4888# 0.497367f
C142 source.n12 a_n1724_n4888# 4.44667f
C143 source.n13 a_n1724_n4888# 2.91137f
C144 source.t22 a_n1724_n4888# 0.497367f
C145 source.t27 a_n1724_n4888# 0.497367f
C146 source.n14 a_n1724_n4888# 4.44668f
C147 source.n15 a_n1724_n4888# 2.91136f
C148 source.t20 a_n1724_n4888# 0.497367f
C149 source.t19 a_n1724_n4888# 0.497367f
C150 source.n16 a_n1724_n4888# 4.44668f
C151 source.n17 a_n1724_n4888# 0.433286f
C152 source.t25 a_n1724_n4888# 0.497367f
C153 source.t21 a_n1724_n4888# 0.497367f
C154 source.n18 a_n1724_n4888# 4.44668f
C155 source.n19 a_n1724_n4888# 0.433286f
C156 source.t16 a_n1724_n4888# 5.68408f
C157 source.n20 a_n1724_n4888# 0.57245f
C158 source.t1 a_n1724_n4888# 0.497367f
C159 source.t13 a_n1724_n4888# 0.497367f
C160 source.n21 a_n1724_n4888# 4.44668f
C161 source.n22 a_n1724_n4888# 0.453392f
C162 source.t8 a_n1724_n4888# 0.497367f
C163 source.t12 a_n1724_n4888# 0.497367f
C164 source.n23 a_n1724_n4888# 4.44668f
C165 source.n24 a_n1724_n4888# 0.433286f
C166 source.t7 a_n1724_n4888# 0.497367f
C167 source.t5 a_n1724_n4888# 0.497367f
C168 source.n25 a_n1724_n4888# 4.44668f
C169 source.n26 a_n1724_n4888# 0.433286f
C170 source.t11 a_n1724_n4888# 5.68408f
C171 source.n27 a_n1724_n4888# 0.72256f
C172 source.n28 a_n1724_n4888# 2.83286f
C173 plus.n0 a_n1724_n4888# 0.052146f
C174 plus.t7 a_n1724_n4888# 0.881211f
C175 plus.t5 a_n1724_n4888# 0.881211f
C176 plus.t13 a_n1724_n4888# 0.881211f
C177 plus.n1 a_n1724_n4888# 0.344647f
C178 plus.n2 a_n1724_n4888# 0.122856f
C179 plus.t9 a_n1724_n4888# 0.881211f
C180 plus.t6 a_n1724_n4888# 0.881211f
C181 plus.t2 a_n1724_n4888# 0.891954f
C182 plus.n3 a_n1724_n4888# 0.344275f
C183 plus.n4 a_n1724_n4888# 0.327349f
C184 plus.n5 a_n1724_n4888# 0.021478f
C185 plus.n6 a_n1724_n4888# 0.327349f
C186 plus.n7 a_n1724_n4888# 0.021478f
C187 plus.n8 a_n1724_n4888# 0.052146f
C188 plus.n9 a_n1724_n4888# 0.052146f
C189 plus.n10 a_n1724_n4888# 0.052146f
C190 plus.n11 a_n1724_n4888# 0.021478f
C191 plus.n12 a_n1724_n4888# 0.327349f
C192 plus.n13 a_n1724_n4888# 0.021478f
C193 plus.n14 a_n1724_n4888# 0.327349f
C194 plus.t12 a_n1724_n4888# 0.891954f
C195 plus.n15 a_n1724_n4888# 0.344192f
C196 plus.n16 a_n1724_n4888# 0.796177f
C197 plus.n17 a_n1724_n4888# 0.052146f
C198 plus.t4 a_n1724_n4888# 0.891954f
C199 plus.t11 a_n1724_n4888# 0.881211f
C200 plus.t3 a_n1724_n4888# 0.881211f
C201 plus.t10 a_n1724_n4888# 0.881211f
C202 plus.n18 a_n1724_n4888# 0.344647f
C203 plus.n19 a_n1724_n4888# 0.122856f
C204 plus.t1 a_n1724_n4888# 0.881211f
C205 plus.t8 a_n1724_n4888# 0.881211f
C206 plus.t0 a_n1724_n4888# 0.891954f
C207 plus.n20 a_n1724_n4888# 0.344275f
C208 plus.n21 a_n1724_n4888# 0.327349f
C209 plus.n22 a_n1724_n4888# 0.021478f
C210 plus.n23 a_n1724_n4888# 0.327349f
C211 plus.n24 a_n1724_n4888# 0.021478f
C212 plus.n25 a_n1724_n4888# 0.052146f
C213 plus.n26 a_n1724_n4888# 0.052146f
C214 plus.n27 a_n1724_n4888# 0.052146f
C215 plus.n28 a_n1724_n4888# 0.021478f
C216 plus.n29 a_n1724_n4888# 0.327349f
C217 plus.n30 a_n1724_n4888# 0.021478f
C218 plus.n31 a_n1724_n4888# 0.327349f
C219 plus.n32 a_n1724_n4888# 0.344192f
C220 plus.n33 a_n1724_n4888# 1.80919f
.ends

