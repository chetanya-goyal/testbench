* NGSPICE file created from diffpair267.ext - technology: sky130A

.subckt diffpair267 minus drain_right drain_left source plus
X0 drain_left.t15 plus.t0 source.t16 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X1 drain_left.t14 plus.t1 source.t31 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X2 drain_left.t13 plus.t2 source.t22 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X3 source.t8 minus.t0 drain_right.t15 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X4 drain_left.t12 plus.t3 source.t26 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X5 source.t2 minus.t1 drain_right.t14 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X6 a_n1760_n2088# a_n1760_n2088# a_n1760_n2088# a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.25
X7 a_n1760_n2088# a_n1760_n2088# a_n1760_n2088# a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X8 source.t25 plus.t4 drain_left.t11 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X9 drain_right.t13 minus.t2 source.t1 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X10 source.t3 minus.t3 drain_right.t12 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X11 drain_right.t11 minus.t4 source.t6 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X12 drain_left.t10 plus.t5 source.t24 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X13 source.t9 minus.t5 drain_right.t10 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X14 source.t11 minus.t6 drain_right.t9 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X15 source.t29 plus.t6 drain_left.t9 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X16 source.t0 minus.t7 drain_right.t8 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X17 source.t28 plus.t7 drain_left.t8 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X18 source.t21 plus.t8 drain_left.t7 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X19 source.t27 plus.t9 drain_left.t6 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X20 source.t20 plus.t10 drain_left.t5 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X21 a_n1760_n2088# a_n1760_n2088# a_n1760_n2088# a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X22 drain_left.t4 plus.t11 source.t18 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X23 drain_right.t7 minus.t8 source.t13 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X24 a_n1760_n2088# a_n1760_n2088# a_n1760_n2088# a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.25
X25 drain_right.t6 minus.t9 source.t4 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X26 source.t12 minus.t10 drain_right.t5 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
X27 drain_right.t4 minus.t11 source.t15 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.25
X28 source.t17 plus.t12 drain_left.t3 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X29 drain_right.t3 minus.t12 source.t5 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X30 drain_left.t2 plus.t13 source.t19 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X31 drain_right.t2 minus.t13 source.t14 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X32 drain_right.t1 minus.t14 source.t7 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X33 source.t10 minus.t15 drain_right.t0 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X34 drain_left.t1 plus.t14 source.t30 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.25
X35 source.t23 plus.t15 drain_left.t0 a_n1760_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.25
R0 plus.n4 plus.t4 744.617
R1 plus.n19 plus.t3 744.617
R2 plus.n25 plus.t11 744.617
R3 plus.n40 plus.t15 744.617
R4 plus.n5 plus.t1 703.721
R5 plus.n3 plus.t10 703.721
R6 plus.n10 plus.t0 703.721
R7 plus.n1 plus.t9 703.721
R8 plus.n16 plus.t14 703.721
R9 plus.n18 plus.t8 703.721
R10 plus.n26 plus.t6 703.721
R11 plus.n24 plus.t2 703.721
R12 plus.n31 plus.t12 703.721
R13 plus.n22 plus.t13 703.721
R14 plus.n37 plus.t7 703.721
R15 plus.n39 plus.t5 703.721
R16 plus.n7 plus.n4 161.489
R17 plus.n28 plus.n25 161.489
R18 plus.n7 plus.n6 161.3
R19 plus.n9 plus.n8 161.3
R20 plus.n11 plus.n2 161.3
R21 plus.n13 plus.n12 161.3
R22 plus.n15 plus.n14 161.3
R23 plus.n17 plus.n0 161.3
R24 plus.n20 plus.n19 161.3
R25 plus.n28 plus.n27 161.3
R26 plus.n30 plus.n29 161.3
R27 plus.n32 plus.n23 161.3
R28 plus.n34 plus.n33 161.3
R29 plus.n36 plus.n35 161.3
R30 plus.n38 plus.n21 161.3
R31 plus.n41 plus.n40 161.3
R32 plus.n12 plus.n11 73.0308
R33 plus.n33 plus.n32 73.0308
R34 plus.n10 plus.n9 67.1884
R35 plus.n15 plus.n1 67.1884
R36 plus.n36 plus.n22 67.1884
R37 plus.n31 plus.n30 67.1884
R38 plus.n6 plus.n3 55.5035
R39 plus.n17 plus.n16 55.5035
R40 plus.n38 plus.n37 55.5035
R41 plus.n27 plus.n24 55.5035
R42 plus.n5 plus.n4 43.8187
R43 plus.n19 plus.n18 43.8187
R44 plus.n40 plus.n39 43.8187
R45 plus.n26 plus.n25 43.8187
R46 plus.n6 plus.n5 29.2126
R47 plus.n18 plus.n17 29.2126
R48 plus.n39 plus.n38 29.2126
R49 plus.n27 plus.n26 29.2126
R50 plus plus.n41 27.3627
R51 plus.n9 plus.n3 17.5278
R52 plus.n16 plus.n15 17.5278
R53 plus.n37 plus.n36 17.5278
R54 plus.n30 plus.n24 17.5278
R55 plus plus.n20 9.83762
R56 plus.n11 plus.n10 5.84292
R57 plus.n12 plus.n1 5.84292
R58 plus.n33 plus.n22 5.84292
R59 plus.n32 plus.n31 5.84292
R60 plus.n8 plus.n7 0.189894
R61 plus.n8 plus.n2 0.189894
R62 plus.n13 plus.n2 0.189894
R63 plus.n14 plus.n13 0.189894
R64 plus.n14 plus.n0 0.189894
R65 plus.n20 plus.n0 0.189894
R66 plus.n41 plus.n21 0.189894
R67 plus.n35 plus.n21 0.189894
R68 plus.n35 plus.n34 0.189894
R69 plus.n34 plus.n23 0.189894
R70 plus.n29 plus.n23 0.189894
R71 plus.n29 plus.n28 0.189894
R72 source.n274 source.n248 289.615
R73 source.n236 source.n210 289.615
R74 source.n204 source.n178 289.615
R75 source.n166 source.n140 289.615
R76 source.n26 source.n0 289.615
R77 source.n64 source.n38 289.615
R78 source.n96 source.n70 289.615
R79 source.n134 source.n108 289.615
R80 source.n259 source.n258 185
R81 source.n256 source.n255 185
R82 source.n265 source.n264 185
R83 source.n267 source.n266 185
R84 source.n252 source.n251 185
R85 source.n273 source.n272 185
R86 source.n275 source.n274 185
R87 source.n221 source.n220 185
R88 source.n218 source.n217 185
R89 source.n227 source.n226 185
R90 source.n229 source.n228 185
R91 source.n214 source.n213 185
R92 source.n235 source.n234 185
R93 source.n237 source.n236 185
R94 source.n189 source.n188 185
R95 source.n186 source.n185 185
R96 source.n195 source.n194 185
R97 source.n197 source.n196 185
R98 source.n182 source.n181 185
R99 source.n203 source.n202 185
R100 source.n205 source.n204 185
R101 source.n151 source.n150 185
R102 source.n148 source.n147 185
R103 source.n157 source.n156 185
R104 source.n159 source.n158 185
R105 source.n144 source.n143 185
R106 source.n165 source.n164 185
R107 source.n167 source.n166 185
R108 source.n27 source.n26 185
R109 source.n25 source.n24 185
R110 source.n4 source.n3 185
R111 source.n19 source.n18 185
R112 source.n17 source.n16 185
R113 source.n8 source.n7 185
R114 source.n11 source.n10 185
R115 source.n65 source.n64 185
R116 source.n63 source.n62 185
R117 source.n42 source.n41 185
R118 source.n57 source.n56 185
R119 source.n55 source.n54 185
R120 source.n46 source.n45 185
R121 source.n49 source.n48 185
R122 source.n97 source.n96 185
R123 source.n95 source.n94 185
R124 source.n74 source.n73 185
R125 source.n89 source.n88 185
R126 source.n87 source.n86 185
R127 source.n78 source.n77 185
R128 source.n81 source.n80 185
R129 source.n135 source.n134 185
R130 source.n133 source.n132 185
R131 source.n112 source.n111 185
R132 source.n127 source.n126 185
R133 source.n125 source.n124 185
R134 source.n116 source.n115 185
R135 source.n119 source.n118 185
R136 source.t6 source.n257 147.661
R137 source.t12 source.n219 147.661
R138 source.t18 source.n187 147.661
R139 source.t23 source.n149 147.661
R140 source.t26 source.n9 147.661
R141 source.t25 source.n47 147.661
R142 source.t15 source.n79 147.661
R143 source.t3 source.n117 147.661
R144 source.n258 source.n255 104.615
R145 source.n265 source.n255 104.615
R146 source.n266 source.n265 104.615
R147 source.n266 source.n251 104.615
R148 source.n273 source.n251 104.615
R149 source.n274 source.n273 104.615
R150 source.n220 source.n217 104.615
R151 source.n227 source.n217 104.615
R152 source.n228 source.n227 104.615
R153 source.n228 source.n213 104.615
R154 source.n235 source.n213 104.615
R155 source.n236 source.n235 104.615
R156 source.n188 source.n185 104.615
R157 source.n195 source.n185 104.615
R158 source.n196 source.n195 104.615
R159 source.n196 source.n181 104.615
R160 source.n203 source.n181 104.615
R161 source.n204 source.n203 104.615
R162 source.n150 source.n147 104.615
R163 source.n157 source.n147 104.615
R164 source.n158 source.n157 104.615
R165 source.n158 source.n143 104.615
R166 source.n165 source.n143 104.615
R167 source.n166 source.n165 104.615
R168 source.n26 source.n25 104.615
R169 source.n25 source.n3 104.615
R170 source.n18 source.n3 104.615
R171 source.n18 source.n17 104.615
R172 source.n17 source.n7 104.615
R173 source.n10 source.n7 104.615
R174 source.n64 source.n63 104.615
R175 source.n63 source.n41 104.615
R176 source.n56 source.n41 104.615
R177 source.n56 source.n55 104.615
R178 source.n55 source.n45 104.615
R179 source.n48 source.n45 104.615
R180 source.n96 source.n95 104.615
R181 source.n95 source.n73 104.615
R182 source.n88 source.n73 104.615
R183 source.n88 source.n87 104.615
R184 source.n87 source.n77 104.615
R185 source.n80 source.n77 104.615
R186 source.n134 source.n133 104.615
R187 source.n133 source.n111 104.615
R188 source.n126 source.n111 104.615
R189 source.n126 source.n125 104.615
R190 source.n125 source.n115 104.615
R191 source.n118 source.n115 104.615
R192 source.n258 source.t6 52.3082
R193 source.n220 source.t12 52.3082
R194 source.n188 source.t18 52.3082
R195 source.n150 source.t23 52.3082
R196 source.n10 source.t26 52.3082
R197 source.n48 source.t25 52.3082
R198 source.n80 source.t15 52.3082
R199 source.n118 source.t3 52.3082
R200 source.n33 source.n32 50.512
R201 source.n35 source.n34 50.512
R202 source.n37 source.n36 50.512
R203 source.n103 source.n102 50.512
R204 source.n105 source.n104 50.512
R205 source.n107 source.n106 50.512
R206 source.n247 source.n246 50.5119
R207 source.n245 source.n244 50.5119
R208 source.n243 source.n242 50.5119
R209 source.n177 source.n176 50.5119
R210 source.n175 source.n174 50.5119
R211 source.n173 source.n172 50.5119
R212 source.n279 source.n278 32.1853
R213 source.n241 source.n240 32.1853
R214 source.n209 source.n208 32.1853
R215 source.n171 source.n170 32.1853
R216 source.n31 source.n30 32.1853
R217 source.n69 source.n68 32.1853
R218 source.n101 source.n100 32.1853
R219 source.n139 source.n138 32.1853
R220 source.n171 source.n139 17.2423
R221 source.n259 source.n257 15.6674
R222 source.n221 source.n219 15.6674
R223 source.n189 source.n187 15.6674
R224 source.n151 source.n149 15.6674
R225 source.n11 source.n9 15.6674
R226 source.n49 source.n47 15.6674
R227 source.n81 source.n79 15.6674
R228 source.n119 source.n117 15.6674
R229 source.n260 source.n256 12.8005
R230 source.n222 source.n218 12.8005
R231 source.n190 source.n186 12.8005
R232 source.n152 source.n148 12.8005
R233 source.n12 source.n8 12.8005
R234 source.n50 source.n46 12.8005
R235 source.n82 source.n78 12.8005
R236 source.n120 source.n116 12.8005
R237 source.n264 source.n263 12.0247
R238 source.n226 source.n225 12.0247
R239 source.n194 source.n193 12.0247
R240 source.n156 source.n155 12.0247
R241 source.n16 source.n15 12.0247
R242 source.n54 source.n53 12.0247
R243 source.n86 source.n85 12.0247
R244 source.n124 source.n123 12.0247
R245 source.n280 source.n31 11.7293
R246 source.n267 source.n254 11.249
R247 source.n229 source.n216 11.249
R248 source.n197 source.n184 11.249
R249 source.n159 source.n146 11.249
R250 source.n19 source.n6 11.249
R251 source.n57 source.n44 11.249
R252 source.n89 source.n76 11.249
R253 source.n127 source.n114 11.249
R254 source.n268 source.n252 10.4732
R255 source.n230 source.n214 10.4732
R256 source.n198 source.n182 10.4732
R257 source.n160 source.n144 10.4732
R258 source.n20 source.n4 10.4732
R259 source.n58 source.n42 10.4732
R260 source.n90 source.n74 10.4732
R261 source.n128 source.n112 10.4732
R262 source.n272 source.n271 9.69747
R263 source.n234 source.n233 9.69747
R264 source.n202 source.n201 9.69747
R265 source.n164 source.n163 9.69747
R266 source.n24 source.n23 9.69747
R267 source.n62 source.n61 9.69747
R268 source.n94 source.n93 9.69747
R269 source.n132 source.n131 9.69747
R270 source.n278 source.n277 9.45567
R271 source.n240 source.n239 9.45567
R272 source.n208 source.n207 9.45567
R273 source.n170 source.n169 9.45567
R274 source.n30 source.n29 9.45567
R275 source.n68 source.n67 9.45567
R276 source.n100 source.n99 9.45567
R277 source.n138 source.n137 9.45567
R278 source.n277 source.n276 9.3005
R279 source.n250 source.n249 9.3005
R280 source.n271 source.n270 9.3005
R281 source.n269 source.n268 9.3005
R282 source.n254 source.n253 9.3005
R283 source.n263 source.n262 9.3005
R284 source.n261 source.n260 9.3005
R285 source.n239 source.n238 9.3005
R286 source.n212 source.n211 9.3005
R287 source.n233 source.n232 9.3005
R288 source.n231 source.n230 9.3005
R289 source.n216 source.n215 9.3005
R290 source.n225 source.n224 9.3005
R291 source.n223 source.n222 9.3005
R292 source.n207 source.n206 9.3005
R293 source.n180 source.n179 9.3005
R294 source.n201 source.n200 9.3005
R295 source.n199 source.n198 9.3005
R296 source.n184 source.n183 9.3005
R297 source.n193 source.n192 9.3005
R298 source.n191 source.n190 9.3005
R299 source.n169 source.n168 9.3005
R300 source.n142 source.n141 9.3005
R301 source.n163 source.n162 9.3005
R302 source.n161 source.n160 9.3005
R303 source.n146 source.n145 9.3005
R304 source.n155 source.n154 9.3005
R305 source.n153 source.n152 9.3005
R306 source.n29 source.n28 9.3005
R307 source.n2 source.n1 9.3005
R308 source.n23 source.n22 9.3005
R309 source.n21 source.n20 9.3005
R310 source.n6 source.n5 9.3005
R311 source.n15 source.n14 9.3005
R312 source.n13 source.n12 9.3005
R313 source.n67 source.n66 9.3005
R314 source.n40 source.n39 9.3005
R315 source.n61 source.n60 9.3005
R316 source.n59 source.n58 9.3005
R317 source.n44 source.n43 9.3005
R318 source.n53 source.n52 9.3005
R319 source.n51 source.n50 9.3005
R320 source.n99 source.n98 9.3005
R321 source.n72 source.n71 9.3005
R322 source.n93 source.n92 9.3005
R323 source.n91 source.n90 9.3005
R324 source.n76 source.n75 9.3005
R325 source.n85 source.n84 9.3005
R326 source.n83 source.n82 9.3005
R327 source.n137 source.n136 9.3005
R328 source.n110 source.n109 9.3005
R329 source.n131 source.n130 9.3005
R330 source.n129 source.n128 9.3005
R331 source.n114 source.n113 9.3005
R332 source.n123 source.n122 9.3005
R333 source.n121 source.n120 9.3005
R334 source.n275 source.n250 8.92171
R335 source.n237 source.n212 8.92171
R336 source.n205 source.n180 8.92171
R337 source.n167 source.n142 8.92171
R338 source.n27 source.n2 8.92171
R339 source.n65 source.n40 8.92171
R340 source.n97 source.n72 8.92171
R341 source.n135 source.n110 8.92171
R342 source.n276 source.n248 8.14595
R343 source.n238 source.n210 8.14595
R344 source.n206 source.n178 8.14595
R345 source.n168 source.n140 8.14595
R346 source.n28 source.n0 8.14595
R347 source.n66 source.n38 8.14595
R348 source.n98 source.n70 8.14595
R349 source.n136 source.n108 8.14595
R350 source.n278 source.n248 5.81868
R351 source.n240 source.n210 5.81868
R352 source.n208 source.n178 5.81868
R353 source.n170 source.n140 5.81868
R354 source.n30 source.n0 5.81868
R355 source.n68 source.n38 5.81868
R356 source.n100 source.n70 5.81868
R357 source.n138 source.n108 5.81868
R358 source.n280 source.n279 5.51343
R359 source.n276 source.n275 5.04292
R360 source.n238 source.n237 5.04292
R361 source.n206 source.n205 5.04292
R362 source.n168 source.n167 5.04292
R363 source.n28 source.n27 5.04292
R364 source.n66 source.n65 5.04292
R365 source.n98 source.n97 5.04292
R366 source.n136 source.n135 5.04292
R367 source.n261 source.n257 4.38594
R368 source.n223 source.n219 4.38594
R369 source.n191 source.n187 4.38594
R370 source.n153 source.n149 4.38594
R371 source.n13 source.n9 4.38594
R372 source.n51 source.n47 4.38594
R373 source.n83 source.n79 4.38594
R374 source.n121 source.n117 4.38594
R375 source.n272 source.n250 4.26717
R376 source.n234 source.n212 4.26717
R377 source.n202 source.n180 4.26717
R378 source.n164 source.n142 4.26717
R379 source.n24 source.n2 4.26717
R380 source.n62 source.n40 4.26717
R381 source.n94 source.n72 4.26717
R382 source.n132 source.n110 4.26717
R383 source.n271 source.n252 3.49141
R384 source.n233 source.n214 3.49141
R385 source.n201 source.n182 3.49141
R386 source.n163 source.n144 3.49141
R387 source.n23 source.n4 3.49141
R388 source.n61 source.n42 3.49141
R389 source.n93 source.n74 3.49141
R390 source.n131 source.n112 3.49141
R391 source.n246 source.t13 3.3005
R392 source.n246 source.t11 3.3005
R393 source.n244 source.t1 3.3005
R394 source.n244 source.t10 3.3005
R395 source.n242 source.t5 3.3005
R396 source.n242 source.t0 3.3005
R397 source.n176 source.t22 3.3005
R398 source.n176 source.t29 3.3005
R399 source.n174 source.t19 3.3005
R400 source.n174 source.t17 3.3005
R401 source.n172 source.t24 3.3005
R402 source.n172 source.t28 3.3005
R403 source.n32 source.t30 3.3005
R404 source.n32 source.t21 3.3005
R405 source.n34 source.t16 3.3005
R406 source.n34 source.t27 3.3005
R407 source.n36 source.t31 3.3005
R408 source.n36 source.t20 3.3005
R409 source.n102 source.t4 3.3005
R410 source.n102 source.t2 3.3005
R411 source.n104 source.t14 3.3005
R412 source.n104 source.t8 3.3005
R413 source.n106 source.t7 3.3005
R414 source.n106 source.t9 3.3005
R415 source.n268 source.n267 2.71565
R416 source.n230 source.n229 2.71565
R417 source.n198 source.n197 2.71565
R418 source.n160 source.n159 2.71565
R419 source.n20 source.n19 2.71565
R420 source.n58 source.n57 2.71565
R421 source.n90 source.n89 2.71565
R422 source.n128 source.n127 2.71565
R423 source.n264 source.n254 1.93989
R424 source.n226 source.n216 1.93989
R425 source.n194 source.n184 1.93989
R426 source.n156 source.n146 1.93989
R427 source.n16 source.n6 1.93989
R428 source.n54 source.n44 1.93989
R429 source.n86 source.n76 1.93989
R430 source.n124 source.n114 1.93989
R431 source.n263 source.n256 1.16414
R432 source.n225 source.n218 1.16414
R433 source.n193 source.n186 1.16414
R434 source.n155 source.n148 1.16414
R435 source.n15 source.n8 1.16414
R436 source.n53 source.n46 1.16414
R437 source.n85 source.n78 1.16414
R438 source.n123 source.n116 1.16414
R439 source.n139 source.n107 0.5005
R440 source.n107 source.n105 0.5005
R441 source.n105 source.n103 0.5005
R442 source.n103 source.n101 0.5005
R443 source.n69 source.n37 0.5005
R444 source.n37 source.n35 0.5005
R445 source.n35 source.n33 0.5005
R446 source.n33 source.n31 0.5005
R447 source.n173 source.n171 0.5005
R448 source.n175 source.n173 0.5005
R449 source.n177 source.n175 0.5005
R450 source.n209 source.n177 0.5005
R451 source.n243 source.n241 0.5005
R452 source.n245 source.n243 0.5005
R453 source.n247 source.n245 0.5005
R454 source.n279 source.n247 0.5005
R455 source.n101 source.n69 0.470328
R456 source.n241 source.n209 0.470328
R457 source.n260 source.n259 0.388379
R458 source.n222 source.n221 0.388379
R459 source.n190 source.n189 0.388379
R460 source.n152 source.n151 0.388379
R461 source.n12 source.n11 0.388379
R462 source.n50 source.n49 0.388379
R463 source.n82 source.n81 0.388379
R464 source.n120 source.n119 0.388379
R465 source source.n280 0.188
R466 source.n262 source.n261 0.155672
R467 source.n262 source.n253 0.155672
R468 source.n269 source.n253 0.155672
R469 source.n270 source.n269 0.155672
R470 source.n270 source.n249 0.155672
R471 source.n277 source.n249 0.155672
R472 source.n224 source.n223 0.155672
R473 source.n224 source.n215 0.155672
R474 source.n231 source.n215 0.155672
R475 source.n232 source.n231 0.155672
R476 source.n232 source.n211 0.155672
R477 source.n239 source.n211 0.155672
R478 source.n192 source.n191 0.155672
R479 source.n192 source.n183 0.155672
R480 source.n199 source.n183 0.155672
R481 source.n200 source.n199 0.155672
R482 source.n200 source.n179 0.155672
R483 source.n207 source.n179 0.155672
R484 source.n154 source.n153 0.155672
R485 source.n154 source.n145 0.155672
R486 source.n161 source.n145 0.155672
R487 source.n162 source.n161 0.155672
R488 source.n162 source.n141 0.155672
R489 source.n169 source.n141 0.155672
R490 source.n29 source.n1 0.155672
R491 source.n22 source.n1 0.155672
R492 source.n22 source.n21 0.155672
R493 source.n21 source.n5 0.155672
R494 source.n14 source.n5 0.155672
R495 source.n14 source.n13 0.155672
R496 source.n67 source.n39 0.155672
R497 source.n60 source.n39 0.155672
R498 source.n60 source.n59 0.155672
R499 source.n59 source.n43 0.155672
R500 source.n52 source.n43 0.155672
R501 source.n52 source.n51 0.155672
R502 source.n99 source.n71 0.155672
R503 source.n92 source.n71 0.155672
R504 source.n92 source.n91 0.155672
R505 source.n91 source.n75 0.155672
R506 source.n84 source.n75 0.155672
R507 source.n84 source.n83 0.155672
R508 source.n137 source.n109 0.155672
R509 source.n130 source.n109 0.155672
R510 source.n130 source.n129 0.155672
R511 source.n129 source.n113 0.155672
R512 source.n122 source.n113 0.155672
R513 source.n122 source.n121 0.155672
R514 drain_left.n9 drain_left.n7 67.6908
R515 drain_left.n5 drain_left.n3 67.6907
R516 drain_left.n2 drain_left.n0 67.6907
R517 drain_left.n11 drain_left.n10 67.1908
R518 drain_left.n9 drain_left.n8 67.1908
R519 drain_left.n13 drain_left.n12 67.1907
R520 drain_left.n5 drain_left.n4 67.1907
R521 drain_left.n2 drain_left.n1 67.1907
R522 drain_left drain_left.n6 26.0716
R523 drain_left drain_left.n13 6.15322
R524 drain_left.n3 drain_left.t9 3.3005
R525 drain_left.n3 drain_left.t4 3.3005
R526 drain_left.n4 drain_left.t3 3.3005
R527 drain_left.n4 drain_left.t13 3.3005
R528 drain_left.n1 drain_left.t8 3.3005
R529 drain_left.n1 drain_left.t2 3.3005
R530 drain_left.n0 drain_left.t0 3.3005
R531 drain_left.n0 drain_left.t10 3.3005
R532 drain_left.n12 drain_left.t7 3.3005
R533 drain_left.n12 drain_left.t12 3.3005
R534 drain_left.n10 drain_left.t6 3.3005
R535 drain_left.n10 drain_left.t1 3.3005
R536 drain_left.n8 drain_left.t5 3.3005
R537 drain_left.n8 drain_left.t15 3.3005
R538 drain_left.n7 drain_left.t11 3.3005
R539 drain_left.n7 drain_left.t14 3.3005
R540 drain_left.n11 drain_left.n9 0.5005
R541 drain_left.n13 drain_left.n11 0.5005
R542 drain_left.n6 drain_left.n5 0.195154
R543 drain_left.n6 drain_left.n2 0.195154
R544 minus.n19 minus.t3 744.617
R545 minus.n4 minus.t11 744.617
R546 minus.n40 minus.t4 744.617
R547 minus.n25 minus.t10 744.617
R548 minus.n18 minus.t14 703.721
R549 minus.n16 minus.t5 703.721
R550 minus.n1 minus.t13 703.721
R551 minus.n10 minus.t0 703.721
R552 minus.n3 minus.t9 703.721
R553 minus.n5 minus.t1 703.721
R554 minus.n39 minus.t6 703.721
R555 minus.n37 minus.t8 703.721
R556 minus.n22 minus.t15 703.721
R557 minus.n31 minus.t2 703.721
R558 minus.n24 minus.t7 703.721
R559 minus.n26 minus.t12 703.721
R560 minus.n7 minus.n4 161.489
R561 minus.n28 minus.n25 161.489
R562 minus.n20 minus.n19 161.3
R563 minus.n17 minus.n0 161.3
R564 minus.n15 minus.n14 161.3
R565 minus.n13 minus.n12 161.3
R566 minus.n11 minus.n2 161.3
R567 minus.n9 minus.n8 161.3
R568 minus.n7 minus.n6 161.3
R569 minus.n41 minus.n40 161.3
R570 minus.n38 minus.n21 161.3
R571 minus.n36 minus.n35 161.3
R572 minus.n34 minus.n33 161.3
R573 minus.n32 minus.n23 161.3
R574 minus.n30 minus.n29 161.3
R575 minus.n28 minus.n27 161.3
R576 minus.n12 minus.n11 73.0308
R577 minus.n33 minus.n32 73.0308
R578 minus.n15 minus.n1 67.1884
R579 minus.n10 minus.n9 67.1884
R580 minus.n31 minus.n30 67.1884
R581 minus.n36 minus.n22 67.1884
R582 minus.n17 minus.n16 55.5035
R583 minus.n6 minus.n3 55.5035
R584 minus.n27 minus.n24 55.5035
R585 minus.n38 minus.n37 55.5035
R586 minus.n19 minus.n18 43.8187
R587 minus.n5 minus.n4 43.8187
R588 minus.n26 minus.n25 43.8187
R589 minus.n40 minus.n39 43.8187
R590 minus.n42 minus.n20 31.2088
R591 minus.n18 minus.n17 29.2126
R592 minus.n6 minus.n5 29.2126
R593 minus.n27 minus.n26 29.2126
R594 minus.n39 minus.n38 29.2126
R595 minus.n16 minus.n15 17.5278
R596 minus.n9 minus.n3 17.5278
R597 minus.n30 minus.n24 17.5278
R598 minus.n37 minus.n36 17.5278
R599 minus.n42 minus.n41 6.46641
R600 minus.n12 minus.n1 5.84292
R601 minus.n11 minus.n10 5.84292
R602 minus.n32 minus.n31 5.84292
R603 minus.n33 minus.n22 5.84292
R604 minus.n20 minus.n0 0.189894
R605 minus.n14 minus.n0 0.189894
R606 minus.n14 minus.n13 0.189894
R607 minus.n13 minus.n2 0.189894
R608 minus.n8 minus.n2 0.189894
R609 minus.n8 minus.n7 0.189894
R610 minus.n29 minus.n28 0.189894
R611 minus.n29 minus.n23 0.189894
R612 minus.n34 minus.n23 0.189894
R613 minus.n35 minus.n34 0.189894
R614 minus.n35 minus.n21 0.189894
R615 minus.n41 minus.n21 0.189894
R616 minus minus.n42 0.188
R617 drain_right.n9 drain_right.n7 67.6907
R618 drain_right.n5 drain_right.n3 67.6907
R619 drain_right.n2 drain_right.n0 67.6907
R620 drain_right.n9 drain_right.n8 67.1908
R621 drain_right.n11 drain_right.n10 67.1908
R622 drain_right.n13 drain_right.n12 67.1908
R623 drain_right.n5 drain_right.n4 67.1907
R624 drain_right.n2 drain_right.n1 67.1907
R625 drain_right drain_right.n6 25.5184
R626 drain_right drain_right.n13 6.15322
R627 drain_right.n3 drain_right.t9 3.3005
R628 drain_right.n3 drain_right.t11 3.3005
R629 drain_right.n4 drain_right.t0 3.3005
R630 drain_right.n4 drain_right.t7 3.3005
R631 drain_right.n1 drain_right.t8 3.3005
R632 drain_right.n1 drain_right.t13 3.3005
R633 drain_right.n0 drain_right.t5 3.3005
R634 drain_right.n0 drain_right.t3 3.3005
R635 drain_right.n7 drain_right.t14 3.3005
R636 drain_right.n7 drain_right.t4 3.3005
R637 drain_right.n8 drain_right.t15 3.3005
R638 drain_right.n8 drain_right.t6 3.3005
R639 drain_right.n10 drain_right.t10 3.3005
R640 drain_right.n10 drain_right.t2 3.3005
R641 drain_right.n12 drain_right.t12 3.3005
R642 drain_right.n12 drain_right.t1 3.3005
R643 drain_right.n13 drain_right.n11 0.5005
R644 drain_right.n11 drain_right.n9 0.5005
R645 drain_right.n6 drain_right.n5 0.195154
R646 drain_right.n6 drain_right.n2 0.195154
C0 minus source 2.79229f
C1 plus source 2.80631f
C2 plus minus 4.23906f
C3 drain_right drain_left 0.897273f
C4 drain_left source 18.0015f
C5 drain_left minus 0.171252f
C6 plus drain_left 3.01638f
C7 drain_right source 18.0015f
C8 drain_right minus 2.84604f
C9 plus drain_right 0.324551f
C10 drain_right a_n1760_n2088# 5.22538f
C11 drain_left a_n1760_n2088# 5.50874f
C12 source a_n1760_n2088# 5.297333f
C13 minus a_n1760_n2088# 6.37946f
C14 plus a_n1760_n2088# 7.97981f
C15 drain_right.t5 a_n1760_n2088# 0.165914f
C16 drain_right.t3 a_n1760_n2088# 0.165914f
C17 drain_right.n0 a_n1760_n2088# 1.38676f
C18 drain_right.t8 a_n1760_n2088# 0.165914f
C19 drain_right.t13 a_n1760_n2088# 0.165914f
C20 drain_right.n1 a_n1760_n2088# 1.38372f
C21 drain_right.n2 a_n1760_n2088# 0.774335f
C22 drain_right.t9 a_n1760_n2088# 0.165914f
C23 drain_right.t11 a_n1760_n2088# 0.165914f
C24 drain_right.n3 a_n1760_n2088# 1.38676f
C25 drain_right.t0 a_n1760_n2088# 0.165914f
C26 drain_right.t7 a_n1760_n2088# 0.165914f
C27 drain_right.n4 a_n1760_n2088# 1.38372f
C28 drain_right.n5 a_n1760_n2088# 0.774335f
C29 drain_right.n6 a_n1760_n2088# 1.15129f
C30 drain_right.t14 a_n1760_n2088# 0.165914f
C31 drain_right.t4 a_n1760_n2088# 0.165914f
C32 drain_right.n7 a_n1760_n2088# 1.38676f
C33 drain_right.t15 a_n1760_n2088# 0.165914f
C34 drain_right.t6 a_n1760_n2088# 0.165914f
C35 drain_right.n8 a_n1760_n2088# 1.38373f
C36 drain_right.n9 a_n1760_n2088# 0.80459f
C37 drain_right.t10 a_n1760_n2088# 0.165914f
C38 drain_right.t2 a_n1760_n2088# 0.165914f
C39 drain_right.n10 a_n1760_n2088# 1.38373f
C40 drain_right.n11 a_n1760_n2088# 0.396762f
C41 drain_right.t12 a_n1760_n2088# 0.165914f
C42 drain_right.t1 a_n1760_n2088# 0.165914f
C43 drain_right.n12 a_n1760_n2088# 1.38373f
C44 drain_right.n13 a_n1760_n2088# 0.685603f
C45 minus.n0 a_n1760_n2088# 0.051532f
C46 minus.t3 a_n1760_n2088# 0.225987f
C47 minus.t14 a_n1760_n2088# 0.220237f
C48 minus.t5 a_n1760_n2088# 0.220237f
C49 minus.t13 a_n1760_n2088# 0.220237f
C50 minus.n1 a_n1760_n2088# 0.10374f
C51 minus.n2 a_n1760_n2088# 0.051532f
C52 minus.t0 a_n1760_n2088# 0.220237f
C53 minus.t9 a_n1760_n2088# 0.220237f
C54 minus.n3 a_n1760_n2088# 0.10374f
C55 minus.t11 a_n1760_n2088# 0.225987f
C56 minus.n4 a_n1760_n2088# 0.118652f
C57 minus.t1 a_n1760_n2088# 0.220237f
C58 minus.n5 a_n1760_n2088# 0.10374f
C59 minus.n6 a_n1760_n2088# 0.019637f
C60 minus.n7 a_n1760_n2088# 0.112842f
C61 minus.n8 a_n1760_n2088# 0.051532f
C62 minus.n9 a_n1760_n2088# 0.019637f
C63 minus.n10 a_n1760_n2088# 0.10374f
C64 minus.n11 a_n1760_n2088# 0.018366f
C65 minus.n12 a_n1760_n2088# 0.018366f
C66 minus.n13 a_n1760_n2088# 0.051532f
C67 minus.n14 a_n1760_n2088# 0.051532f
C68 minus.n15 a_n1760_n2088# 0.019637f
C69 minus.n16 a_n1760_n2088# 0.10374f
C70 minus.n17 a_n1760_n2088# 0.019637f
C71 minus.n18 a_n1760_n2088# 0.10374f
C72 minus.n19 a_n1760_n2088# 0.11858f
C73 minus.n20 a_n1760_n2088# 1.43162f
C74 minus.n21 a_n1760_n2088# 0.051532f
C75 minus.t6 a_n1760_n2088# 0.220237f
C76 minus.t8 a_n1760_n2088# 0.220237f
C77 minus.t15 a_n1760_n2088# 0.220237f
C78 minus.n22 a_n1760_n2088# 0.10374f
C79 minus.n23 a_n1760_n2088# 0.051532f
C80 minus.t2 a_n1760_n2088# 0.220237f
C81 minus.t7 a_n1760_n2088# 0.220237f
C82 minus.n24 a_n1760_n2088# 0.10374f
C83 minus.t10 a_n1760_n2088# 0.225987f
C84 minus.n25 a_n1760_n2088# 0.118652f
C85 minus.t12 a_n1760_n2088# 0.220237f
C86 minus.n26 a_n1760_n2088# 0.10374f
C87 minus.n27 a_n1760_n2088# 0.019637f
C88 minus.n28 a_n1760_n2088# 0.112842f
C89 minus.n29 a_n1760_n2088# 0.051532f
C90 minus.n30 a_n1760_n2088# 0.019637f
C91 minus.n31 a_n1760_n2088# 0.10374f
C92 minus.n32 a_n1760_n2088# 0.018366f
C93 minus.n33 a_n1760_n2088# 0.018366f
C94 minus.n34 a_n1760_n2088# 0.051532f
C95 minus.n35 a_n1760_n2088# 0.051532f
C96 minus.n36 a_n1760_n2088# 0.019637f
C97 minus.n37 a_n1760_n2088# 0.10374f
C98 minus.n38 a_n1760_n2088# 0.019637f
C99 minus.n39 a_n1760_n2088# 0.10374f
C100 minus.t4 a_n1760_n2088# 0.225987f
C101 minus.n40 a_n1760_n2088# 0.11858f
C102 minus.n41 a_n1760_n2088# 0.33282f
C103 minus.n42 a_n1760_n2088# 1.76403f
C104 drain_left.t0 a_n1760_n2088# 0.166414f
C105 drain_left.t10 a_n1760_n2088# 0.166414f
C106 drain_left.n0 a_n1760_n2088# 1.39094f
C107 drain_left.t8 a_n1760_n2088# 0.166414f
C108 drain_left.t2 a_n1760_n2088# 0.166414f
C109 drain_left.n1 a_n1760_n2088# 1.3879f
C110 drain_left.n2 a_n1760_n2088# 0.776669f
C111 drain_left.t9 a_n1760_n2088# 0.166414f
C112 drain_left.t4 a_n1760_n2088# 0.166414f
C113 drain_left.n3 a_n1760_n2088# 1.39094f
C114 drain_left.t3 a_n1760_n2088# 0.166414f
C115 drain_left.t13 a_n1760_n2088# 0.166414f
C116 drain_left.n4 a_n1760_n2088# 1.3879f
C117 drain_left.n5 a_n1760_n2088# 0.776669f
C118 drain_left.n6 a_n1760_n2088# 1.2261f
C119 drain_left.t11 a_n1760_n2088# 0.166414f
C120 drain_left.t14 a_n1760_n2088# 0.166414f
C121 drain_left.n7 a_n1760_n2088# 1.39095f
C122 drain_left.t5 a_n1760_n2088# 0.166414f
C123 drain_left.t15 a_n1760_n2088# 0.166414f
C124 drain_left.n8 a_n1760_n2088# 1.3879f
C125 drain_left.n9 a_n1760_n2088# 0.807008f
C126 drain_left.t6 a_n1760_n2088# 0.166414f
C127 drain_left.t1 a_n1760_n2088# 0.166414f
C128 drain_left.n10 a_n1760_n2088# 1.3879f
C129 drain_left.n11 a_n1760_n2088# 0.397958f
C130 drain_left.t7 a_n1760_n2088# 0.166414f
C131 drain_left.t12 a_n1760_n2088# 0.166414f
C132 drain_left.n12 a_n1760_n2088# 1.3879f
C133 drain_left.n13 a_n1760_n2088# 0.687677f
C134 source.n0 a_n1760_n2088# 0.043614f
C135 source.n1 a_n1760_n2088# 0.031029f
C136 source.n2 a_n1760_n2088# 0.016674f
C137 source.n3 a_n1760_n2088# 0.039411f
C138 source.n4 a_n1760_n2088# 0.017655f
C139 source.n5 a_n1760_n2088# 0.031029f
C140 source.n6 a_n1760_n2088# 0.016674f
C141 source.n7 a_n1760_n2088# 0.039411f
C142 source.n8 a_n1760_n2088# 0.017655f
C143 source.n9 a_n1760_n2088# 0.132784f
C144 source.t26 a_n1760_n2088# 0.064235f
C145 source.n10 a_n1760_n2088# 0.029558f
C146 source.n11 a_n1760_n2088# 0.02328f
C147 source.n12 a_n1760_n2088# 0.016674f
C148 source.n13 a_n1760_n2088# 0.738314f
C149 source.n14 a_n1760_n2088# 0.031029f
C150 source.n15 a_n1760_n2088# 0.016674f
C151 source.n16 a_n1760_n2088# 0.017655f
C152 source.n17 a_n1760_n2088# 0.039411f
C153 source.n18 a_n1760_n2088# 0.039411f
C154 source.n19 a_n1760_n2088# 0.017655f
C155 source.n20 a_n1760_n2088# 0.016674f
C156 source.n21 a_n1760_n2088# 0.031029f
C157 source.n22 a_n1760_n2088# 0.031029f
C158 source.n23 a_n1760_n2088# 0.016674f
C159 source.n24 a_n1760_n2088# 0.017655f
C160 source.n25 a_n1760_n2088# 0.039411f
C161 source.n26 a_n1760_n2088# 0.085318f
C162 source.n27 a_n1760_n2088# 0.017655f
C163 source.n28 a_n1760_n2088# 0.016674f
C164 source.n29 a_n1760_n2088# 0.071723f
C165 source.n30 a_n1760_n2088# 0.047739f
C166 source.n31 a_n1760_n2088# 0.744203f
C167 source.t30 a_n1760_n2088# 0.147122f
C168 source.t21 a_n1760_n2088# 0.147122f
C169 source.n32 a_n1760_n2088# 1.1458f
C170 source.n33 a_n1760_n2088# 0.390854f
C171 source.t16 a_n1760_n2088# 0.147122f
C172 source.t27 a_n1760_n2088# 0.147122f
C173 source.n34 a_n1760_n2088# 1.1458f
C174 source.n35 a_n1760_n2088# 0.390854f
C175 source.t31 a_n1760_n2088# 0.147122f
C176 source.t20 a_n1760_n2088# 0.147122f
C177 source.n36 a_n1760_n2088# 1.1458f
C178 source.n37 a_n1760_n2088# 0.390854f
C179 source.n38 a_n1760_n2088# 0.043614f
C180 source.n39 a_n1760_n2088# 0.031029f
C181 source.n40 a_n1760_n2088# 0.016674f
C182 source.n41 a_n1760_n2088# 0.039411f
C183 source.n42 a_n1760_n2088# 0.017655f
C184 source.n43 a_n1760_n2088# 0.031029f
C185 source.n44 a_n1760_n2088# 0.016674f
C186 source.n45 a_n1760_n2088# 0.039411f
C187 source.n46 a_n1760_n2088# 0.017655f
C188 source.n47 a_n1760_n2088# 0.132784f
C189 source.t25 a_n1760_n2088# 0.064235f
C190 source.n48 a_n1760_n2088# 0.029558f
C191 source.n49 a_n1760_n2088# 0.02328f
C192 source.n50 a_n1760_n2088# 0.016674f
C193 source.n51 a_n1760_n2088# 0.738314f
C194 source.n52 a_n1760_n2088# 0.031029f
C195 source.n53 a_n1760_n2088# 0.016674f
C196 source.n54 a_n1760_n2088# 0.017655f
C197 source.n55 a_n1760_n2088# 0.039411f
C198 source.n56 a_n1760_n2088# 0.039411f
C199 source.n57 a_n1760_n2088# 0.017655f
C200 source.n58 a_n1760_n2088# 0.016674f
C201 source.n59 a_n1760_n2088# 0.031029f
C202 source.n60 a_n1760_n2088# 0.031029f
C203 source.n61 a_n1760_n2088# 0.016674f
C204 source.n62 a_n1760_n2088# 0.017655f
C205 source.n63 a_n1760_n2088# 0.039411f
C206 source.n64 a_n1760_n2088# 0.085318f
C207 source.n65 a_n1760_n2088# 0.017655f
C208 source.n66 a_n1760_n2088# 0.016674f
C209 source.n67 a_n1760_n2088# 0.071723f
C210 source.n68 a_n1760_n2088# 0.047739f
C211 source.n69 a_n1760_n2088# 0.123468f
C212 source.n70 a_n1760_n2088# 0.043614f
C213 source.n71 a_n1760_n2088# 0.031029f
C214 source.n72 a_n1760_n2088# 0.016674f
C215 source.n73 a_n1760_n2088# 0.039411f
C216 source.n74 a_n1760_n2088# 0.017655f
C217 source.n75 a_n1760_n2088# 0.031029f
C218 source.n76 a_n1760_n2088# 0.016674f
C219 source.n77 a_n1760_n2088# 0.039411f
C220 source.n78 a_n1760_n2088# 0.017655f
C221 source.n79 a_n1760_n2088# 0.132784f
C222 source.t15 a_n1760_n2088# 0.064235f
C223 source.n80 a_n1760_n2088# 0.029558f
C224 source.n81 a_n1760_n2088# 0.02328f
C225 source.n82 a_n1760_n2088# 0.016674f
C226 source.n83 a_n1760_n2088# 0.738314f
C227 source.n84 a_n1760_n2088# 0.031029f
C228 source.n85 a_n1760_n2088# 0.016674f
C229 source.n86 a_n1760_n2088# 0.017655f
C230 source.n87 a_n1760_n2088# 0.039411f
C231 source.n88 a_n1760_n2088# 0.039411f
C232 source.n89 a_n1760_n2088# 0.017655f
C233 source.n90 a_n1760_n2088# 0.016674f
C234 source.n91 a_n1760_n2088# 0.031029f
C235 source.n92 a_n1760_n2088# 0.031029f
C236 source.n93 a_n1760_n2088# 0.016674f
C237 source.n94 a_n1760_n2088# 0.017655f
C238 source.n95 a_n1760_n2088# 0.039411f
C239 source.n96 a_n1760_n2088# 0.085318f
C240 source.n97 a_n1760_n2088# 0.017655f
C241 source.n98 a_n1760_n2088# 0.016674f
C242 source.n99 a_n1760_n2088# 0.071723f
C243 source.n100 a_n1760_n2088# 0.047739f
C244 source.n101 a_n1760_n2088# 0.123468f
C245 source.t4 a_n1760_n2088# 0.147122f
C246 source.t2 a_n1760_n2088# 0.147122f
C247 source.n102 a_n1760_n2088# 1.1458f
C248 source.n103 a_n1760_n2088# 0.390854f
C249 source.t14 a_n1760_n2088# 0.147122f
C250 source.t8 a_n1760_n2088# 0.147122f
C251 source.n104 a_n1760_n2088# 1.1458f
C252 source.n105 a_n1760_n2088# 0.390854f
C253 source.t7 a_n1760_n2088# 0.147122f
C254 source.t9 a_n1760_n2088# 0.147122f
C255 source.n106 a_n1760_n2088# 1.1458f
C256 source.n107 a_n1760_n2088# 0.390854f
C257 source.n108 a_n1760_n2088# 0.043614f
C258 source.n109 a_n1760_n2088# 0.031029f
C259 source.n110 a_n1760_n2088# 0.016674f
C260 source.n111 a_n1760_n2088# 0.039411f
C261 source.n112 a_n1760_n2088# 0.017655f
C262 source.n113 a_n1760_n2088# 0.031029f
C263 source.n114 a_n1760_n2088# 0.016674f
C264 source.n115 a_n1760_n2088# 0.039411f
C265 source.n116 a_n1760_n2088# 0.017655f
C266 source.n117 a_n1760_n2088# 0.132784f
C267 source.t3 a_n1760_n2088# 0.064235f
C268 source.n118 a_n1760_n2088# 0.029558f
C269 source.n119 a_n1760_n2088# 0.02328f
C270 source.n120 a_n1760_n2088# 0.016674f
C271 source.n121 a_n1760_n2088# 0.738314f
C272 source.n122 a_n1760_n2088# 0.031029f
C273 source.n123 a_n1760_n2088# 0.016674f
C274 source.n124 a_n1760_n2088# 0.017655f
C275 source.n125 a_n1760_n2088# 0.039411f
C276 source.n126 a_n1760_n2088# 0.039411f
C277 source.n127 a_n1760_n2088# 0.017655f
C278 source.n128 a_n1760_n2088# 0.016674f
C279 source.n129 a_n1760_n2088# 0.031029f
C280 source.n130 a_n1760_n2088# 0.031029f
C281 source.n131 a_n1760_n2088# 0.016674f
C282 source.n132 a_n1760_n2088# 0.017655f
C283 source.n133 a_n1760_n2088# 0.039411f
C284 source.n134 a_n1760_n2088# 0.085318f
C285 source.n135 a_n1760_n2088# 0.017655f
C286 source.n136 a_n1760_n2088# 0.016674f
C287 source.n137 a_n1760_n2088# 0.071723f
C288 source.n138 a_n1760_n2088# 0.047739f
C289 source.n139 a_n1760_n2088# 1.14244f
C290 source.n140 a_n1760_n2088# 0.043614f
C291 source.n141 a_n1760_n2088# 0.031029f
C292 source.n142 a_n1760_n2088# 0.016674f
C293 source.n143 a_n1760_n2088# 0.039411f
C294 source.n144 a_n1760_n2088# 0.017655f
C295 source.n145 a_n1760_n2088# 0.031029f
C296 source.n146 a_n1760_n2088# 0.016674f
C297 source.n147 a_n1760_n2088# 0.039411f
C298 source.n148 a_n1760_n2088# 0.017655f
C299 source.n149 a_n1760_n2088# 0.132784f
C300 source.t23 a_n1760_n2088# 0.064235f
C301 source.n150 a_n1760_n2088# 0.029558f
C302 source.n151 a_n1760_n2088# 0.02328f
C303 source.n152 a_n1760_n2088# 0.016674f
C304 source.n153 a_n1760_n2088# 0.738314f
C305 source.n154 a_n1760_n2088# 0.031029f
C306 source.n155 a_n1760_n2088# 0.016674f
C307 source.n156 a_n1760_n2088# 0.017655f
C308 source.n157 a_n1760_n2088# 0.039411f
C309 source.n158 a_n1760_n2088# 0.039411f
C310 source.n159 a_n1760_n2088# 0.017655f
C311 source.n160 a_n1760_n2088# 0.016674f
C312 source.n161 a_n1760_n2088# 0.031029f
C313 source.n162 a_n1760_n2088# 0.031029f
C314 source.n163 a_n1760_n2088# 0.016674f
C315 source.n164 a_n1760_n2088# 0.017655f
C316 source.n165 a_n1760_n2088# 0.039411f
C317 source.n166 a_n1760_n2088# 0.085318f
C318 source.n167 a_n1760_n2088# 0.017655f
C319 source.n168 a_n1760_n2088# 0.016674f
C320 source.n169 a_n1760_n2088# 0.071723f
C321 source.n170 a_n1760_n2088# 0.047739f
C322 source.n171 a_n1760_n2088# 1.14244f
C323 source.t24 a_n1760_n2088# 0.147122f
C324 source.t28 a_n1760_n2088# 0.147122f
C325 source.n172 a_n1760_n2088# 1.14579f
C326 source.n173 a_n1760_n2088# 0.390862f
C327 source.t19 a_n1760_n2088# 0.147122f
C328 source.t17 a_n1760_n2088# 0.147122f
C329 source.n174 a_n1760_n2088# 1.14579f
C330 source.n175 a_n1760_n2088# 0.390862f
C331 source.t22 a_n1760_n2088# 0.147122f
C332 source.t29 a_n1760_n2088# 0.147122f
C333 source.n176 a_n1760_n2088# 1.14579f
C334 source.n177 a_n1760_n2088# 0.390862f
C335 source.n178 a_n1760_n2088# 0.043614f
C336 source.n179 a_n1760_n2088# 0.031029f
C337 source.n180 a_n1760_n2088# 0.016674f
C338 source.n181 a_n1760_n2088# 0.039411f
C339 source.n182 a_n1760_n2088# 0.017655f
C340 source.n183 a_n1760_n2088# 0.031029f
C341 source.n184 a_n1760_n2088# 0.016674f
C342 source.n185 a_n1760_n2088# 0.039411f
C343 source.n186 a_n1760_n2088# 0.017655f
C344 source.n187 a_n1760_n2088# 0.132784f
C345 source.t18 a_n1760_n2088# 0.064235f
C346 source.n188 a_n1760_n2088# 0.029558f
C347 source.n189 a_n1760_n2088# 0.02328f
C348 source.n190 a_n1760_n2088# 0.016674f
C349 source.n191 a_n1760_n2088# 0.738314f
C350 source.n192 a_n1760_n2088# 0.031029f
C351 source.n193 a_n1760_n2088# 0.016674f
C352 source.n194 a_n1760_n2088# 0.017655f
C353 source.n195 a_n1760_n2088# 0.039411f
C354 source.n196 a_n1760_n2088# 0.039411f
C355 source.n197 a_n1760_n2088# 0.017655f
C356 source.n198 a_n1760_n2088# 0.016674f
C357 source.n199 a_n1760_n2088# 0.031029f
C358 source.n200 a_n1760_n2088# 0.031029f
C359 source.n201 a_n1760_n2088# 0.016674f
C360 source.n202 a_n1760_n2088# 0.017655f
C361 source.n203 a_n1760_n2088# 0.039411f
C362 source.n204 a_n1760_n2088# 0.085318f
C363 source.n205 a_n1760_n2088# 0.017655f
C364 source.n206 a_n1760_n2088# 0.016674f
C365 source.n207 a_n1760_n2088# 0.071723f
C366 source.n208 a_n1760_n2088# 0.047739f
C367 source.n209 a_n1760_n2088# 0.123468f
C368 source.n210 a_n1760_n2088# 0.043614f
C369 source.n211 a_n1760_n2088# 0.031029f
C370 source.n212 a_n1760_n2088# 0.016674f
C371 source.n213 a_n1760_n2088# 0.039411f
C372 source.n214 a_n1760_n2088# 0.017655f
C373 source.n215 a_n1760_n2088# 0.031029f
C374 source.n216 a_n1760_n2088# 0.016674f
C375 source.n217 a_n1760_n2088# 0.039411f
C376 source.n218 a_n1760_n2088# 0.017655f
C377 source.n219 a_n1760_n2088# 0.132784f
C378 source.t12 a_n1760_n2088# 0.064235f
C379 source.n220 a_n1760_n2088# 0.029558f
C380 source.n221 a_n1760_n2088# 0.02328f
C381 source.n222 a_n1760_n2088# 0.016674f
C382 source.n223 a_n1760_n2088# 0.738314f
C383 source.n224 a_n1760_n2088# 0.031029f
C384 source.n225 a_n1760_n2088# 0.016674f
C385 source.n226 a_n1760_n2088# 0.017655f
C386 source.n227 a_n1760_n2088# 0.039411f
C387 source.n228 a_n1760_n2088# 0.039411f
C388 source.n229 a_n1760_n2088# 0.017655f
C389 source.n230 a_n1760_n2088# 0.016674f
C390 source.n231 a_n1760_n2088# 0.031029f
C391 source.n232 a_n1760_n2088# 0.031029f
C392 source.n233 a_n1760_n2088# 0.016674f
C393 source.n234 a_n1760_n2088# 0.017655f
C394 source.n235 a_n1760_n2088# 0.039411f
C395 source.n236 a_n1760_n2088# 0.085318f
C396 source.n237 a_n1760_n2088# 0.017655f
C397 source.n238 a_n1760_n2088# 0.016674f
C398 source.n239 a_n1760_n2088# 0.071723f
C399 source.n240 a_n1760_n2088# 0.047739f
C400 source.n241 a_n1760_n2088# 0.123468f
C401 source.t5 a_n1760_n2088# 0.147122f
C402 source.t0 a_n1760_n2088# 0.147122f
C403 source.n242 a_n1760_n2088# 1.14579f
C404 source.n243 a_n1760_n2088# 0.390862f
C405 source.t1 a_n1760_n2088# 0.147122f
C406 source.t10 a_n1760_n2088# 0.147122f
C407 source.n244 a_n1760_n2088# 1.14579f
C408 source.n245 a_n1760_n2088# 0.390862f
C409 source.t13 a_n1760_n2088# 0.147122f
C410 source.t11 a_n1760_n2088# 0.147122f
C411 source.n246 a_n1760_n2088# 1.14579f
C412 source.n247 a_n1760_n2088# 0.390862f
C413 source.n248 a_n1760_n2088# 0.043614f
C414 source.n249 a_n1760_n2088# 0.031029f
C415 source.n250 a_n1760_n2088# 0.016674f
C416 source.n251 a_n1760_n2088# 0.039411f
C417 source.n252 a_n1760_n2088# 0.017655f
C418 source.n253 a_n1760_n2088# 0.031029f
C419 source.n254 a_n1760_n2088# 0.016674f
C420 source.n255 a_n1760_n2088# 0.039411f
C421 source.n256 a_n1760_n2088# 0.017655f
C422 source.n257 a_n1760_n2088# 0.132784f
C423 source.t6 a_n1760_n2088# 0.064235f
C424 source.n258 a_n1760_n2088# 0.029558f
C425 source.n259 a_n1760_n2088# 0.02328f
C426 source.n260 a_n1760_n2088# 0.016674f
C427 source.n261 a_n1760_n2088# 0.738314f
C428 source.n262 a_n1760_n2088# 0.031029f
C429 source.n263 a_n1760_n2088# 0.016674f
C430 source.n264 a_n1760_n2088# 0.017655f
C431 source.n265 a_n1760_n2088# 0.039411f
C432 source.n266 a_n1760_n2088# 0.039411f
C433 source.n267 a_n1760_n2088# 0.017655f
C434 source.n268 a_n1760_n2088# 0.016674f
C435 source.n269 a_n1760_n2088# 0.031029f
C436 source.n270 a_n1760_n2088# 0.031029f
C437 source.n271 a_n1760_n2088# 0.016674f
C438 source.n272 a_n1760_n2088# 0.017655f
C439 source.n273 a_n1760_n2088# 0.039411f
C440 source.n274 a_n1760_n2088# 0.085318f
C441 source.n275 a_n1760_n2088# 0.017655f
C442 source.n276 a_n1760_n2088# 0.016674f
C443 source.n277 a_n1760_n2088# 0.071723f
C444 source.n278 a_n1760_n2088# 0.047739f
C445 source.n279 a_n1760_n2088# 0.295179f
C446 source.n280 a_n1760_n2088# 1.26758f
C447 plus.n0 a_n1760_n2088# 0.053149f
C448 plus.t8 a_n1760_n2088# 0.227147f
C449 plus.t14 a_n1760_n2088# 0.227147f
C450 plus.t9 a_n1760_n2088# 0.227147f
C451 plus.n1 a_n1760_n2088# 0.106995f
C452 plus.n2 a_n1760_n2088# 0.053149f
C453 plus.t0 a_n1760_n2088# 0.227147f
C454 plus.t10 a_n1760_n2088# 0.227147f
C455 plus.n3 a_n1760_n2088# 0.106995f
C456 plus.t4 a_n1760_n2088# 0.233077f
C457 plus.n4 a_n1760_n2088# 0.122374f
C458 plus.t1 a_n1760_n2088# 0.227147f
C459 plus.n5 a_n1760_n2088# 0.106995f
C460 plus.n6 a_n1760_n2088# 0.020253f
C461 plus.n7 a_n1760_n2088# 0.116382f
C462 plus.n8 a_n1760_n2088# 0.053149f
C463 plus.n9 a_n1760_n2088# 0.020253f
C464 plus.n10 a_n1760_n2088# 0.106995f
C465 plus.n11 a_n1760_n2088# 0.018942f
C466 plus.n12 a_n1760_n2088# 0.018942f
C467 plus.n13 a_n1760_n2088# 0.053149f
C468 plus.n14 a_n1760_n2088# 0.053149f
C469 plus.n15 a_n1760_n2088# 0.020253f
C470 plus.n16 a_n1760_n2088# 0.106995f
C471 plus.n17 a_n1760_n2088# 0.020253f
C472 plus.n18 a_n1760_n2088# 0.106995f
C473 plus.t3 a_n1760_n2088# 0.233077f
C474 plus.n19 a_n1760_n2088# 0.1223f
C475 plus.n20 a_n1760_n2088# 0.45104f
C476 plus.n21 a_n1760_n2088# 0.053149f
C477 plus.t15 a_n1760_n2088# 0.233077f
C478 plus.t5 a_n1760_n2088# 0.227147f
C479 plus.t7 a_n1760_n2088# 0.227147f
C480 plus.t13 a_n1760_n2088# 0.227147f
C481 plus.n22 a_n1760_n2088# 0.106995f
C482 plus.n23 a_n1760_n2088# 0.053149f
C483 plus.t12 a_n1760_n2088# 0.227147f
C484 plus.t2 a_n1760_n2088# 0.227147f
C485 plus.n24 a_n1760_n2088# 0.106995f
C486 plus.t11 a_n1760_n2088# 0.233077f
C487 plus.n25 a_n1760_n2088# 0.122374f
C488 plus.t6 a_n1760_n2088# 0.227147f
C489 plus.n26 a_n1760_n2088# 0.106995f
C490 plus.n27 a_n1760_n2088# 0.020253f
C491 plus.n28 a_n1760_n2088# 0.116382f
C492 plus.n29 a_n1760_n2088# 0.053149f
C493 plus.n30 a_n1760_n2088# 0.020253f
C494 plus.n31 a_n1760_n2088# 0.106995f
C495 plus.n32 a_n1760_n2088# 0.018942f
C496 plus.n33 a_n1760_n2088# 0.018942f
C497 plus.n34 a_n1760_n2088# 0.053149f
C498 plus.n35 a_n1760_n2088# 0.053149f
C499 plus.n36 a_n1760_n2088# 0.020253f
C500 plus.n37 a_n1760_n2088# 0.106995f
C501 plus.n38 a_n1760_n2088# 0.020253f
C502 plus.n39 a_n1760_n2088# 0.106995f
C503 plus.n40 a_n1760_n2088# 0.1223f
C504 plus.n41 a_n1760_n2088# 1.33349f
.ends

