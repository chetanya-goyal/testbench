* NGSPICE file created from diffpair75.ext - technology: sky130A

.subckt diffpair75 minus drain_right drain_left source plus
X0 source.t23 minus.t0 drain_right.t3 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X1 a_n2298_n1088# a_n2298_n1088# a_n2298_n1088# a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=3.12 ps=22.24 w=1 l=0.8
X2 drain_left.t11 plus.t0 source.t2 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X3 a_n2298_n1088# a_n2298_n1088# a_n2298_n1088# a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X4 source.t22 minus.t1 drain_right.t2 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X5 source.t21 minus.t2 drain_right.t4 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X6 a_n2298_n1088# a_n2298_n1088# a_n2298_n1088# a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X7 drain_right.t11 minus.t3 source.t20 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X8 drain_left.t10 plus.t1 source.t4 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X9 drain_left.t9 plus.t2 source.t1 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X10 source.t19 minus.t4 drain_right.t8 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X11 drain_right.t9 minus.t5 source.t18 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X12 source.t17 minus.t6 drain_right.t10 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X13 source.t16 minus.t7 drain_right.t1 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X14 a_n2298_n1088# a_n2298_n1088# a_n2298_n1088# a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.8
X15 drain_right.t7 minus.t8 source.t15 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X16 drain_left.t8 plus.t3 source.t3 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X17 drain_left.t7 plus.t4 source.t7 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X18 drain_right.t5 minus.t9 source.t14 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X19 drain_right.t6 minus.t10 source.t13 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X20 source.t9 plus.t5 drain_left.t6 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X21 source.t11 plus.t6 drain_left.t5 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X22 drain_left.t4 plus.t7 source.t0 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X23 drain_right.t0 minus.t11 source.t12 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.8
X24 source.t5 plus.t8 drain_left.t3 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X25 source.t6 plus.t9 drain_left.t2 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
X26 source.t8 plus.t10 drain_left.t1 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.8
X27 source.t10 plus.t11 drain_left.t0 a_n2298_n1088# sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.8
R0 minus.n15 minus.n14 161.3
R1 minus.n13 minus.n0 161.3
R2 minus.n12 minus.n11 161.3
R3 minus.n10 minus.n1 161.3
R4 minus.n6 minus.n5 161.3
R5 minus.n31 minus.n30 161.3
R6 minus.n29 minus.n16 161.3
R7 minus.n28 minus.n27 161.3
R8 minus.n26 minus.n17 161.3
R9 minus.n22 minus.n21 161.3
R10 minus.n4 minus.t5 100.626
R11 minus.n20 minus.t2 100.626
R12 minus.n9 minus.n8 80.6037
R13 minus.n7 minus.n2 80.6037
R14 minus.n25 minus.n24 80.6037
R15 minus.n23 minus.n18 80.6037
R16 minus.n3 minus.t4 79.2293
R17 minus.n7 minus.t3 79.2293
R18 minus.n8 minus.t7 79.2293
R19 minus.n12 minus.t8 79.2293
R20 minus.n14 minus.t6 79.2293
R21 minus.n19 minus.t10 79.2293
R22 minus.n23 minus.t1 79.2293
R23 minus.n24 minus.t9 79.2293
R24 minus.n28 minus.t0 79.2293
R25 minus.n30 minus.t11 79.2293
R26 minus.n8 minus.n7 48.2005
R27 minus.n24 minus.n23 48.2005
R28 minus.n5 minus.n4 44.853
R29 minus.n21 minus.n20 44.853
R30 minus.n7 minus.n6 41.6278
R31 minus.n8 minus.n1 41.6278
R32 minus.n23 minus.n22 41.6278
R33 minus.n24 minus.n17 41.6278
R34 minus.n32 minus.n15 29.6937
R35 minus.n14 minus.n13 25.5611
R36 minus.n30 minus.n29 25.5611
R37 minus.n13 minus.n12 22.6399
R38 minus.n29 minus.n28 22.6399
R39 minus.n4 minus.n3 20.5405
R40 minus.n20 minus.n19 20.5405
R41 minus.n32 minus.n31 6.70126
R42 minus.n6 minus.n3 6.57323
R43 minus.n12 minus.n1 6.57323
R44 minus.n22 minus.n19 6.57323
R45 minus.n28 minus.n17 6.57323
R46 minus.n9 minus.n2 0.380177
R47 minus.n25 minus.n18 0.380177
R48 minus.n10 minus.n9 0.285035
R49 minus.n5 minus.n2 0.285035
R50 minus.n21 minus.n18 0.285035
R51 minus.n26 minus.n25 0.285035
R52 minus.n15 minus.n0 0.189894
R53 minus.n11 minus.n0 0.189894
R54 minus.n11 minus.n10 0.189894
R55 minus.n27 minus.n26 0.189894
R56 minus.n27 minus.n16 0.189894
R57 minus.n31 minus.n16 0.189894
R58 minus minus.n32 0.188
R59 drain_right.n6 drain_right.n4 241.107
R60 drain_right.n3 drain_right.n2 241.05
R61 drain_right.n3 drain_right.n0 241.05
R62 drain_right.n6 drain_right.n5 240.132
R63 drain_right.n8 drain_right.n7 240.132
R64 drain_right.n3 drain_right.n1 240.131
R65 drain_right drain_right.n3 23.3512
R66 drain_right.n1 drain_right.t2 19.8005
R67 drain_right.n1 drain_right.t5 19.8005
R68 drain_right.n2 drain_right.t3 19.8005
R69 drain_right.n2 drain_right.t0 19.8005
R70 drain_right.n0 drain_right.t4 19.8005
R71 drain_right.n0 drain_right.t6 19.8005
R72 drain_right.n4 drain_right.t8 19.8005
R73 drain_right.n4 drain_right.t9 19.8005
R74 drain_right.n5 drain_right.t1 19.8005
R75 drain_right.n5 drain_right.t11 19.8005
R76 drain_right.n7 drain_right.t10 19.8005
R77 drain_right.n7 drain_right.t7 19.8005
R78 drain_right drain_right.n8 6.62735
R79 drain_right.n8 drain_right.n6 0.974638
R80 source.n0 source.t3 243.255
R81 source.n5 source.t6 243.255
R82 source.n6 source.t18 243.255
R83 source.n11 source.t17 243.255
R84 source.n23 source.t12 243.254
R85 source.n18 source.t21 243.254
R86 source.n17 source.t4 243.254
R87 source.n12 source.t10 243.254
R88 source.n2 source.n1 223.454
R89 source.n4 source.n3 223.454
R90 source.n8 source.n7 223.454
R91 source.n10 source.n9 223.454
R92 source.n22 source.n21 223.453
R93 source.n20 source.n19 223.453
R94 source.n16 source.n15 223.453
R95 source.n14 source.n13 223.453
R96 source.n21 source.t14 19.8005
R97 source.n21 source.t23 19.8005
R98 source.n19 source.t13 19.8005
R99 source.n19 source.t22 19.8005
R100 source.n15 source.t1 19.8005
R101 source.n15 source.t5 19.8005
R102 source.n13 source.t2 19.8005
R103 source.n13 source.t8 19.8005
R104 source.n1 source.t7 19.8005
R105 source.n1 source.t11 19.8005
R106 source.n3 source.t0 19.8005
R107 source.n3 source.t9 19.8005
R108 source.n7 source.t20 19.8005
R109 source.n7 source.t19 19.8005
R110 source.n9 source.t15 19.8005
R111 source.n9 source.t16 19.8005
R112 source.n12 source.n11 13.9285
R113 source.n24 source.n0 8.17853
R114 source.n24 source.n23 5.7505
R115 source.n11 source.n10 0.974638
R116 source.n10 source.n8 0.974638
R117 source.n8 source.n6 0.974638
R118 source.n5 source.n4 0.974638
R119 source.n4 source.n2 0.974638
R120 source.n2 source.n0 0.974638
R121 source.n14 source.n12 0.974638
R122 source.n16 source.n14 0.974638
R123 source.n17 source.n16 0.974638
R124 source.n20 source.n18 0.974638
R125 source.n22 source.n20 0.974638
R126 source.n23 source.n22 0.974638
R127 source.n6 source.n5 0.470328
R128 source.n18 source.n17 0.470328
R129 source source.n24 0.188
R130 plus.n6 plus.n3 161.3
R131 plus.n11 plus.n10 161.3
R132 plus.n12 plus.n1 161.3
R133 plus.n13 plus.n0 161.3
R134 plus.n15 plus.n14 161.3
R135 plus.n22 plus.n19 161.3
R136 plus.n27 plus.n26 161.3
R137 plus.n28 plus.n17 161.3
R138 plus.n29 plus.n16 161.3
R139 plus.n31 plus.n30 161.3
R140 plus.n4 plus.t9 100.626
R141 plus.n20 plus.t1 100.626
R142 plus.n8 plus.n7 80.6037
R143 plus.n9 plus.n2 80.6037
R144 plus.n24 plus.n23 80.6037
R145 plus.n25 plus.n18 80.6037
R146 plus.n14 plus.t3 79.2293
R147 plus.n12 plus.t6 79.2293
R148 plus.n2 plus.t4 79.2293
R149 plus.n7 plus.t5 79.2293
R150 plus.n5 plus.t7 79.2293
R151 plus.n30 plus.t11 79.2293
R152 plus.n28 plus.t0 79.2293
R153 plus.n18 plus.t10 79.2293
R154 plus.n23 plus.t2 79.2293
R155 plus.n21 plus.t8 79.2293
R156 plus.n7 plus.n2 48.2005
R157 plus.n23 plus.n18 48.2005
R158 plus.n4 plus.n3 44.853
R159 plus.n20 plus.n19 44.853
R160 plus.n11 plus.n2 41.6278
R161 plus.n7 plus.n6 41.6278
R162 plus.n27 plus.n18 41.6278
R163 plus.n23 plus.n22 41.6278
R164 plus plus.n31 27.7414
R165 plus.n14 plus.n13 25.5611
R166 plus.n30 plus.n29 25.5611
R167 plus.n13 plus.n12 22.6399
R168 plus.n29 plus.n28 22.6399
R169 plus.n5 plus.n4 20.5405
R170 plus.n21 plus.n20 20.5405
R171 plus plus.n15 8.17853
R172 plus.n12 plus.n11 6.57323
R173 plus.n6 plus.n5 6.57323
R174 plus.n28 plus.n27 6.57323
R175 plus.n22 plus.n21 6.57323
R176 plus.n9 plus.n8 0.380177
R177 plus.n25 plus.n24 0.380177
R178 plus.n8 plus.n3 0.285035
R179 plus.n10 plus.n9 0.285035
R180 plus.n26 plus.n25 0.285035
R181 plus.n24 plus.n19 0.285035
R182 plus.n10 plus.n1 0.189894
R183 plus.n1 plus.n0 0.189894
R184 plus.n15 plus.n0 0.189894
R185 plus.n31 plus.n16 0.189894
R186 plus.n17 plus.n16 0.189894
R187 plus.n26 plus.n17 0.189894
R188 drain_left.n6 drain_left.n4 241.107
R189 drain_left.n3 drain_left.n2 241.05
R190 drain_left.n3 drain_left.n0 241.05
R191 drain_left.n8 drain_left.n7 240.132
R192 drain_left.n6 drain_left.n5 240.132
R193 drain_left.n3 drain_left.n1 240.131
R194 drain_left drain_left.n3 23.9044
R195 drain_left.n1 drain_left.t1 19.8005
R196 drain_left.n1 drain_left.t9 19.8005
R197 drain_left.n2 drain_left.t3 19.8005
R198 drain_left.n2 drain_left.t10 19.8005
R199 drain_left.n0 drain_left.t0 19.8005
R200 drain_left.n0 drain_left.t11 19.8005
R201 drain_left.n7 drain_left.t5 19.8005
R202 drain_left.n7 drain_left.t8 19.8005
R203 drain_left.n5 drain_left.t6 19.8005
R204 drain_left.n5 drain_left.t7 19.8005
R205 drain_left.n4 drain_left.t2 19.8005
R206 drain_left.n4 drain_left.t4 19.8005
R207 drain_left drain_left.n8 6.62735
R208 drain_left.n8 drain_left.n6 0.974638
C0 source drain_left 3.91551f
C1 drain_left plus 1.39493f
C2 source drain_right 3.91805f
C3 drain_right plus 0.39034f
C4 minus drain_left 0.179384f
C5 source plus 1.76774f
C6 minus drain_right 1.16881f
C7 drain_left drain_right 1.16235f
C8 minus source 1.75387f
C9 minus plus 3.9779f
C10 drain_right a_n2298_n1088# 3.81724f
C11 drain_left a_n2298_n1088# 4.09981f
C12 source a_n2298_n1088# 2.638721f
C13 minus a_n2298_n1088# 8.149334f
C14 plus a_n2298_n1088# 8.753612f
C15 drain_left.t0 a_n2298_n1088# 0.015159f
C16 drain_left.t11 a_n2298_n1088# 0.015159f
C17 drain_left.n0 a_n2298_n1088# 0.059894f
C18 drain_left.t1 a_n2298_n1088# 0.015159f
C19 drain_left.t9 a_n2298_n1088# 0.015159f
C20 drain_left.n1 a_n2298_n1088# 0.058905f
C21 drain_left.t3 a_n2298_n1088# 0.015159f
C22 drain_left.t10 a_n2298_n1088# 0.015159f
C23 drain_left.n2 a_n2298_n1088# 0.059894f
C24 drain_left.n3 a_n2298_n1088# 1.33515f
C25 drain_left.t2 a_n2298_n1088# 0.015159f
C26 drain_left.t4 a_n2298_n1088# 0.015159f
C27 drain_left.n4 a_n2298_n1088# 0.059965f
C28 drain_left.t6 a_n2298_n1088# 0.015159f
C29 drain_left.t7 a_n2298_n1088# 0.015159f
C30 drain_left.n5 a_n2298_n1088# 0.058905f
C31 drain_left.n6 a_n2298_n1088# 0.515833f
C32 drain_left.t5 a_n2298_n1088# 0.015159f
C33 drain_left.t8 a_n2298_n1088# 0.015159f
C34 drain_left.n7 a_n2298_n1088# 0.058905f
C35 drain_left.n8 a_n2298_n1088# 0.426601f
C36 plus.n0 a_n2298_n1088# 0.026284f
C37 plus.t3 a_n2298_n1088# 0.071304f
C38 plus.t6 a_n2298_n1088# 0.071304f
C39 plus.n1 a_n2298_n1088# 0.026284f
C40 plus.t4 a_n2298_n1088# 0.071304f
C41 plus.n2 a_n2298_n1088# 0.075825f
C42 plus.n3 a_n2298_n1088# 0.120665f
C43 plus.t5 a_n2298_n1088# 0.071304f
C44 plus.t7 a_n2298_n1088# 0.071304f
C45 plus.t9 a_n2298_n1088# 0.086173f
C46 plus.n4 a_n2298_n1088# 0.057678f
C47 plus.n5 a_n2298_n1088# 0.07053f
C48 plus.n6 a_n2298_n1088# 0.005964f
C49 plus.n7 a_n2298_n1088# 0.075825f
C50 plus.n8 a_n2298_n1088# 0.04378f
C51 plus.n9 a_n2298_n1088# 0.04378f
C52 plus.n10 a_n2298_n1088# 0.035073f
C53 plus.n11 a_n2298_n1088# 0.005964f
C54 plus.n12 a_n2298_n1088# 0.068483f
C55 plus.n13 a_n2298_n1088# 0.005964f
C56 plus.n14 a_n2298_n1088# 0.068078f
C57 plus.n15 a_n2298_n1088# 0.193226f
C58 plus.n16 a_n2298_n1088# 0.026284f
C59 plus.t11 a_n2298_n1088# 0.071304f
C60 plus.n17 a_n2298_n1088# 0.026284f
C61 plus.t0 a_n2298_n1088# 0.071304f
C62 plus.t10 a_n2298_n1088# 0.071304f
C63 plus.n18 a_n2298_n1088# 0.075825f
C64 plus.n19 a_n2298_n1088# 0.120665f
C65 plus.t2 a_n2298_n1088# 0.071304f
C66 plus.t1 a_n2298_n1088# 0.086173f
C67 plus.n20 a_n2298_n1088# 0.057678f
C68 plus.t8 a_n2298_n1088# 0.071304f
C69 plus.n21 a_n2298_n1088# 0.07053f
C70 plus.n22 a_n2298_n1088# 0.005964f
C71 plus.n23 a_n2298_n1088# 0.075825f
C72 plus.n24 a_n2298_n1088# 0.04378f
C73 plus.n25 a_n2298_n1088# 0.04378f
C74 plus.n26 a_n2298_n1088# 0.035073f
C75 plus.n27 a_n2298_n1088# 0.005964f
C76 plus.n28 a_n2298_n1088# 0.068483f
C77 plus.n29 a_n2298_n1088# 0.005964f
C78 plus.n30 a_n2298_n1088# 0.068078f
C79 plus.n31 a_n2298_n1088# 0.654038f
C80 source.t3 a_n2298_n1088# 0.102948f
C81 source.n0 a_n2298_n1088# 0.500045f
C82 source.t7 a_n2298_n1088# 0.018496f
C83 source.t11 a_n2298_n1088# 0.018496f
C84 source.n1 a_n2298_n1088# 0.059986f
C85 source.n2 a_n2298_n1088# 0.290692f
C86 source.t0 a_n2298_n1088# 0.018496f
C87 source.t9 a_n2298_n1088# 0.018496f
C88 source.n3 a_n2298_n1088# 0.059986f
C89 source.n4 a_n2298_n1088# 0.290692f
C90 source.t6 a_n2298_n1088# 0.102948f
C91 source.n5 a_n2298_n1088# 0.26014f
C92 source.t18 a_n2298_n1088# 0.102948f
C93 source.n6 a_n2298_n1088# 0.26014f
C94 source.t20 a_n2298_n1088# 0.018496f
C95 source.t19 a_n2298_n1088# 0.018496f
C96 source.n7 a_n2298_n1088# 0.059986f
C97 source.n8 a_n2298_n1088# 0.290692f
C98 source.t15 a_n2298_n1088# 0.018496f
C99 source.t16 a_n2298_n1088# 0.018496f
C100 source.n9 a_n2298_n1088# 0.059986f
C101 source.n10 a_n2298_n1088# 0.290692f
C102 source.t17 a_n2298_n1088# 0.102948f
C103 source.n11 a_n2298_n1088# 0.694612f
C104 source.t10 a_n2298_n1088# 0.102947f
C105 source.n12 a_n2298_n1088# 0.694612f
C106 source.t2 a_n2298_n1088# 0.018496f
C107 source.t8 a_n2298_n1088# 0.018496f
C108 source.n13 a_n2298_n1088# 0.059986f
C109 source.n14 a_n2298_n1088# 0.290692f
C110 source.t1 a_n2298_n1088# 0.018496f
C111 source.t5 a_n2298_n1088# 0.018496f
C112 source.n15 a_n2298_n1088# 0.059986f
C113 source.n16 a_n2298_n1088# 0.290692f
C114 source.t4 a_n2298_n1088# 0.102947f
C115 source.n17 a_n2298_n1088# 0.26014f
C116 source.t21 a_n2298_n1088# 0.102947f
C117 source.n18 a_n2298_n1088# 0.26014f
C118 source.t13 a_n2298_n1088# 0.018496f
C119 source.t22 a_n2298_n1088# 0.018496f
C120 source.n19 a_n2298_n1088# 0.059986f
C121 source.n20 a_n2298_n1088# 0.290692f
C122 source.t14 a_n2298_n1088# 0.018496f
C123 source.t23 a_n2298_n1088# 0.018496f
C124 source.n21 a_n2298_n1088# 0.059986f
C125 source.n22 a_n2298_n1088# 0.290692f
C126 source.t12 a_n2298_n1088# 0.102947f
C127 source.n23 a_n2298_n1088# 0.417887f
C128 source.n24 a_n2298_n1088# 0.48794f
C129 drain_right.t4 a_n2298_n1088# 0.015457f
C130 drain_right.t6 a_n2298_n1088# 0.015457f
C131 drain_right.n0 a_n2298_n1088# 0.061069f
C132 drain_right.t2 a_n2298_n1088# 0.015457f
C133 drain_right.t5 a_n2298_n1088# 0.015457f
C134 drain_right.n1 a_n2298_n1088# 0.060061f
C135 drain_right.t3 a_n2298_n1088# 0.015457f
C136 drain_right.t0 a_n2298_n1088# 0.015457f
C137 drain_right.n2 a_n2298_n1088# 0.061069f
C138 drain_right.n3 a_n2298_n1088# 1.32365f
C139 drain_right.t8 a_n2298_n1088# 0.015457f
C140 drain_right.t9 a_n2298_n1088# 0.015457f
C141 drain_right.n4 a_n2298_n1088# 0.061141f
C142 drain_right.t1 a_n2298_n1088# 0.015457f
C143 drain_right.t11 a_n2298_n1088# 0.015457f
C144 drain_right.n5 a_n2298_n1088# 0.060061f
C145 drain_right.n6 a_n2298_n1088# 0.525953f
C146 drain_right.t10 a_n2298_n1088# 0.015457f
C147 drain_right.t7 a_n2298_n1088# 0.015457f
C148 drain_right.n7 a_n2298_n1088# 0.060061f
C149 drain_right.n8 a_n2298_n1088# 0.434971f
C150 minus.n0 a_n2298_n1088# 0.025939f
C151 minus.n1 a_n2298_n1088# 0.005886f
C152 minus.t8 a_n2298_n1088# 0.070368f
C153 minus.n2 a_n2298_n1088# 0.043206f
C154 minus.t4 a_n2298_n1088# 0.070368f
C155 minus.n3 a_n2298_n1088# 0.069605f
C156 minus.t5 a_n2298_n1088# 0.085043f
C157 minus.n4 a_n2298_n1088# 0.056921f
C158 minus.n5 a_n2298_n1088# 0.119082f
C159 minus.n6 a_n2298_n1088# 0.005886f
C160 minus.t3 a_n2298_n1088# 0.070368f
C161 minus.n7 a_n2298_n1088# 0.07483f
C162 minus.t7 a_n2298_n1088# 0.070368f
C163 minus.n8 a_n2298_n1088# 0.07483f
C164 minus.n9 a_n2298_n1088# 0.043206f
C165 minus.n10 a_n2298_n1088# 0.034613f
C166 minus.n11 a_n2298_n1088# 0.025939f
C167 minus.n12 a_n2298_n1088# 0.067585f
C168 minus.n13 a_n2298_n1088# 0.005886f
C169 minus.t6 a_n2298_n1088# 0.070368f
C170 minus.n14 a_n2298_n1088# 0.067185f
C171 minus.n15 a_n2298_n1088# 0.667951f
C172 minus.n16 a_n2298_n1088# 0.025939f
C173 minus.n17 a_n2298_n1088# 0.005886f
C174 minus.n18 a_n2298_n1088# 0.043206f
C175 minus.t10 a_n2298_n1088# 0.070368f
C176 minus.n19 a_n2298_n1088# 0.069605f
C177 minus.t2 a_n2298_n1088# 0.085043f
C178 minus.n20 a_n2298_n1088# 0.056921f
C179 minus.n21 a_n2298_n1088# 0.119082f
C180 minus.n22 a_n2298_n1088# 0.005886f
C181 minus.t1 a_n2298_n1088# 0.070368f
C182 minus.n23 a_n2298_n1088# 0.07483f
C183 minus.t9 a_n2298_n1088# 0.070368f
C184 minus.n24 a_n2298_n1088# 0.07483f
C185 minus.n25 a_n2298_n1088# 0.043206f
C186 minus.n26 a_n2298_n1088# 0.034613f
C187 minus.n27 a_n2298_n1088# 0.025939f
C188 minus.t0 a_n2298_n1088# 0.070368f
C189 minus.n28 a_n2298_n1088# 0.067585f
C190 minus.n29 a_n2298_n1088# 0.005886f
C191 minus.t11 a_n2298_n1088# 0.070368f
C192 minus.n30 a_n2298_n1088# 0.067185f
C193 minus.n31 a_n2298_n1088# 0.181771f
C194 minus.n32 a_n2298_n1088# 0.818272f
.ends

