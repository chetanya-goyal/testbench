* NGSPICE file created from diffpair191.ext - technology: sky130A

.subckt diffpair191 minus drain_right drain_left source plus
X0 drain_right.t3 minus.t0 source.t4 a_n1094_n1492# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X1 a_n1094_n1492# a_n1094_n1492# a_n1094_n1492# a_n1094_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.3
X2 source.t5 minus.t1 drain_right.t2 a_n1094_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X3 a_n1094_n1492# a_n1094_n1492# a_n1094_n1492# a_n1094_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X4 source.t3 plus.t0 drain_left.t3 a_n1094_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X5 drain_right.t1 minus.t2 source.t6 a_n1094_n1492# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X6 a_n1094_n1492# a_n1094_n1492# a_n1094_n1492# a_n1094_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X7 source.t2 plus.t1 drain_left.t2 a_n1094_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
X8 drain_left.t1 plus.t2 source.t1 a_n1094_n1492# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X9 a_n1094_n1492# a_n1094_n1492# a_n1094_n1492# a_n1094_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.3
X10 drain_left.t0 plus.t3 source.t0 a_n1094_n1492# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.3
X11 source.t7 minus.t3 drain_right.t0 a_n1094_n1492# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.3
R0 minus.n0 minus.t1 391.442
R1 minus.n0 minus.t0 391.442
R2 minus.n1 minus.t2 391.442
R3 minus.n1 minus.t3 391.442
R4 minus.n2 minus.n0 187.77
R5 minus.n2 minus.n1 167.809
R6 minus minus.n2 0.188
R7 source.n0 source.t0 69.6943
R8 source.n1 source.t2 69.6943
R9 source.n2 source.t4 69.6943
R10 source.n3 source.t5 69.6943
R11 source.n7 source.t6 69.6942
R12 source.n6 source.t7 69.6942
R13 source.n5 source.t1 69.6942
R14 source.n4 source.t3 69.6942
R15 source.n4 source.n3 15.0278
R16 source.n8 source.n0 9.49332
R17 source.n8 source.n7 5.53498
R18 source.n3 source.n2 0.543603
R19 source.n1 source.n0 0.543603
R20 source.n5 source.n4 0.543603
R21 source.n7 source.n6 0.543603
R22 source.n2 source.n1 0.470328
R23 source.n6 source.n5 0.470328
R24 source source.n8 0.188
R25 drain_right drain_right.n0 100.87
R26 drain_right drain_right.n1 85.9689
R27 drain_right.n0 drain_right.t0 6.6005
R28 drain_right.n0 drain_right.t1 6.6005
R29 drain_right.n1 drain_right.t2 6.6005
R30 drain_right.n1 drain_right.t3 6.6005
R31 plus.n0 plus.t1 391.442
R32 plus.n0 plus.t3 391.442
R33 plus.n1 plus.t2 391.442
R34 plus.n1 plus.t0 391.442
R35 plus plus.n1 185.06
R36 plus plus.n0 170.042
R37 drain_left drain_left.n0 101.422
R38 drain_left drain_left.n1 85.9689
R39 drain_left.n0 drain_left.t3 6.6005
R40 drain_left.n0 drain_left.t1 6.6005
R41 drain_left.n1 drain_left.t2 6.6005
R42 drain_left.n1 drain_left.t0 6.6005
C0 drain_left source 3.3878f
C1 drain_left minus 0.1762f
C2 source drain_right 3.38634f
C3 minus drain_right 0.732285f
C4 source minus 0.667038f
C5 plus drain_left 0.833259f
C6 plus drain_right 0.260363f
C7 plus source 0.681036f
C8 plus minus 2.84821f
C9 drain_left drain_right 0.477436f
C10 drain_right a_n1094_n1492# 3.87053f
C11 drain_left a_n1094_n1492# 3.99988f
C12 source a_n1094_n1492# 3.385202f
C13 minus a_n1094_n1492# 3.456714f
C14 plus a_n1094_n1492# 5.26674f
C15 drain_left.t3 a_n1094_n1492# 0.056278f
C16 drain_left.t1 a_n1094_n1492# 0.056278f
C17 drain_left.n0 a_n1094_n1492# 0.542948f
C18 drain_left.t2 a_n1094_n1492# 0.056278f
C19 drain_left.t0 a_n1094_n1492# 0.056278f
C20 drain_left.n1 a_n1094_n1492# 0.440485f
C21 plus.t1 a_n1094_n1492# 0.11181f
C22 plus.t3 a_n1094_n1492# 0.11181f
C23 plus.n0 a_n1094_n1492# 0.144408f
C24 plus.t0 a_n1094_n1492# 0.11181f
C25 plus.t2 a_n1094_n1492# 0.11181f
C26 plus.n1 a_n1094_n1492# 0.231569f
C27 drain_right.t0 a_n1094_n1492# 0.057858f
C28 drain_right.t1 a_n1094_n1492# 0.057858f
C29 drain_right.n0 a_n1094_n1492# 0.545129f
C30 drain_right.t2 a_n1094_n1492# 0.057858f
C31 drain_right.t3 a_n1094_n1492# 0.057858f
C32 drain_right.n1 a_n1094_n1492# 0.452854f
C33 source.t0 a_n1094_n1492# 0.367347f
C34 source.n0 a_n1094_n1492# 0.501986f
C35 source.t2 a_n1094_n1492# 0.367347f
C36 source.n1 a_n1094_n1492# 0.257262f
C37 source.t4 a_n1094_n1492# 0.367347f
C38 source.n2 a_n1094_n1492# 0.257262f
C39 source.t5 a_n1094_n1492# 0.367347f
C40 source.n3 a_n1094_n1492# 0.696874f
C41 source.t3 a_n1094_n1492# 0.367345f
C42 source.n4 a_n1094_n1492# 0.696876f
C43 source.t1 a_n1094_n1492# 0.367345f
C44 source.n5 a_n1094_n1492# 0.257264f
C45 source.t7 a_n1094_n1492# 0.367345f
C46 source.n6 a_n1094_n1492# 0.257264f
C47 source.t6 a_n1094_n1492# 0.367345f
C48 source.n7 a_n1094_n1492# 0.362602f
C49 source.n8 a_n1094_n1492# 0.542434f
C50 minus.t1 a_n1094_n1492# 0.108667f
C51 minus.t0 a_n1094_n1492# 0.108667f
C52 minus.n0 a_n1094_n1492# 0.240705f
C53 minus.t3 a_n1094_n1492# 0.108667f
C54 minus.t2 a_n1094_n1492# 0.108667f
C55 minus.n1 a_n1094_n1492# 0.135129f
C56 minus.n2 a_n1094_n1492# 1.96394f
.ends

