* NGSPICE file created from diffpair167.ext - technology: sky130A

.subckt diffpair167 minus drain_right drain_left source plus
X0 source.t31 plus.t0 drain_left.t14 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X1 drain_right.t15 minus.t0 source.t3 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X2 a_n1886_n1488# a_n1886_n1488# a_n1886_n1488# a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=11.4 ps=55.6 w=3 l=0.15
X3 drain_right.t14 minus.t1 source.t7 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X4 source.t30 plus.t1 drain_left.t13 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X5 source.t9 minus.t2 drain_right.t13 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X6 drain_left.t12 plus.t2 source.t29 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X7 drain_right.t12 minus.t3 source.t0 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X8 drain_left.t11 plus.t3 source.t28 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X9 source.t13 minus.t4 drain_right.t11 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X10 a_n1886_n1488# a_n1886_n1488# a_n1886_n1488# a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X11 a_n1886_n1488# a_n1886_n1488# a_n1886_n1488# a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X12 source.t1 minus.t5 drain_right.t10 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X13 source.t11 minus.t6 drain_right.t9 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X14 source.t27 plus.t4 drain_left.t6 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X15 drain_right.t8 minus.t7 source.t15 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X16 drain_right.t7 minus.t8 source.t2 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X17 source.t14 minus.t9 drain_right.t6 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X18 drain_left.t9 plus.t5 source.t26 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X19 source.t25 plus.t6 drain_left.t15 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X20 drain_left.t5 plus.t7 source.t24 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
X21 source.t23 plus.t8 drain_left.t10 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X22 drain_right.t5 minus.t10 source.t4 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X23 drain_right.t4 minus.t11 source.t8 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X24 a_n1886_n1488# a_n1886_n1488# a_n1886_n1488# a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X25 source.t10 minus.t12 drain_right.t3 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
X26 drain_left.t7 plus.t9 source.t22 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X27 source.t5 minus.t13 drain_right.t2 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X28 drain_right.t1 minus.t14 source.t12 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X29 source.t21 plus.t10 drain_left.t0 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X30 source.t20 plus.t11 drain_left.t4 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X31 drain_left.t1 plus.t12 source.t19 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X32 drain_left.t8 plus.t13 source.t18 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X33 drain_left.t2 plus.t14 source.t17 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X34 source.t6 minus.t15 drain_right.t0 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
X35 source.t16 plus.t15 drain_left.t3 a_n1886_n1488# sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.15
R0 plus.n5 plus.t8 731.034
R1 plus.n21 plus.t7 731.034
R2 plus.n28 plus.t2 731.034
R3 plus.n44 plus.t6 731.034
R4 plus.n6 plus.t14 690.867
R5 plus.n3 plus.t11 690.867
R6 plus.n12 plus.t9 690.867
R7 plus.n14 plus.t15 690.867
R8 plus.n1 plus.t13 690.867
R9 plus.n20 plus.t10 690.867
R10 plus.n29 plus.t1 690.867
R11 plus.n26 plus.t5 690.867
R12 plus.n35 plus.t4 690.867
R13 plus.n37 plus.t3 690.867
R14 plus.n24 plus.t0 690.867
R15 plus.n43 plus.t12 690.867
R16 plus.n5 plus.n4 161.489
R17 plus.n28 plus.n27 161.489
R18 plus.n7 plus.n4 161.3
R19 plus.n9 plus.n8 161.3
R20 plus.n11 plus.n10 161.3
R21 plus.n13 plus.n2 161.3
R22 plus.n16 plus.n15 161.3
R23 plus.n18 plus.n17 161.3
R24 plus.n19 plus.n0 161.3
R25 plus.n22 plus.n21 161.3
R26 plus.n30 plus.n27 161.3
R27 plus.n32 plus.n31 161.3
R28 plus.n34 plus.n33 161.3
R29 plus.n36 plus.n25 161.3
R30 plus.n39 plus.n38 161.3
R31 plus.n41 plus.n40 161.3
R32 plus.n42 plus.n23 161.3
R33 plus.n45 plus.n44 161.3
R34 plus.n8 plus.n7 73.0308
R35 plus.n19 plus.n18 73.0308
R36 plus.n42 plus.n41 73.0308
R37 plus.n31 plus.n30 73.0308
R38 plus.n11 plus.n3 69.3793
R39 plus.n15 plus.n1 69.3793
R40 plus.n38 plus.n24 69.3793
R41 plus.n34 plus.n26 69.3793
R42 plus.n6 plus.n5 54.7732
R43 plus.n21 plus.n20 54.7732
R44 plus.n44 plus.n43 54.7732
R45 plus.n29 plus.n28 54.7732
R46 plus.n13 plus.n12 47.4702
R47 plus.n14 plus.n13 47.4702
R48 plus.n37 plus.n36 47.4702
R49 plus.n36 plus.n35 47.4702
R50 plus plus.n45 26.7414
R51 plus.n12 plus.n11 25.5611
R52 plus.n15 plus.n14 25.5611
R53 plus.n38 plus.n37 25.5611
R54 plus.n35 plus.n34 25.5611
R55 plus.n7 plus.n6 18.2581
R56 plus.n20 plus.n19 18.2581
R57 plus.n43 plus.n42 18.2581
R58 plus.n30 plus.n29 18.2581
R59 plus plus.n22 8.73914
R60 plus.n8 plus.n3 3.65202
R61 plus.n18 plus.n1 3.65202
R62 plus.n41 plus.n24 3.65202
R63 plus.n31 plus.n26 3.65202
R64 plus.n9 plus.n4 0.189894
R65 plus.n10 plus.n9 0.189894
R66 plus.n10 plus.n2 0.189894
R67 plus.n16 plus.n2 0.189894
R68 plus.n17 plus.n16 0.189894
R69 plus.n17 plus.n0 0.189894
R70 plus.n22 plus.n0 0.189894
R71 plus.n45 plus.n23 0.189894
R72 plus.n40 plus.n23 0.189894
R73 plus.n40 plus.n39 0.189894
R74 plus.n39 plus.n25 0.189894
R75 plus.n33 plus.n25 0.189894
R76 plus.n33 plus.n32 0.189894
R77 plus.n32 plus.n27 0.189894
R78 drain_left.n9 drain_left.n7 80.3335
R79 drain_left.n5 drain_left.n3 80.3334
R80 drain_left.n2 drain_left.n0 80.3334
R81 drain_left.n13 drain_left.n12 79.7731
R82 drain_left.n11 drain_left.n10 79.7731
R83 drain_left.n9 drain_left.n8 79.7731
R84 drain_left.n5 drain_left.n4 79.773
R85 drain_left.n2 drain_left.n1 79.773
R86 drain_left drain_left.n6 24.1911
R87 drain_left.n3 drain_left.t13 10.0005
R88 drain_left.n3 drain_left.t12 10.0005
R89 drain_left.n4 drain_left.t6 10.0005
R90 drain_left.n4 drain_left.t9 10.0005
R91 drain_left.n1 drain_left.t14 10.0005
R92 drain_left.n1 drain_left.t11 10.0005
R93 drain_left.n0 drain_left.t15 10.0005
R94 drain_left.n0 drain_left.t1 10.0005
R95 drain_left.n12 drain_left.t0 10.0005
R96 drain_left.n12 drain_left.t5 10.0005
R97 drain_left.n10 drain_left.t3 10.0005
R98 drain_left.n10 drain_left.t8 10.0005
R99 drain_left.n8 drain_left.t4 10.0005
R100 drain_left.n8 drain_left.t7 10.0005
R101 drain_left.n7 drain_left.t10 10.0005
R102 drain_left.n7 drain_left.t2 10.0005
R103 drain_left drain_left.n13 6.21356
R104 drain_left.n11 drain_left.n9 0.560845
R105 drain_left.n13 drain_left.n11 0.560845
R106 drain_left.n6 drain_left.n5 0.225326
R107 drain_left.n6 drain_left.n2 0.225326
R108 source.n0 source.t24 73.0943
R109 source.n7 source.t23 73.0943
R110 source.n8 source.t15 73.0943
R111 source.n15 source.t10 73.0943
R112 source.n31 source.t3 73.0942
R113 source.n24 source.t1 73.0942
R114 source.n23 source.t29 73.0942
R115 source.n16 source.t25 73.0942
R116 source.n2 source.n1 63.0943
R117 source.n4 source.n3 63.0943
R118 source.n6 source.n5 63.0943
R119 source.n10 source.n9 63.0943
R120 source.n12 source.n11 63.0943
R121 source.n14 source.n13 63.0943
R122 source.n30 source.n29 63.0942
R123 source.n28 source.n27 63.0942
R124 source.n26 source.n25 63.0942
R125 source.n22 source.n21 63.0942
R126 source.n20 source.n19 63.0942
R127 source.n18 source.n17 63.0942
R128 source.n16 source.n15 15.0299
R129 source.n29 source.t0 10.0005
R130 source.n29 source.t9 10.0005
R131 source.n27 source.t12 10.0005
R132 source.n27 source.t13 10.0005
R133 source.n25 source.t7 10.0005
R134 source.n25 source.t6 10.0005
R135 source.n21 source.t26 10.0005
R136 source.n21 source.t30 10.0005
R137 source.n19 source.t28 10.0005
R138 source.n19 source.t27 10.0005
R139 source.n17 source.t19 10.0005
R140 source.n17 source.t31 10.0005
R141 source.n1 source.t18 10.0005
R142 source.n1 source.t21 10.0005
R143 source.n3 source.t22 10.0005
R144 source.n3 source.t16 10.0005
R145 source.n5 source.t17 10.0005
R146 source.n5 source.t20 10.0005
R147 source.n9 source.t4 10.0005
R148 source.n9 source.t11 10.0005
R149 source.n11 source.t2 10.0005
R150 source.n11 source.t14 10.0005
R151 source.n13 source.t8 10.0005
R152 source.n13 source.t5 10.0005
R153 source.n32 source.n0 9.48679
R154 source.n32 source.n31 5.5436
R155 source.n15 source.n14 0.560845
R156 source.n14 source.n12 0.560845
R157 source.n12 source.n10 0.560845
R158 source.n10 source.n8 0.560845
R159 source.n7 source.n6 0.560845
R160 source.n6 source.n4 0.560845
R161 source.n4 source.n2 0.560845
R162 source.n2 source.n0 0.560845
R163 source.n18 source.n16 0.560845
R164 source.n20 source.n18 0.560845
R165 source.n22 source.n20 0.560845
R166 source.n23 source.n22 0.560845
R167 source.n26 source.n24 0.560845
R168 source.n28 source.n26 0.560845
R169 source.n30 source.n28 0.560845
R170 source.n31 source.n30 0.560845
R171 source.n8 source.n7 0.470328
R172 source.n24 source.n23 0.470328
R173 source source.n32 0.188
R174 minus.n21 minus.t12 731.034
R175 minus.n5 minus.t7 731.034
R176 minus.n44 minus.t0 731.034
R177 minus.n28 minus.t5 731.034
R178 minus.n20 minus.t11 690.867
R179 minus.n1 minus.t13 690.867
R180 minus.n14 minus.t8 690.867
R181 minus.n12 minus.t9 690.867
R182 minus.n3 minus.t10 690.867
R183 minus.n6 minus.t6 690.867
R184 minus.n43 minus.t2 690.867
R185 minus.n24 minus.t3 690.867
R186 minus.n37 minus.t4 690.867
R187 minus.n35 minus.t14 690.867
R188 minus.n26 minus.t15 690.867
R189 minus.n29 minus.t1 690.867
R190 minus.n5 minus.n4 161.489
R191 minus.n28 minus.n27 161.489
R192 minus.n22 minus.n21 161.3
R193 minus.n19 minus.n0 161.3
R194 minus.n18 minus.n17 161.3
R195 minus.n16 minus.n15 161.3
R196 minus.n13 minus.n2 161.3
R197 minus.n11 minus.n10 161.3
R198 minus.n9 minus.n8 161.3
R199 minus.n7 minus.n4 161.3
R200 minus.n45 minus.n44 161.3
R201 minus.n42 minus.n23 161.3
R202 minus.n41 minus.n40 161.3
R203 minus.n39 minus.n38 161.3
R204 minus.n36 minus.n25 161.3
R205 minus.n34 minus.n33 161.3
R206 minus.n32 minus.n31 161.3
R207 minus.n30 minus.n27 161.3
R208 minus.n19 minus.n18 73.0308
R209 minus.n8 minus.n7 73.0308
R210 minus.n31 minus.n30 73.0308
R211 minus.n42 minus.n41 73.0308
R212 minus.n15 minus.n1 69.3793
R213 minus.n11 minus.n3 69.3793
R214 minus.n34 minus.n26 69.3793
R215 minus.n38 minus.n24 69.3793
R216 minus.n21 minus.n20 54.7732
R217 minus.n6 minus.n5 54.7732
R218 minus.n29 minus.n28 54.7732
R219 minus.n44 minus.n43 54.7732
R220 minus.n14 minus.n13 47.4702
R221 minus.n13 minus.n12 47.4702
R222 minus.n36 minus.n35 47.4702
R223 minus.n37 minus.n36 47.4702
R224 minus.n46 minus.n22 29.4513
R225 minus.n15 minus.n14 25.5611
R226 minus.n12 minus.n11 25.5611
R227 minus.n35 minus.n34 25.5611
R228 minus.n38 minus.n37 25.5611
R229 minus.n20 minus.n19 18.2581
R230 minus.n7 minus.n6 18.2581
R231 minus.n30 minus.n29 18.2581
R232 minus.n43 minus.n42 18.2581
R233 minus.n46 minus.n45 6.50429
R234 minus.n18 minus.n1 3.65202
R235 minus.n8 minus.n3 3.65202
R236 minus.n31 minus.n26 3.65202
R237 minus.n41 minus.n24 3.65202
R238 minus.n22 minus.n0 0.189894
R239 minus.n17 minus.n0 0.189894
R240 minus.n17 minus.n16 0.189894
R241 minus.n16 minus.n2 0.189894
R242 minus.n10 minus.n2 0.189894
R243 minus.n10 minus.n9 0.189894
R244 minus.n9 minus.n4 0.189894
R245 minus.n32 minus.n27 0.189894
R246 minus.n33 minus.n32 0.189894
R247 minus.n33 minus.n25 0.189894
R248 minus.n39 minus.n25 0.189894
R249 minus.n40 minus.n39 0.189894
R250 minus.n40 minus.n23 0.189894
R251 minus.n45 minus.n23 0.189894
R252 minus minus.n46 0.188
R253 drain_right.n9 drain_right.n7 80.3335
R254 drain_right.n5 drain_right.n3 80.3334
R255 drain_right.n2 drain_right.n0 80.3334
R256 drain_right.n9 drain_right.n8 79.7731
R257 drain_right.n11 drain_right.n10 79.7731
R258 drain_right.n13 drain_right.n12 79.7731
R259 drain_right.n5 drain_right.n4 79.773
R260 drain_right.n2 drain_right.n1 79.773
R261 drain_right drain_right.n6 23.6379
R262 drain_right.n3 drain_right.t13 10.0005
R263 drain_right.n3 drain_right.t15 10.0005
R264 drain_right.n4 drain_right.t11 10.0005
R265 drain_right.n4 drain_right.t12 10.0005
R266 drain_right.n1 drain_right.t0 10.0005
R267 drain_right.n1 drain_right.t1 10.0005
R268 drain_right.n0 drain_right.t10 10.0005
R269 drain_right.n0 drain_right.t14 10.0005
R270 drain_right.n7 drain_right.t9 10.0005
R271 drain_right.n7 drain_right.t8 10.0005
R272 drain_right.n8 drain_right.t6 10.0005
R273 drain_right.n8 drain_right.t5 10.0005
R274 drain_right.n10 drain_right.t2 10.0005
R275 drain_right.n10 drain_right.t7 10.0005
R276 drain_right.n12 drain_right.t3 10.0005
R277 drain_right.n12 drain_right.t4 10.0005
R278 drain_right drain_right.n13 6.21356
R279 drain_right.n13 drain_right.n11 0.560845
R280 drain_right.n11 drain_right.n9 0.560845
R281 drain_right.n6 drain_right.n5 0.225326
R282 drain_right.n6 drain_right.n2 0.225326
C0 drain_left minus 0.176066f
C1 drain_right source 9.94735f
C2 plus source 1.31511f
C3 minus source 1.30111f
C4 drain_right plus 0.342914f
C5 drain_left source 9.947001f
C6 drain_right minus 1.27334f
C7 drain_right drain_left 0.96779f
C8 plus minus 3.83258f
C9 plus drain_left 1.45691f
C10 drain_right a_n1886_n1488# 4.098259f
C11 drain_left a_n1886_n1488# 4.35584f
C12 source a_n1886_n1488# 3.769038f
C13 minus a_n1886_n1488# 6.244088f
C14 plus a_n1886_n1488# 7.015201f
C15 drain_right.t10 a_n1886_n1488# 0.088466f
C16 drain_right.t14 a_n1886_n1488# 0.088466f
C17 drain_right.n0 a_n1886_n1488# 0.483308f
C18 drain_right.t0 a_n1886_n1488# 0.088466f
C19 drain_right.t1 a_n1886_n1488# 0.088466f
C20 drain_right.n1 a_n1886_n1488# 0.481243f
C21 drain_right.n2 a_n1886_n1488# 0.555946f
C22 drain_right.t13 a_n1886_n1488# 0.088466f
C23 drain_right.t15 a_n1886_n1488# 0.088466f
C24 drain_right.n3 a_n1886_n1488# 0.483308f
C25 drain_right.t11 a_n1886_n1488# 0.088466f
C26 drain_right.t12 a_n1886_n1488# 0.088466f
C27 drain_right.n4 a_n1886_n1488# 0.481243f
C28 drain_right.n5 a_n1886_n1488# 0.555946f
C29 drain_right.n6 a_n1886_n1488# 0.707533f
C30 drain_right.t9 a_n1886_n1488# 0.088466f
C31 drain_right.t8 a_n1886_n1488# 0.088466f
C32 drain_right.n7 a_n1886_n1488# 0.48331f
C33 drain_right.t6 a_n1886_n1488# 0.088466f
C34 drain_right.t5 a_n1886_n1488# 0.088466f
C35 drain_right.n8 a_n1886_n1488# 0.481245f
C36 drain_right.n9 a_n1886_n1488# 0.580029f
C37 drain_right.t2 a_n1886_n1488# 0.088466f
C38 drain_right.t7 a_n1886_n1488# 0.088466f
C39 drain_right.n10 a_n1886_n1488# 0.481245f
C40 drain_right.n11 a_n1886_n1488# 0.286087f
C41 drain_right.t3 a_n1886_n1488# 0.088466f
C42 drain_right.t4 a_n1886_n1488# 0.088466f
C43 drain_right.n12 a_n1886_n1488# 0.481245f
C44 drain_right.n13 a_n1886_n1488# 0.491765f
C45 minus.n0 a_n1886_n1488# 0.031076f
C46 minus.t12 a_n1886_n1488# 0.041973f
C47 minus.t11 a_n1886_n1488# 0.040497f
C48 minus.t13 a_n1886_n1488# 0.040497f
C49 minus.n1 a_n1886_n1488# 0.028304f
C50 minus.n2 a_n1886_n1488# 0.031076f
C51 minus.t8 a_n1886_n1488# 0.040497f
C52 minus.t9 a_n1886_n1488# 0.040497f
C53 minus.t10 a_n1886_n1488# 0.040497f
C54 minus.n3 a_n1886_n1488# 0.028304f
C55 minus.n4 a_n1886_n1488# 0.065943f
C56 minus.t6 a_n1886_n1488# 0.040497f
C57 minus.t7 a_n1886_n1488# 0.041973f
C58 minus.n5 a_n1886_n1488# 0.038615f
C59 minus.n6 a_n1886_n1488# 0.028304f
C60 minus.n7 a_n1886_n1488# 0.012704f
C61 minus.n8 a_n1886_n1488# 0.010788f
C62 minus.n9 a_n1886_n1488# 0.031076f
C63 minus.n10 a_n1886_n1488# 0.031076f
C64 minus.n11 a_n1886_n1488# 0.013183f
C65 minus.n12 a_n1886_n1488# 0.028304f
C66 minus.n13 a_n1886_n1488# 0.013183f
C67 minus.n14 a_n1886_n1488# 0.028304f
C68 minus.n15 a_n1886_n1488# 0.013183f
C69 minus.n16 a_n1886_n1488# 0.031076f
C70 minus.n17 a_n1886_n1488# 0.031076f
C71 minus.n18 a_n1886_n1488# 0.010788f
C72 minus.n19 a_n1886_n1488# 0.012704f
C73 minus.n20 a_n1886_n1488# 0.028304f
C74 minus.n21 a_n1886_n1488# 0.038574f
C75 minus.n22 a_n1886_n1488# 0.783345f
C76 minus.n23 a_n1886_n1488# 0.031076f
C77 minus.t2 a_n1886_n1488# 0.040497f
C78 minus.t3 a_n1886_n1488# 0.040497f
C79 minus.n24 a_n1886_n1488# 0.028304f
C80 minus.n25 a_n1886_n1488# 0.031076f
C81 minus.t4 a_n1886_n1488# 0.040497f
C82 minus.t14 a_n1886_n1488# 0.040497f
C83 minus.t15 a_n1886_n1488# 0.040497f
C84 minus.n26 a_n1886_n1488# 0.028304f
C85 minus.n27 a_n1886_n1488# 0.065943f
C86 minus.t1 a_n1886_n1488# 0.040497f
C87 minus.t5 a_n1886_n1488# 0.041973f
C88 minus.n28 a_n1886_n1488# 0.038615f
C89 minus.n29 a_n1886_n1488# 0.028304f
C90 minus.n30 a_n1886_n1488# 0.012704f
C91 minus.n31 a_n1886_n1488# 0.010788f
C92 minus.n32 a_n1886_n1488# 0.031076f
C93 minus.n33 a_n1886_n1488# 0.031076f
C94 minus.n34 a_n1886_n1488# 0.013183f
C95 minus.n35 a_n1886_n1488# 0.028304f
C96 minus.n36 a_n1886_n1488# 0.013183f
C97 minus.n37 a_n1886_n1488# 0.028304f
C98 minus.n38 a_n1886_n1488# 0.013183f
C99 minus.n39 a_n1886_n1488# 0.031076f
C100 minus.n40 a_n1886_n1488# 0.031076f
C101 minus.n41 a_n1886_n1488# 0.010788f
C102 minus.n42 a_n1886_n1488# 0.012704f
C103 minus.n43 a_n1886_n1488# 0.028304f
C104 minus.t0 a_n1886_n1488# 0.041973f
C105 minus.n44 a_n1886_n1488# 0.038574f
C106 minus.n45 a_n1886_n1488# 0.203482f
C107 minus.n46 a_n1886_n1488# 0.967018f
C108 source.t24 a_n1886_n1488# 0.505824f
C109 source.n0 a_n1886_n1488# 0.667751f
C110 source.t18 a_n1886_n1488# 0.085882f
C111 source.t21 a_n1886_n1488# 0.085882f
C112 source.n1 a_n1886_n1488# 0.417795f
C113 source.n2 a_n1886_n1488# 0.294622f
C114 source.t22 a_n1886_n1488# 0.085882f
C115 source.t16 a_n1886_n1488# 0.085882f
C116 source.n3 a_n1886_n1488# 0.417795f
C117 source.n4 a_n1886_n1488# 0.294622f
C118 source.t17 a_n1886_n1488# 0.085882f
C119 source.t20 a_n1886_n1488# 0.085882f
C120 source.n5 a_n1886_n1488# 0.417795f
C121 source.n6 a_n1886_n1488# 0.294622f
C122 source.t23 a_n1886_n1488# 0.505824f
C123 source.n7 a_n1886_n1488# 0.354206f
C124 source.t15 a_n1886_n1488# 0.505824f
C125 source.n8 a_n1886_n1488# 0.354206f
C126 source.t4 a_n1886_n1488# 0.085882f
C127 source.t11 a_n1886_n1488# 0.085882f
C128 source.n9 a_n1886_n1488# 0.417795f
C129 source.n10 a_n1886_n1488# 0.294622f
C130 source.t2 a_n1886_n1488# 0.085882f
C131 source.t14 a_n1886_n1488# 0.085882f
C132 source.n11 a_n1886_n1488# 0.417795f
C133 source.n12 a_n1886_n1488# 0.294622f
C134 source.t8 a_n1886_n1488# 0.085882f
C135 source.t5 a_n1886_n1488# 0.085882f
C136 source.n13 a_n1886_n1488# 0.417795f
C137 source.n14 a_n1886_n1488# 0.294622f
C138 source.t10 a_n1886_n1488# 0.505824f
C139 source.n15 a_n1886_n1488# 0.917292f
C140 source.t25 a_n1886_n1488# 0.505821f
C141 source.n16 a_n1886_n1488# 0.917295f
C142 source.t19 a_n1886_n1488# 0.085882f
C143 source.t31 a_n1886_n1488# 0.085882f
C144 source.n17 a_n1886_n1488# 0.417793f
C145 source.n18 a_n1886_n1488# 0.294624f
C146 source.t28 a_n1886_n1488# 0.085882f
C147 source.t27 a_n1886_n1488# 0.085882f
C148 source.n19 a_n1886_n1488# 0.417793f
C149 source.n20 a_n1886_n1488# 0.294624f
C150 source.t26 a_n1886_n1488# 0.085882f
C151 source.t30 a_n1886_n1488# 0.085882f
C152 source.n21 a_n1886_n1488# 0.417793f
C153 source.n22 a_n1886_n1488# 0.294624f
C154 source.t29 a_n1886_n1488# 0.505821f
C155 source.n23 a_n1886_n1488# 0.354209f
C156 source.t1 a_n1886_n1488# 0.505821f
C157 source.n24 a_n1886_n1488# 0.354209f
C158 source.t7 a_n1886_n1488# 0.085882f
C159 source.t6 a_n1886_n1488# 0.085882f
C160 source.n25 a_n1886_n1488# 0.417793f
C161 source.n26 a_n1886_n1488# 0.294624f
C162 source.t12 a_n1886_n1488# 0.085882f
C163 source.t13 a_n1886_n1488# 0.085882f
C164 source.n27 a_n1886_n1488# 0.417793f
C165 source.n28 a_n1886_n1488# 0.294624f
C166 source.t0 a_n1886_n1488# 0.085882f
C167 source.t9 a_n1886_n1488# 0.085882f
C168 source.n29 a_n1886_n1488# 0.417793f
C169 source.n30 a_n1886_n1488# 0.294624f
C170 source.t3 a_n1886_n1488# 0.505821f
C171 source.n31 a_n1886_n1488# 0.490238f
C172 source.n32 a_n1886_n1488# 0.693604f
C173 drain_left.t15 a_n1886_n1488# 0.087614f
C174 drain_left.t1 a_n1886_n1488# 0.087614f
C175 drain_left.n0 a_n1886_n1488# 0.478649f
C176 drain_left.t14 a_n1886_n1488# 0.087614f
C177 drain_left.t11 a_n1886_n1488# 0.087614f
C178 drain_left.n1 a_n1886_n1488# 0.476604f
C179 drain_left.n2 a_n1886_n1488# 0.550588f
C180 drain_left.t13 a_n1886_n1488# 0.087614f
C181 drain_left.t12 a_n1886_n1488# 0.087614f
C182 drain_left.n3 a_n1886_n1488# 0.478649f
C183 drain_left.t6 a_n1886_n1488# 0.087614f
C184 drain_left.t9 a_n1886_n1488# 0.087614f
C185 drain_left.n4 a_n1886_n1488# 0.476604f
C186 drain_left.n5 a_n1886_n1488# 0.550588f
C187 drain_left.n6 a_n1886_n1488# 0.749015f
C188 drain_left.t10 a_n1886_n1488# 0.087614f
C189 drain_left.t2 a_n1886_n1488# 0.087614f
C190 drain_left.n7 a_n1886_n1488# 0.478651f
C191 drain_left.t4 a_n1886_n1488# 0.087614f
C192 drain_left.t7 a_n1886_n1488# 0.087614f
C193 drain_left.n8 a_n1886_n1488# 0.476607f
C194 drain_left.n9 a_n1886_n1488# 0.574439f
C195 drain_left.t3 a_n1886_n1488# 0.087614f
C196 drain_left.t8 a_n1886_n1488# 0.087614f
C197 drain_left.n10 a_n1886_n1488# 0.476607f
C198 drain_left.n11 a_n1886_n1488# 0.28333f
C199 drain_left.t0 a_n1886_n1488# 0.087614f
C200 drain_left.t5 a_n1886_n1488# 0.087614f
C201 drain_left.n12 a_n1886_n1488# 0.476607f
C202 drain_left.n13 a_n1886_n1488# 0.487025f
C203 plus.n0 a_n1886_n1488# 0.031599f
C204 plus.t10 a_n1886_n1488# 0.041178f
C205 plus.t13 a_n1886_n1488# 0.041178f
C206 plus.n1 a_n1886_n1488# 0.02878f
C207 plus.n2 a_n1886_n1488# 0.031599f
C208 plus.t15 a_n1886_n1488# 0.041178f
C209 plus.t9 a_n1886_n1488# 0.041178f
C210 plus.t11 a_n1886_n1488# 0.041178f
C211 plus.n3 a_n1886_n1488# 0.02878f
C212 plus.n4 a_n1886_n1488# 0.067052f
C213 plus.t14 a_n1886_n1488# 0.041178f
C214 plus.t8 a_n1886_n1488# 0.042679f
C215 plus.n5 a_n1886_n1488# 0.039264f
C216 plus.n6 a_n1886_n1488# 0.02878f
C217 plus.n7 a_n1886_n1488# 0.012918f
C218 plus.n8 a_n1886_n1488# 0.010969f
C219 plus.n9 a_n1886_n1488# 0.031599f
C220 plus.n10 a_n1886_n1488# 0.031599f
C221 plus.n11 a_n1886_n1488# 0.013405f
C222 plus.n12 a_n1886_n1488# 0.02878f
C223 plus.n13 a_n1886_n1488# 0.013405f
C224 plus.n14 a_n1886_n1488# 0.02878f
C225 plus.n15 a_n1886_n1488# 0.013405f
C226 plus.n16 a_n1886_n1488# 0.031599f
C227 plus.n17 a_n1886_n1488# 0.031599f
C228 plus.n18 a_n1886_n1488# 0.010969f
C229 plus.n19 a_n1886_n1488# 0.012918f
C230 plus.n20 a_n1886_n1488# 0.02878f
C231 plus.t7 a_n1886_n1488# 0.042679f
C232 plus.n21 a_n1886_n1488# 0.039223f
C233 plus.n22 a_n1886_n1488# 0.236375f
C234 plus.n23 a_n1886_n1488# 0.031599f
C235 plus.t6 a_n1886_n1488# 0.042679f
C236 plus.t12 a_n1886_n1488# 0.041178f
C237 plus.t0 a_n1886_n1488# 0.041178f
C238 plus.n24 a_n1886_n1488# 0.02878f
C239 plus.n25 a_n1886_n1488# 0.031599f
C240 plus.t3 a_n1886_n1488# 0.041178f
C241 plus.t4 a_n1886_n1488# 0.041178f
C242 plus.t5 a_n1886_n1488# 0.041178f
C243 plus.n26 a_n1886_n1488# 0.02878f
C244 plus.n27 a_n1886_n1488# 0.067052f
C245 plus.t1 a_n1886_n1488# 0.041178f
C246 plus.t2 a_n1886_n1488# 0.042679f
C247 plus.n28 a_n1886_n1488# 0.039264f
C248 plus.n29 a_n1886_n1488# 0.02878f
C249 plus.n30 a_n1886_n1488# 0.012918f
C250 plus.n31 a_n1886_n1488# 0.010969f
C251 plus.n32 a_n1886_n1488# 0.031599f
C252 plus.n33 a_n1886_n1488# 0.031599f
C253 plus.n34 a_n1886_n1488# 0.013405f
C254 plus.n35 a_n1886_n1488# 0.02878f
C255 plus.n36 a_n1886_n1488# 0.013405f
C256 plus.n37 a_n1886_n1488# 0.02878f
C257 plus.n38 a_n1886_n1488# 0.013405f
C258 plus.n39 a_n1886_n1488# 0.031599f
C259 plus.n40 a_n1886_n1488# 0.031599f
C260 plus.n41 a_n1886_n1488# 0.010969f
C261 plus.n42 a_n1886_n1488# 0.012918f
C262 plus.n43 a_n1886_n1488# 0.02878f
C263 plus.n44 a_n1886_n1488# 0.039223f
C264 plus.n45 a_n1886_n1488# 0.749064f
.ends

