* NGSPICE file created from diffpair123.ext - technology: sky130A

.subckt diffpair123 minus drain_right drain_left source plus
X0 drain_right.t7 minus.t0 source.t8 a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X1 source.t6 plus.t0 drain_left.t7 a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X2 source.t11 minus.t1 drain_right.t6 a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X3 source.t5 plus.t1 drain_left.t6 a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X4 source.t2 plus.t2 drain_left.t5 a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X5 a_n1546_n1288# a_n1546_n1288# a_n1546_n1288# a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.5
X6 drain_right.t5 minus.t2 source.t9 a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X7 drain_left.t4 plus.t3 source.t4 a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X8 drain_right.t4 minus.t3 source.t15 a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X9 drain_left.t3 plus.t4 source.t3 a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X10 source.t13 minus.t4 drain_right.t3 a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X11 source.t10 minus.t5 drain_right.t2 a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X12 a_n1546_n1288# a_n1546_n1288# a_n1546_n1288# a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X13 drain_left.t2 plus.t5 source.t7 a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X14 a_n1546_n1288# a_n1546_n1288# a_n1546_n1288# a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X15 source.t12 minus.t6 drain_right.t1 a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.5
X16 a_n1546_n1288# a_n1546_n1288# a_n1546_n1288# a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.5
X17 drain_right.t0 minus.t7 source.t14 a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
X18 source.t0 plus.t6 drain_left.t1 a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.5
X19 drain_left.t0 plus.t7 source.t1 a_n1546_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.5
R0 minus.n2 minus.t3 195.948
R1 minus.n10 minus.t6 195.948
R2 minus.n1 minus.t1 174.966
R3 minus.n5 minus.t2 174.966
R4 minus.n6 minus.t5 174.966
R5 minus.n9 minus.t0 174.966
R6 minus.n13 minus.t4 174.966
R7 minus.n14 minus.t7 174.966
R8 minus.n7 minus.n6 161.3
R9 minus.n5 minus.n0 161.3
R10 minus.n4 minus.n3 161.3
R11 minus.n15 minus.n14 161.3
R12 minus.n13 minus.n8 161.3
R13 minus.n12 minus.n11 161.3
R14 minus.n3 minus.n2 70.4033
R15 minus.n11 minus.n10 70.4033
R16 minus.n6 minus.n5 48.2005
R17 minus.n14 minus.n13 48.2005
R18 minus.n16 minus.n7 27.4967
R19 minus.n5 minus.n4 24.1005
R20 minus.n4 minus.n1 24.1005
R21 minus.n12 minus.n9 24.1005
R22 minus.n13 minus.n12 24.1005
R23 minus.n2 minus.n1 20.9576
R24 minus.n10 minus.n9 20.9576
R25 minus.n16 minus.n15 6.5952
R26 minus.n7 minus.n0 0.189894
R27 minus.n3 minus.n0 0.189894
R28 minus.n11 minus.n8 0.189894
R29 minus.n15 minus.n8 0.189894
R30 minus minus.n16 0.188
R31 source.n66 source.n64 289.615
R32 source.n56 source.n54 289.615
R33 source.n48 source.n46 289.615
R34 source.n38 source.n36 289.615
R35 source.n2 source.n0 289.615
R36 source.n12 source.n10 289.615
R37 source.n20 source.n18 289.615
R38 source.n30 source.n28 289.615
R39 source.n67 source.n66 185
R40 source.n57 source.n56 185
R41 source.n49 source.n48 185
R42 source.n39 source.n38 185
R43 source.n3 source.n2 185
R44 source.n13 source.n12 185
R45 source.n21 source.n20 185
R46 source.n31 source.n30 185
R47 source.t14 source.n65 167.117
R48 source.t12 source.n55 167.117
R49 source.t1 source.n47 167.117
R50 source.t2 source.n37 167.117
R51 source.t4 source.n1 167.117
R52 source.t5 source.n11 167.117
R53 source.t15 source.n19 167.117
R54 source.t10 source.n29 167.117
R55 source.n9 source.n8 84.1169
R56 source.n27 source.n26 84.1169
R57 source.n63 source.n62 84.1168
R58 source.n45 source.n44 84.1168
R59 source.n66 source.t14 52.3082
R60 source.n56 source.t12 52.3082
R61 source.n48 source.t1 52.3082
R62 source.n38 source.t2 52.3082
R63 source.n2 source.t4 52.3082
R64 source.n12 source.t5 52.3082
R65 source.n20 source.t15 52.3082
R66 source.n30 source.t10 52.3082
R67 source.n71 source.n70 31.4096
R68 source.n61 source.n60 31.4096
R69 source.n53 source.n52 31.4096
R70 source.n43 source.n42 31.4096
R71 source.n7 source.n6 31.4096
R72 source.n17 source.n16 31.4096
R73 source.n25 source.n24 31.4096
R74 source.n35 source.n34 31.4096
R75 source.n43 source.n35 14.4275
R76 source.n62 source.t8 9.9005
R77 source.n62 source.t13 9.9005
R78 source.n44 source.t7 9.9005
R79 source.n44 source.t6 9.9005
R80 source.n8 source.t3 9.9005
R81 source.n8 source.t0 9.9005
R82 source.n26 source.t9 9.9005
R83 source.n26 source.t11 9.9005
R84 source.n67 source.n65 9.71174
R85 source.n57 source.n55 9.71174
R86 source.n49 source.n47 9.71174
R87 source.n39 source.n37 9.71174
R88 source.n3 source.n1 9.71174
R89 source.n13 source.n11 9.71174
R90 source.n21 source.n19 9.71174
R91 source.n31 source.n29 9.71174
R92 source.n70 source.n69 9.45567
R93 source.n60 source.n59 9.45567
R94 source.n52 source.n51 9.45567
R95 source.n42 source.n41 9.45567
R96 source.n6 source.n5 9.45567
R97 source.n16 source.n15 9.45567
R98 source.n24 source.n23 9.45567
R99 source.n34 source.n33 9.45567
R100 source.n69 source.n68 9.3005
R101 source.n59 source.n58 9.3005
R102 source.n51 source.n50 9.3005
R103 source.n41 source.n40 9.3005
R104 source.n5 source.n4 9.3005
R105 source.n15 source.n14 9.3005
R106 source.n23 source.n22 9.3005
R107 source.n33 source.n32 9.3005
R108 source.n72 source.n7 8.8068
R109 source.n70 source.n64 8.14595
R110 source.n60 source.n54 8.14595
R111 source.n52 source.n46 8.14595
R112 source.n42 source.n36 8.14595
R113 source.n6 source.n0 8.14595
R114 source.n16 source.n10 8.14595
R115 source.n24 source.n18 8.14595
R116 source.n34 source.n28 8.14595
R117 source.n68 source.n67 7.3702
R118 source.n58 source.n57 7.3702
R119 source.n50 source.n49 7.3702
R120 source.n40 source.n39 7.3702
R121 source.n4 source.n3 7.3702
R122 source.n14 source.n13 7.3702
R123 source.n22 source.n21 7.3702
R124 source.n32 source.n31 7.3702
R125 source.n68 source.n64 5.81868
R126 source.n58 source.n54 5.81868
R127 source.n50 source.n46 5.81868
R128 source.n40 source.n36 5.81868
R129 source.n4 source.n0 5.81868
R130 source.n14 source.n10 5.81868
R131 source.n22 source.n18 5.81868
R132 source.n32 source.n28 5.81868
R133 source.n72 source.n71 5.62119
R134 source.n69 source.n65 3.44771
R135 source.n59 source.n55 3.44771
R136 source.n51 source.n47 3.44771
R137 source.n41 source.n37 3.44771
R138 source.n5 source.n1 3.44771
R139 source.n15 source.n11 3.44771
R140 source.n23 source.n19 3.44771
R141 source.n33 source.n29 3.44771
R142 source.n35 source.n27 0.716017
R143 source.n27 source.n25 0.716017
R144 source.n17 source.n9 0.716017
R145 source.n9 source.n7 0.716017
R146 source.n45 source.n43 0.716017
R147 source.n53 source.n45 0.716017
R148 source.n63 source.n61 0.716017
R149 source.n71 source.n63 0.716017
R150 source.n25 source.n17 0.470328
R151 source.n61 source.n53 0.470328
R152 source source.n72 0.188
R153 drain_right.n5 drain_right.n3 101.511
R154 drain_right.n2 drain_right.n1 101.099
R155 drain_right.n2 drain_right.n0 101.099
R156 drain_right.n5 drain_right.n4 100.796
R157 drain_right drain_right.n2 21.7424
R158 drain_right.n1 drain_right.t3 9.9005
R159 drain_right.n1 drain_right.t0 9.9005
R160 drain_right.n0 drain_right.t1 9.9005
R161 drain_right.n0 drain_right.t7 9.9005
R162 drain_right.n3 drain_right.t6 9.9005
R163 drain_right.n3 drain_right.t4 9.9005
R164 drain_right.n4 drain_right.t2 9.9005
R165 drain_right.n4 drain_right.t5 9.9005
R166 drain_right drain_right.n5 6.36873
R167 plus.n2 plus.t1 195.948
R168 plus.n10 plus.t7 195.948
R169 plus.n6 plus.t3 174.966
R170 plus.n5 plus.t6 174.966
R171 plus.n1 plus.t4 174.966
R172 plus.n14 plus.t2 174.966
R173 plus.n13 plus.t5 174.966
R174 plus.n9 plus.t0 174.966
R175 plus.n4 plus.n3 161.3
R176 plus.n5 plus.n0 161.3
R177 plus.n7 plus.n6 161.3
R178 plus.n12 plus.n11 161.3
R179 plus.n13 plus.n8 161.3
R180 plus.n15 plus.n14 161.3
R181 plus.n3 plus.n2 70.4033
R182 plus.n11 plus.n10 70.4033
R183 plus.n6 plus.n5 48.2005
R184 plus.n14 plus.n13 48.2005
R185 plus plus.n15 25.1657
R186 plus.n4 plus.n1 24.1005
R187 plus.n5 plus.n4 24.1005
R188 plus.n13 plus.n12 24.1005
R189 plus.n12 plus.n9 24.1005
R190 plus.n2 plus.n1 20.9576
R191 plus.n10 plus.n9 20.9576
R192 plus plus.n7 8.45126
R193 plus.n3 plus.n0 0.189894
R194 plus.n7 plus.n0 0.189894
R195 plus.n15 plus.n8 0.189894
R196 plus.n11 plus.n8 0.189894
R197 drain_left.n5 drain_left.n3 101.511
R198 drain_left.n2 drain_left.n1 101.099
R199 drain_left.n2 drain_left.n0 101.099
R200 drain_left.n5 drain_left.n4 100.796
R201 drain_left drain_left.n2 22.2956
R202 drain_left.n1 drain_left.t7 9.9005
R203 drain_left.n1 drain_left.t0 9.9005
R204 drain_left.n0 drain_left.t5 9.9005
R205 drain_left.n0 drain_left.t2 9.9005
R206 drain_left.n4 drain_left.t1 9.9005
R207 drain_left.n4 drain_left.t4 9.9005
R208 drain_left.n3 drain_left.t6 9.9005
R209 drain_left.n3 drain_left.t3 9.9005
R210 drain_left drain_left.n5 6.36873
C0 drain_left source 3.8364f
C1 source minus 1.25807f
C2 drain_left minus 0.176992f
C3 drain_right source 3.83689f
C4 drain_left drain_right 0.727126f
C5 drain_right minus 1.07242f
C6 plus source 1.27203f
C7 drain_left plus 1.22043f
C8 plus minus 3.22742f
C9 drain_right plus 0.308666f
C10 drain_right a_n1546_n1288# 3.15935f
C11 drain_left a_n1546_n1288# 3.35511f
C12 source a_n1546_n1288# 2.968916f
C13 minus a_n1546_n1288# 5.156103f
C14 plus a_n1546_n1288# 5.762223f
C15 drain_left.t5 a_n1546_n1288# 0.032043f
C16 drain_left.t2 a_n1546_n1288# 0.032043f
C17 drain_left.n0 a_n1546_n1288# 0.201999f
C18 drain_left.t7 a_n1546_n1288# 0.032043f
C19 drain_left.t0 a_n1546_n1288# 0.032043f
C20 drain_left.n1 a_n1546_n1288# 0.201999f
C21 drain_left.n2 a_n1546_n1288# 0.990118f
C22 drain_left.t6 a_n1546_n1288# 0.032043f
C23 drain_left.t3 a_n1546_n1288# 0.032043f
C24 drain_left.n3 a_n1546_n1288# 0.203118f
C25 drain_left.t1 a_n1546_n1288# 0.032043f
C26 drain_left.t4 a_n1546_n1288# 0.032043f
C27 drain_left.n4 a_n1546_n1288# 0.201308f
C28 drain_left.n5 a_n1546_n1288# 0.677883f
C29 plus.n0 a_n1546_n1288# 0.029761f
C30 plus.t3 a_n1546_n1288# 0.092161f
C31 plus.t6 a_n1546_n1288# 0.092161f
C32 plus.t4 a_n1546_n1288# 0.092161f
C33 plus.n1 a_n1546_n1288# 0.069414f
C34 plus.t1 a_n1546_n1288# 0.099274f
C35 plus.n2 a_n1546_n1288# 0.059503f
C36 plus.n3 a_n1546_n1288# 0.098043f
C37 plus.n4 a_n1546_n1288# 0.006753f
C38 plus.n5 a_n1546_n1288# 0.069414f
C39 plus.n6 a_n1546_n1288# 0.066386f
C40 plus.n7 a_n1546_n1288# 0.219762f
C41 plus.n8 a_n1546_n1288# 0.029761f
C42 plus.t2 a_n1546_n1288# 0.092161f
C43 plus.t5 a_n1546_n1288# 0.092161f
C44 plus.t0 a_n1546_n1288# 0.092161f
C45 plus.n9 a_n1546_n1288# 0.069414f
C46 plus.t7 a_n1546_n1288# 0.099274f
C47 plus.n10 a_n1546_n1288# 0.059503f
C48 plus.n11 a_n1546_n1288# 0.098043f
C49 plus.n12 a_n1546_n1288# 0.006753f
C50 plus.n13 a_n1546_n1288# 0.069414f
C51 plus.n14 a_n1546_n1288# 0.066386f
C52 plus.n15 a_n1546_n1288# 0.639707f
C53 drain_right.t1 a_n1546_n1288# 0.032727f
C54 drain_right.t7 a_n1546_n1288# 0.032727f
C55 drain_right.n0 a_n1546_n1288# 0.206305f
C56 drain_right.t3 a_n1546_n1288# 0.032727f
C57 drain_right.t0 a_n1546_n1288# 0.032727f
C58 drain_right.n1 a_n1546_n1288# 0.206305f
C59 drain_right.n2 a_n1546_n1288# 0.97053f
C60 drain_right.t6 a_n1546_n1288# 0.032727f
C61 drain_right.t4 a_n1546_n1288# 0.032727f
C62 drain_right.n3 a_n1546_n1288# 0.207448f
C63 drain_right.t2 a_n1546_n1288# 0.032727f
C64 drain_right.t5 a_n1546_n1288# 0.032727f
C65 drain_right.n4 a_n1546_n1288# 0.205599f
C66 drain_right.n5 a_n1546_n1288# 0.692333f
C67 source.n0 a_n1546_n1288# 0.029442f
C68 source.n1 a_n1546_n1288# 0.065144f
C69 source.t4 a_n1546_n1288# 0.048887f
C70 source.n2 a_n1546_n1288# 0.050984f
C71 source.n3 a_n1546_n1288# 0.016435f
C72 source.n4 a_n1546_n1288# 0.010839f
C73 source.n5 a_n1546_n1288# 0.143593f
C74 source.n6 a_n1546_n1288# 0.032275f
C75 source.n7 a_n1546_n1288# 0.324446f
C76 source.t3 a_n1546_n1288# 0.031881f
C77 source.t0 a_n1546_n1288# 0.031881f
C78 source.n8 a_n1546_n1288# 0.170433f
C79 source.n9 a_n1546_n1288# 0.249841f
C80 source.n10 a_n1546_n1288# 0.029442f
C81 source.n11 a_n1546_n1288# 0.065144f
C82 source.t5 a_n1546_n1288# 0.048887f
C83 source.n12 a_n1546_n1288# 0.050984f
C84 source.n13 a_n1546_n1288# 0.016435f
C85 source.n14 a_n1546_n1288# 0.010839f
C86 source.n15 a_n1546_n1288# 0.143593f
C87 source.n16 a_n1546_n1288# 0.032275f
C88 source.n17 a_n1546_n1288# 0.093651f
C89 source.n18 a_n1546_n1288# 0.029442f
C90 source.n19 a_n1546_n1288# 0.065144f
C91 source.t15 a_n1546_n1288# 0.048887f
C92 source.n20 a_n1546_n1288# 0.050984f
C93 source.n21 a_n1546_n1288# 0.016435f
C94 source.n22 a_n1546_n1288# 0.010839f
C95 source.n23 a_n1546_n1288# 0.143593f
C96 source.n24 a_n1546_n1288# 0.032275f
C97 source.n25 a_n1546_n1288# 0.093651f
C98 source.t9 a_n1546_n1288# 0.031881f
C99 source.t11 a_n1546_n1288# 0.031881f
C100 source.n26 a_n1546_n1288# 0.170433f
C101 source.n27 a_n1546_n1288# 0.249841f
C102 source.n28 a_n1546_n1288# 0.029442f
C103 source.n29 a_n1546_n1288# 0.065144f
C104 source.t10 a_n1546_n1288# 0.048887f
C105 source.n30 a_n1546_n1288# 0.050984f
C106 source.n31 a_n1546_n1288# 0.016435f
C107 source.n32 a_n1546_n1288# 0.010839f
C108 source.n33 a_n1546_n1288# 0.143593f
C109 source.n34 a_n1546_n1288# 0.032275f
C110 source.n35 a_n1546_n1288# 0.515036f
C111 source.n36 a_n1546_n1288# 0.029442f
C112 source.n37 a_n1546_n1288# 0.065144f
C113 source.t2 a_n1546_n1288# 0.048887f
C114 source.n38 a_n1546_n1288# 0.050984f
C115 source.n39 a_n1546_n1288# 0.016435f
C116 source.n40 a_n1546_n1288# 0.010839f
C117 source.n41 a_n1546_n1288# 0.143593f
C118 source.n42 a_n1546_n1288# 0.032275f
C119 source.n43 a_n1546_n1288# 0.515036f
C120 source.t7 a_n1546_n1288# 0.031881f
C121 source.t6 a_n1546_n1288# 0.031881f
C122 source.n44 a_n1546_n1288# 0.170432f
C123 source.n45 a_n1546_n1288# 0.249842f
C124 source.n46 a_n1546_n1288# 0.029442f
C125 source.n47 a_n1546_n1288# 0.065144f
C126 source.t1 a_n1546_n1288# 0.048887f
C127 source.n48 a_n1546_n1288# 0.050984f
C128 source.n49 a_n1546_n1288# 0.016435f
C129 source.n50 a_n1546_n1288# 0.010839f
C130 source.n51 a_n1546_n1288# 0.143593f
C131 source.n52 a_n1546_n1288# 0.032275f
C132 source.n53 a_n1546_n1288# 0.093651f
C133 source.n54 a_n1546_n1288# 0.029442f
C134 source.n55 a_n1546_n1288# 0.065144f
C135 source.t12 a_n1546_n1288# 0.048887f
C136 source.n56 a_n1546_n1288# 0.050984f
C137 source.n57 a_n1546_n1288# 0.016435f
C138 source.n58 a_n1546_n1288# 0.010839f
C139 source.n59 a_n1546_n1288# 0.143593f
C140 source.n60 a_n1546_n1288# 0.032275f
C141 source.n61 a_n1546_n1288# 0.093651f
C142 source.t8 a_n1546_n1288# 0.031881f
C143 source.t13 a_n1546_n1288# 0.031881f
C144 source.n62 a_n1546_n1288# 0.170432f
C145 source.n63 a_n1546_n1288# 0.249842f
C146 source.n64 a_n1546_n1288# 0.029442f
C147 source.n65 a_n1546_n1288# 0.065144f
C148 source.t14 a_n1546_n1288# 0.048887f
C149 source.n66 a_n1546_n1288# 0.050984f
C150 source.n67 a_n1546_n1288# 0.016435f
C151 source.n68 a_n1546_n1288# 0.010839f
C152 source.n69 a_n1546_n1288# 0.143593f
C153 source.n70 a_n1546_n1288# 0.032275f
C154 source.n71 a_n1546_n1288# 0.216426f
C155 source.n72 a_n1546_n1288# 0.503548f
C156 minus.n0 a_n1546_n1288# 0.029211f
C157 minus.t1 a_n1546_n1288# 0.090459f
C158 minus.n1 a_n1546_n1288# 0.068133f
C159 minus.t3 a_n1546_n1288# 0.097441f
C160 minus.n2 a_n1546_n1288# 0.058404f
C161 minus.n3 a_n1546_n1288# 0.096233f
C162 minus.n4 a_n1546_n1288# 0.006629f
C163 minus.t2 a_n1546_n1288# 0.090459f
C164 minus.n5 a_n1546_n1288# 0.068133f
C165 minus.t5 a_n1546_n1288# 0.090459f
C166 minus.n6 a_n1546_n1288# 0.065161f
C167 minus.n7 a_n1546_n1288# 0.655434f
C168 minus.n8 a_n1546_n1288# 0.029211f
C169 minus.t0 a_n1546_n1288# 0.090459f
C170 minus.n9 a_n1546_n1288# 0.068133f
C171 minus.t6 a_n1546_n1288# 0.097441f
C172 minus.n10 a_n1546_n1288# 0.058404f
C173 minus.n11 a_n1546_n1288# 0.096233f
C174 minus.n12 a_n1546_n1288# 0.006629f
C175 minus.t4 a_n1546_n1288# 0.090459f
C176 minus.n13 a_n1546_n1288# 0.068133f
C177 minus.t7 a_n1546_n1288# 0.090459f
C178 minus.n14 a_n1546_n1288# 0.065161f
C179 minus.n15 a_n1546_n1288# 0.197497f
C180 minus.n16 a_n1546_n1288# 0.806441f
.ends

