* NGSPICE file created from diffpair259.ext - technology: sky130A

.subckt diffpair259 minus drain_right drain_left source plus
X0 source.t47 minus.t0 drain_right.t0 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X1 source.t46 minus.t1 drain_right.t1 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X2 source.t22 plus.t0 drain_left.t23 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X3 source.t21 plus.t1 drain_left.t22 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X4 drain_right.t15 minus.t2 source.t45 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X5 drain_right.t22 minus.t3 source.t44 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X6 source.t43 minus.t4 drain_right.t20 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X7 drain_left.t21 plus.t2 source.t16 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X8 a_n2094_n2088# a_n2094_n2088# a_n2094_n2088# a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=0.2
X9 source.t42 minus.t5 drain_right.t19 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X10 a_n2094_n2088# a_n2094_n2088# a_n2094_n2088# a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X11 source.t15 plus.t3 drain_left.t20 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X12 drain_left.t19 plus.t4 source.t20 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X13 source.t17 plus.t5 drain_left.t18 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X14 drain_left.t17 plus.t6 source.t8 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X15 source.t11 plus.t7 drain_left.t16 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X16 source.t41 minus.t6 drain_right.t13 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X17 source.t0 plus.t8 drain_left.t15 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X18 source.t40 minus.t7 drain_right.t14 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X19 drain_left.t14 plus.t9 source.t1 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X20 source.t4 plus.t10 drain_left.t13 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X21 source.t39 minus.t8 drain_right.t23 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X22 drain_right.t5 minus.t9 source.t38 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X23 drain_left.t12 plus.t11 source.t7 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X24 drain_left.t11 plus.t12 source.t10 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X25 source.t5 plus.t13 drain_left.t10 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X26 a_n2094_n2088# a_n2094_n2088# a_n2094_n2088# a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X27 drain_left.t9 plus.t14 source.t13 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X28 drain_left.t8 plus.t15 source.t6 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X29 drain_left.t7 plus.t16 source.t18 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X30 drain_right.t8 minus.t10 source.t37 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X31 drain_right.t11 minus.t11 source.t36 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X32 drain_right.t17 minus.t12 source.t35 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X33 source.t23 plus.t17 drain_left.t6 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X34 source.t12 plus.t18 drain_left.t5 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X35 a_n2094_n2088# a_n2094_n2088# a_n2094_n2088# a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=0.2
X36 source.t2 plus.t19 drain_left.t4 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X37 drain_left.t3 plus.t20 source.t3 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X38 source.t34 minus.t13 drain_right.t6 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X39 source.t33 minus.t14 drain_right.t9 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X40 source.t32 minus.t15 drain_right.t2 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=0.2
X41 source.t31 minus.t16 drain_right.t16 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X42 source.t30 minus.t17 drain_right.t12 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X43 drain_right.t21 minus.t18 source.t29 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X44 drain_left.t2 plus.t21 source.t9 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=0.2
X45 drain_right.t18 minus.t19 source.t28 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X46 drain_right.t7 minus.t20 source.t27 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X47 drain_right.t10 minus.t21 source.t26 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X48 drain_left.t1 plus.t22 source.t14 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X49 source.t19 plus.t23 drain_left.t0 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X50 drain_right.t4 minus.t22 source.t25 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
X51 drain_right.t3 minus.t23 source.t24 a_n2094_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.2
R0 minus.n29 minus.t5 940.265
R1 minus.n6 minus.t11 940.265
R2 minus.n60 minus.t18 940.265
R3 minus.n37 minus.t15 940.265
R4 minus.n28 minus.t9 879.65
R5 minus.n26 minus.t8 879.65
R6 minus.n1 minus.t10 879.65
R7 minus.n21 minus.t17 879.65
R8 minus.n19 minus.t3 879.65
R9 minus.n3 minus.t6 879.65
R10 minus.n14 minus.t12 879.65
R11 minus.n12 minus.t16 879.65
R12 minus.n5 minus.t2 879.65
R13 minus.n7 minus.t7 879.65
R14 minus.n59 minus.t13 879.65
R15 minus.n57 minus.t19 879.65
R16 minus.n32 minus.t0 879.65
R17 minus.n52 minus.t22 879.65
R18 minus.n50 minus.t1 879.65
R19 minus.n34 minus.t23 879.65
R20 minus.n45 minus.t4 879.65
R21 minus.n43 minus.t20 879.65
R22 minus.n36 minus.t14 879.65
R23 minus.n38 minus.t21 879.65
R24 minus.n9 minus.n6 161.489
R25 minus.n40 minus.n37 161.489
R26 minus.n30 minus.n29 161.3
R27 minus.n27 minus.n0 161.3
R28 minus.n25 minus.n24 161.3
R29 minus.n23 minus.n22 161.3
R30 minus.n20 minus.n2 161.3
R31 minus.n18 minus.n17 161.3
R32 minus.n16 minus.n15 161.3
R33 minus.n13 minus.n4 161.3
R34 minus.n11 minus.n10 161.3
R35 minus.n9 minus.n8 161.3
R36 minus.n61 minus.n60 161.3
R37 minus.n58 minus.n31 161.3
R38 minus.n56 minus.n55 161.3
R39 minus.n54 minus.n53 161.3
R40 minus.n51 minus.n33 161.3
R41 minus.n49 minus.n48 161.3
R42 minus.n47 minus.n46 161.3
R43 minus.n44 minus.n35 161.3
R44 minus.n42 minus.n41 161.3
R45 minus.n40 minus.n39 161.3
R46 minus.n28 minus.n27 56.2338
R47 minus.n8 minus.n7 56.2338
R48 minus.n39 minus.n38 56.2338
R49 minus.n59 minus.n58 56.2338
R50 minus.n26 minus.n25 51.852
R51 minus.n11 minus.n5 51.852
R52 minus.n42 minus.n36 51.852
R53 minus.n57 minus.n56 51.852
R54 minus.n22 minus.n1 47.4702
R55 minus.n13 minus.n12 47.4702
R56 minus.n44 minus.n43 47.4702
R57 minus.n53 minus.n32 47.4702
R58 minus.n21 minus.n20 43.0884
R59 minus.n15 minus.n14 43.0884
R60 minus.n46 minus.n45 43.0884
R61 minus.n52 minus.n51 43.0884
R62 minus.n19 minus.n18 38.7066
R63 minus.n18 minus.n3 38.7066
R64 minus.n49 minus.n34 38.7066
R65 minus.n50 minus.n49 38.7066
R66 minus.n20 minus.n19 34.3247
R67 minus.n15 minus.n3 34.3247
R68 minus.n46 minus.n34 34.3247
R69 minus.n51 minus.n50 34.3247
R70 minus.n62 minus.n30 32.4967
R71 minus.n22 minus.n21 29.9429
R72 minus.n14 minus.n13 29.9429
R73 minus.n45 minus.n44 29.9429
R74 minus.n53 minus.n52 29.9429
R75 minus.n25 minus.n1 25.5611
R76 minus.n12 minus.n11 25.5611
R77 minus.n43 minus.n42 25.5611
R78 minus.n56 minus.n32 25.5611
R79 minus.n27 minus.n26 21.1793
R80 minus.n8 minus.n5 21.1793
R81 minus.n39 minus.n36 21.1793
R82 minus.n58 minus.n57 21.1793
R83 minus.n29 minus.n28 16.7975
R84 minus.n7 minus.n6 16.7975
R85 minus.n38 minus.n37 16.7975
R86 minus.n60 minus.n59 16.7975
R87 minus.n62 minus.n61 6.48914
R88 minus.n30 minus.n0 0.189894
R89 minus.n24 minus.n0 0.189894
R90 minus.n24 minus.n23 0.189894
R91 minus.n23 minus.n2 0.189894
R92 minus.n17 minus.n2 0.189894
R93 minus.n17 minus.n16 0.189894
R94 minus.n16 minus.n4 0.189894
R95 minus.n10 minus.n4 0.189894
R96 minus.n10 minus.n9 0.189894
R97 minus.n41 minus.n40 0.189894
R98 minus.n41 minus.n35 0.189894
R99 minus.n47 minus.n35 0.189894
R100 minus.n48 minus.n47 0.189894
R101 minus.n48 minus.n33 0.189894
R102 minus.n54 minus.n33 0.189894
R103 minus.n55 minus.n54 0.189894
R104 minus.n55 minus.n31 0.189894
R105 minus.n61 minus.n31 0.189894
R106 minus minus.n62 0.188
R107 drain_right.n7 drain_right.n5 67.6476
R108 drain_right.n2 drain_right.n0 67.6476
R109 drain_right.n13 drain_right.n11 67.6476
R110 drain_right.n13 drain_right.n12 67.1908
R111 drain_right.n15 drain_right.n14 67.1908
R112 drain_right.n17 drain_right.n16 67.1908
R113 drain_right.n19 drain_right.n18 67.1908
R114 drain_right.n21 drain_right.n20 67.1908
R115 drain_right.n7 drain_right.n6 67.1907
R116 drain_right.n9 drain_right.n8 67.1907
R117 drain_right.n4 drain_right.n3 67.1907
R118 drain_right.n2 drain_right.n1 67.1907
R119 drain_right drain_right.n10 26.6089
R120 drain_right drain_right.n21 6.11011
R121 drain_right.n5 drain_right.t6 3.3005
R122 drain_right.n5 drain_right.t21 3.3005
R123 drain_right.n6 drain_right.t0 3.3005
R124 drain_right.n6 drain_right.t18 3.3005
R125 drain_right.n8 drain_right.t1 3.3005
R126 drain_right.n8 drain_right.t4 3.3005
R127 drain_right.n3 drain_right.t20 3.3005
R128 drain_right.n3 drain_right.t3 3.3005
R129 drain_right.n1 drain_right.t9 3.3005
R130 drain_right.n1 drain_right.t7 3.3005
R131 drain_right.n0 drain_right.t2 3.3005
R132 drain_right.n0 drain_right.t10 3.3005
R133 drain_right.n11 drain_right.t14 3.3005
R134 drain_right.n11 drain_right.t11 3.3005
R135 drain_right.n12 drain_right.t16 3.3005
R136 drain_right.n12 drain_right.t15 3.3005
R137 drain_right.n14 drain_right.t13 3.3005
R138 drain_right.n14 drain_right.t17 3.3005
R139 drain_right.n16 drain_right.t12 3.3005
R140 drain_right.n16 drain_right.t22 3.3005
R141 drain_right.n18 drain_right.t23 3.3005
R142 drain_right.n18 drain_right.t8 3.3005
R143 drain_right.n20 drain_right.t19 3.3005
R144 drain_right.n20 drain_right.t5 3.3005
R145 drain_right.n9 drain_right.n7 0.457397
R146 drain_right.n4 drain_right.n2 0.457397
R147 drain_right.n21 drain_right.n19 0.457397
R148 drain_right.n19 drain_right.n17 0.457397
R149 drain_right.n17 drain_right.n15 0.457397
R150 drain_right.n15 drain_right.n13 0.457397
R151 drain_right.n10 drain_right.n9 0.173602
R152 drain_right.n10 drain_right.n4 0.173602
R153 source.n290 source.n264 289.615
R154 source.n248 source.n222 289.615
R155 source.n216 source.n190 289.615
R156 source.n174 source.n148 289.615
R157 source.n26 source.n0 289.615
R158 source.n68 source.n42 289.615
R159 source.n100 source.n74 289.615
R160 source.n142 source.n116 289.615
R161 source.n275 source.n274 185
R162 source.n272 source.n271 185
R163 source.n281 source.n280 185
R164 source.n283 source.n282 185
R165 source.n268 source.n267 185
R166 source.n289 source.n288 185
R167 source.n291 source.n290 185
R168 source.n233 source.n232 185
R169 source.n230 source.n229 185
R170 source.n239 source.n238 185
R171 source.n241 source.n240 185
R172 source.n226 source.n225 185
R173 source.n247 source.n246 185
R174 source.n249 source.n248 185
R175 source.n201 source.n200 185
R176 source.n198 source.n197 185
R177 source.n207 source.n206 185
R178 source.n209 source.n208 185
R179 source.n194 source.n193 185
R180 source.n215 source.n214 185
R181 source.n217 source.n216 185
R182 source.n159 source.n158 185
R183 source.n156 source.n155 185
R184 source.n165 source.n164 185
R185 source.n167 source.n166 185
R186 source.n152 source.n151 185
R187 source.n173 source.n172 185
R188 source.n175 source.n174 185
R189 source.n27 source.n26 185
R190 source.n25 source.n24 185
R191 source.n4 source.n3 185
R192 source.n19 source.n18 185
R193 source.n17 source.n16 185
R194 source.n8 source.n7 185
R195 source.n11 source.n10 185
R196 source.n69 source.n68 185
R197 source.n67 source.n66 185
R198 source.n46 source.n45 185
R199 source.n61 source.n60 185
R200 source.n59 source.n58 185
R201 source.n50 source.n49 185
R202 source.n53 source.n52 185
R203 source.n101 source.n100 185
R204 source.n99 source.n98 185
R205 source.n78 source.n77 185
R206 source.n93 source.n92 185
R207 source.n91 source.n90 185
R208 source.n82 source.n81 185
R209 source.n85 source.n84 185
R210 source.n143 source.n142 185
R211 source.n141 source.n140 185
R212 source.n120 source.n119 185
R213 source.n135 source.n134 185
R214 source.n133 source.n132 185
R215 source.n124 source.n123 185
R216 source.n127 source.n126 185
R217 source.t29 source.n273 147.661
R218 source.t32 source.n231 147.661
R219 source.t18 source.n199 147.661
R220 source.t4 source.n157 147.661
R221 source.t9 source.n9 147.661
R222 source.t5 source.n51 147.661
R223 source.t36 source.n83 147.661
R224 source.t42 source.n125 147.661
R225 source.n274 source.n271 104.615
R226 source.n281 source.n271 104.615
R227 source.n282 source.n281 104.615
R228 source.n282 source.n267 104.615
R229 source.n289 source.n267 104.615
R230 source.n290 source.n289 104.615
R231 source.n232 source.n229 104.615
R232 source.n239 source.n229 104.615
R233 source.n240 source.n239 104.615
R234 source.n240 source.n225 104.615
R235 source.n247 source.n225 104.615
R236 source.n248 source.n247 104.615
R237 source.n200 source.n197 104.615
R238 source.n207 source.n197 104.615
R239 source.n208 source.n207 104.615
R240 source.n208 source.n193 104.615
R241 source.n215 source.n193 104.615
R242 source.n216 source.n215 104.615
R243 source.n158 source.n155 104.615
R244 source.n165 source.n155 104.615
R245 source.n166 source.n165 104.615
R246 source.n166 source.n151 104.615
R247 source.n173 source.n151 104.615
R248 source.n174 source.n173 104.615
R249 source.n26 source.n25 104.615
R250 source.n25 source.n3 104.615
R251 source.n18 source.n3 104.615
R252 source.n18 source.n17 104.615
R253 source.n17 source.n7 104.615
R254 source.n10 source.n7 104.615
R255 source.n68 source.n67 104.615
R256 source.n67 source.n45 104.615
R257 source.n60 source.n45 104.615
R258 source.n60 source.n59 104.615
R259 source.n59 source.n49 104.615
R260 source.n52 source.n49 104.615
R261 source.n100 source.n99 104.615
R262 source.n99 source.n77 104.615
R263 source.n92 source.n77 104.615
R264 source.n92 source.n91 104.615
R265 source.n91 source.n81 104.615
R266 source.n84 source.n81 104.615
R267 source.n142 source.n141 104.615
R268 source.n141 source.n119 104.615
R269 source.n134 source.n119 104.615
R270 source.n134 source.n133 104.615
R271 source.n133 source.n123 104.615
R272 source.n126 source.n123 104.615
R273 source.n274 source.t29 52.3082
R274 source.n232 source.t32 52.3082
R275 source.n200 source.t18 52.3082
R276 source.n158 source.t4 52.3082
R277 source.n10 source.t9 52.3082
R278 source.n52 source.t5 52.3082
R279 source.n84 source.t36 52.3082
R280 source.n126 source.t42 52.3082
R281 source.n33 source.n32 50.512
R282 source.n35 source.n34 50.512
R283 source.n37 source.n36 50.512
R284 source.n39 source.n38 50.512
R285 source.n41 source.n40 50.512
R286 source.n107 source.n106 50.512
R287 source.n109 source.n108 50.512
R288 source.n111 source.n110 50.512
R289 source.n113 source.n112 50.512
R290 source.n115 source.n114 50.512
R291 source.n263 source.n262 50.5119
R292 source.n261 source.n260 50.5119
R293 source.n259 source.n258 50.5119
R294 source.n257 source.n256 50.5119
R295 source.n255 source.n254 50.5119
R296 source.n189 source.n188 50.5119
R297 source.n187 source.n186 50.5119
R298 source.n185 source.n184 50.5119
R299 source.n183 source.n182 50.5119
R300 source.n181 source.n180 50.5119
R301 source.n295 source.n294 32.1853
R302 source.n253 source.n252 32.1853
R303 source.n221 source.n220 32.1853
R304 source.n179 source.n178 32.1853
R305 source.n31 source.n30 32.1853
R306 source.n73 source.n72 32.1853
R307 source.n105 source.n104 32.1853
R308 source.n147 source.n146 32.1853
R309 source.n179 source.n147 17.1992
R310 source.n275 source.n273 15.6674
R311 source.n233 source.n231 15.6674
R312 source.n201 source.n199 15.6674
R313 source.n159 source.n157 15.6674
R314 source.n11 source.n9 15.6674
R315 source.n53 source.n51 15.6674
R316 source.n85 source.n83 15.6674
R317 source.n127 source.n125 15.6674
R318 source.n276 source.n272 12.8005
R319 source.n234 source.n230 12.8005
R320 source.n202 source.n198 12.8005
R321 source.n160 source.n156 12.8005
R322 source.n12 source.n8 12.8005
R323 source.n54 source.n50 12.8005
R324 source.n86 source.n82 12.8005
R325 source.n128 source.n124 12.8005
R326 source.n280 source.n279 12.0247
R327 source.n238 source.n237 12.0247
R328 source.n206 source.n205 12.0247
R329 source.n164 source.n163 12.0247
R330 source.n16 source.n15 12.0247
R331 source.n58 source.n57 12.0247
R332 source.n90 source.n89 12.0247
R333 source.n132 source.n131 12.0247
R334 source.n296 source.n31 11.7078
R335 source.n283 source.n270 11.249
R336 source.n241 source.n228 11.249
R337 source.n209 source.n196 11.249
R338 source.n167 source.n154 11.249
R339 source.n19 source.n6 11.249
R340 source.n61 source.n48 11.249
R341 source.n93 source.n80 11.249
R342 source.n135 source.n122 11.249
R343 source.n284 source.n268 10.4732
R344 source.n242 source.n226 10.4732
R345 source.n210 source.n194 10.4732
R346 source.n168 source.n152 10.4732
R347 source.n20 source.n4 10.4732
R348 source.n62 source.n46 10.4732
R349 source.n94 source.n78 10.4732
R350 source.n136 source.n120 10.4732
R351 source.n288 source.n287 9.69747
R352 source.n246 source.n245 9.69747
R353 source.n214 source.n213 9.69747
R354 source.n172 source.n171 9.69747
R355 source.n24 source.n23 9.69747
R356 source.n66 source.n65 9.69747
R357 source.n98 source.n97 9.69747
R358 source.n140 source.n139 9.69747
R359 source.n294 source.n293 9.45567
R360 source.n252 source.n251 9.45567
R361 source.n220 source.n219 9.45567
R362 source.n178 source.n177 9.45567
R363 source.n30 source.n29 9.45567
R364 source.n72 source.n71 9.45567
R365 source.n104 source.n103 9.45567
R366 source.n146 source.n145 9.45567
R367 source.n293 source.n292 9.3005
R368 source.n266 source.n265 9.3005
R369 source.n287 source.n286 9.3005
R370 source.n285 source.n284 9.3005
R371 source.n270 source.n269 9.3005
R372 source.n279 source.n278 9.3005
R373 source.n277 source.n276 9.3005
R374 source.n251 source.n250 9.3005
R375 source.n224 source.n223 9.3005
R376 source.n245 source.n244 9.3005
R377 source.n243 source.n242 9.3005
R378 source.n228 source.n227 9.3005
R379 source.n237 source.n236 9.3005
R380 source.n235 source.n234 9.3005
R381 source.n219 source.n218 9.3005
R382 source.n192 source.n191 9.3005
R383 source.n213 source.n212 9.3005
R384 source.n211 source.n210 9.3005
R385 source.n196 source.n195 9.3005
R386 source.n205 source.n204 9.3005
R387 source.n203 source.n202 9.3005
R388 source.n177 source.n176 9.3005
R389 source.n150 source.n149 9.3005
R390 source.n171 source.n170 9.3005
R391 source.n169 source.n168 9.3005
R392 source.n154 source.n153 9.3005
R393 source.n163 source.n162 9.3005
R394 source.n161 source.n160 9.3005
R395 source.n29 source.n28 9.3005
R396 source.n2 source.n1 9.3005
R397 source.n23 source.n22 9.3005
R398 source.n21 source.n20 9.3005
R399 source.n6 source.n5 9.3005
R400 source.n15 source.n14 9.3005
R401 source.n13 source.n12 9.3005
R402 source.n71 source.n70 9.3005
R403 source.n44 source.n43 9.3005
R404 source.n65 source.n64 9.3005
R405 source.n63 source.n62 9.3005
R406 source.n48 source.n47 9.3005
R407 source.n57 source.n56 9.3005
R408 source.n55 source.n54 9.3005
R409 source.n103 source.n102 9.3005
R410 source.n76 source.n75 9.3005
R411 source.n97 source.n96 9.3005
R412 source.n95 source.n94 9.3005
R413 source.n80 source.n79 9.3005
R414 source.n89 source.n88 9.3005
R415 source.n87 source.n86 9.3005
R416 source.n145 source.n144 9.3005
R417 source.n118 source.n117 9.3005
R418 source.n139 source.n138 9.3005
R419 source.n137 source.n136 9.3005
R420 source.n122 source.n121 9.3005
R421 source.n131 source.n130 9.3005
R422 source.n129 source.n128 9.3005
R423 source.n291 source.n266 8.92171
R424 source.n249 source.n224 8.92171
R425 source.n217 source.n192 8.92171
R426 source.n175 source.n150 8.92171
R427 source.n27 source.n2 8.92171
R428 source.n69 source.n44 8.92171
R429 source.n101 source.n76 8.92171
R430 source.n143 source.n118 8.92171
R431 source.n292 source.n264 8.14595
R432 source.n250 source.n222 8.14595
R433 source.n218 source.n190 8.14595
R434 source.n176 source.n148 8.14595
R435 source.n28 source.n0 8.14595
R436 source.n70 source.n42 8.14595
R437 source.n102 source.n74 8.14595
R438 source.n144 source.n116 8.14595
R439 source.n294 source.n264 5.81868
R440 source.n252 source.n222 5.81868
R441 source.n220 source.n190 5.81868
R442 source.n178 source.n148 5.81868
R443 source.n30 source.n0 5.81868
R444 source.n72 source.n42 5.81868
R445 source.n104 source.n74 5.81868
R446 source.n146 source.n116 5.81868
R447 source.n296 source.n295 5.49188
R448 source.n292 source.n291 5.04292
R449 source.n250 source.n249 5.04292
R450 source.n218 source.n217 5.04292
R451 source.n176 source.n175 5.04292
R452 source.n28 source.n27 5.04292
R453 source.n70 source.n69 5.04292
R454 source.n102 source.n101 5.04292
R455 source.n144 source.n143 5.04292
R456 source.n277 source.n273 4.38594
R457 source.n235 source.n231 4.38594
R458 source.n203 source.n199 4.38594
R459 source.n161 source.n157 4.38594
R460 source.n13 source.n9 4.38594
R461 source.n55 source.n51 4.38594
R462 source.n87 source.n83 4.38594
R463 source.n129 source.n125 4.38594
R464 source.n288 source.n266 4.26717
R465 source.n246 source.n224 4.26717
R466 source.n214 source.n192 4.26717
R467 source.n172 source.n150 4.26717
R468 source.n24 source.n2 4.26717
R469 source.n66 source.n44 4.26717
R470 source.n98 source.n76 4.26717
R471 source.n140 source.n118 4.26717
R472 source.n287 source.n268 3.49141
R473 source.n245 source.n226 3.49141
R474 source.n213 source.n194 3.49141
R475 source.n171 source.n152 3.49141
R476 source.n23 source.n4 3.49141
R477 source.n65 source.n46 3.49141
R478 source.n97 source.n78 3.49141
R479 source.n139 source.n120 3.49141
R480 source.n262 source.t28 3.3005
R481 source.n262 source.t34 3.3005
R482 source.n260 source.t25 3.3005
R483 source.n260 source.t47 3.3005
R484 source.n258 source.t24 3.3005
R485 source.n258 source.t46 3.3005
R486 source.n256 source.t27 3.3005
R487 source.n256 source.t43 3.3005
R488 source.n254 source.t26 3.3005
R489 source.n254 source.t33 3.3005
R490 source.n188 source.t13 3.3005
R491 source.n188 source.t23 3.3005
R492 source.n186 source.t6 3.3005
R493 source.n186 source.t0 3.3005
R494 source.n184 source.t7 3.3005
R495 source.n184 source.t11 3.3005
R496 source.n182 source.t16 3.3005
R497 source.n182 source.t17 3.3005
R498 source.n180 source.t8 3.3005
R499 source.n180 source.t22 3.3005
R500 source.n32 source.t1 3.3005
R501 source.n32 source.t21 3.3005
R502 source.n34 source.t14 3.3005
R503 source.n34 source.t12 3.3005
R504 source.n36 source.t10 3.3005
R505 source.n36 source.t15 3.3005
R506 source.n38 source.t3 3.3005
R507 source.n38 source.t2 3.3005
R508 source.n40 source.t20 3.3005
R509 source.n40 source.t19 3.3005
R510 source.n106 source.t45 3.3005
R511 source.n106 source.t40 3.3005
R512 source.n108 source.t35 3.3005
R513 source.n108 source.t31 3.3005
R514 source.n110 source.t44 3.3005
R515 source.n110 source.t41 3.3005
R516 source.n112 source.t37 3.3005
R517 source.n112 source.t30 3.3005
R518 source.n114 source.t38 3.3005
R519 source.n114 source.t39 3.3005
R520 source.n284 source.n283 2.71565
R521 source.n242 source.n241 2.71565
R522 source.n210 source.n209 2.71565
R523 source.n168 source.n167 2.71565
R524 source.n20 source.n19 2.71565
R525 source.n62 source.n61 2.71565
R526 source.n94 source.n93 2.71565
R527 source.n136 source.n135 2.71565
R528 source.n280 source.n270 1.93989
R529 source.n238 source.n228 1.93989
R530 source.n206 source.n196 1.93989
R531 source.n164 source.n154 1.93989
R532 source.n16 source.n6 1.93989
R533 source.n58 source.n48 1.93989
R534 source.n90 source.n80 1.93989
R535 source.n132 source.n122 1.93989
R536 source.n279 source.n272 1.16414
R537 source.n237 source.n230 1.16414
R538 source.n205 source.n198 1.16414
R539 source.n163 source.n156 1.16414
R540 source.n15 source.n8 1.16414
R541 source.n57 source.n50 1.16414
R542 source.n89 source.n82 1.16414
R543 source.n131 source.n124 1.16414
R544 source.n105 source.n73 0.470328
R545 source.n253 source.n221 0.470328
R546 source.n147 source.n115 0.457397
R547 source.n115 source.n113 0.457397
R548 source.n113 source.n111 0.457397
R549 source.n111 source.n109 0.457397
R550 source.n109 source.n107 0.457397
R551 source.n107 source.n105 0.457397
R552 source.n73 source.n41 0.457397
R553 source.n41 source.n39 0.457397
R554 source.n39 source.n37 0.457397
R555 source.n37 source.n35 0.457397
R556 source.n35 source.n33 0.457397
R557 source.n33 source.n31 0.457397
R558 source.n181 source.n179 0.457397
R559 source.n183 source.n181 0.457397
R560 source.n185 source.n183 0.457397
R561 source.n187 source.n185 0.457397
R562 source.n189 source.n187 0.457397
R563 source.n221 source.n189 0.457397
R564 source.n255 source.n253 0.457397
R565 source.n257 source.n255 0.457397
R566 source.n259 source.n257 0.457397
R567 source.n261 source.n259 0.457397
R568 source.n263 source.n261 0.457397
R569 source.n295 source.n263 0.457397
R570 source.n276 source.n275 0.388379
R571 source.n234 source.n233 0.388379
R572 source.n202 source.n201 0.388379
R573 source.n160 source.n159 0.388379
R574 source.n12 source.n11 0.388379
R575 source.n54 source.n53 0.388379
R576 source.n86 source.n85 0.388379
R577 source.n128 source.n127 0.388379
R578 source source.n296 0.188
R579 source.n278 source.n277 0.155672
R580 source.n278 source.n269 0.155672
R581 source.n285 source.n269 0.155672
R582 source.n286 source.n285 0.155672
R583 source.n286 source.n265 0.155672
R584 source.n293 source.n265 0.155672
R585 source.n236 source.n235 0.155672
R586 source.n236 source.n227 0.155672
R587 source.n243 source.n227 0.155672
R588 source.n244 source.n243 0.155672
R589 source.n244 source.n223 0.155672
R590 source.n251 source.n223 0.155672
R591 source.n204 source.n203 0.155672
R592 source.n204 source.n195 0.155672
R593 source.n211 source.n195 0.155672
R594 source.n212 source.n211 0.155672
R595 source.n212 source.n191 0.155672
R596 source.n219 source.n191 0.155672
R597 source.n162 source.n161 0.155672
R598 source.n162 source.n153 0.155672
R599 source.n169 source.n153 0.155672
R600 source.n170 source.n169 0.155672
R601 source.n170 source.n149 0.155672
R602 source.n177 source.n149 0.155672
R603 source.n29 source.n1 0.155672
R604 source.n22 source.n1 0.155672
R605 source.n22 source.n21 0.155672
R606 source.n21 source.n5 0.155672
R607 source.n14 source.n5 0.155672
R608 source.n14 source.n13 0.155672
R609 source.n71 source.n43 0.155672
R610 source.n64 source.n43 0.155672
R611 source.n64 source.n63 0.155672
R612 source.n63 source.n47 0.155672
R613 source.n56 source.n47 0.155672
R614 source.n56 source.n55 0.155672
R615 source.n103 source.n75 0.155672
R616 source.n96 source.n75 0.155672
R617 source.n96 source.n95 0.155672
R618 source.n95 source.n79 0.155672
R619 source.n88 source.n79 0.155672
R620 source.n88 source.n87 0.155672
R621 source.n145 source.n117 0.155672
R622 source.n138 source.n117 0.155672
R623 source.n138 source.n137 0.155672
R624 source.n137 source.n121 0.155672
R625 source.n130 source.n121 0.155672
R626 source.n130 source.n129 0.155672
R627 plus.n6 plus.t13 940.265
R628 plus.n29 plus.t21 940.265
R629 plus.n37 plus.t16 940.265
R630 plus.n60 plus.t10 940.265
R631 plus.n7 plus.t4 879.65
R632 plus.n5 plus.t23 879.65
R633 plus.n12 plus.t20 879.65
R634 plus.n14 plus.t19 879.65
R635 plus.n3 plus.t12 879.65
R636 plus.n19 plus.t3 879.65
R637 plus.n21 plus.t22 879.65
R638 plus.n1 plus.t18 879.65
R639 plus.n26 plus.t9 879.65
R640 plus.n28 plus.t1 879.65
R641 plus.n38 plus.t17 879.65
R642 plus.n36 plus.t14 879.65
R643 plus.n43 plus.t8 879.65
R644 plus.n45 plus.t15 879.65
R645 plus.n34 plus.t7 879.65
R646 plus.n50 plus.t11 879.65
R647 plus.n52 plus.t5 879.65
R648 plus.n32 plus.t2 879.65
R649 plus.n57 plus.t0 879.65
R650 plus.n59 plus.t6 879.65
R651 plus.n9 plus.n6 161.489
R652 plus.n40 plus.n37 161.489
R653 plus.n9 plus.n8 161.3
R654 plus.n11 plus.n10 161.3
R655 plus.n13 plus.n4 161.3
R656 plus.n16 plus.n15 161.3
R657 plus.n18 plus.n17 161.3
R658 plus.n20 plus.n2 161.3
R659 plus.n23 plus.n22 161.3
R660 plus.n25 plus.n24 161.3
R661 plus.n27 plus.n0 161.3
R662 plus.n30 plus.n29 161.3
R663 plus.n40 plus.n39 161.3
R664 plus.n42 plus.n41 161.3
R665 plus.n44 plus.n35 161.3
R666 plus.n47 plus.n46 161.3
R667 plus.n49 plus.n48 161.3
R668 plus.n51 plus.n33 161.3
R669 plus.n54 plus.n53 161.3
R670 plus.n56 plus.n55 161.3
R671 plus.n58 plus.n31 161.3
R672 plus.n61 plus.n60 161.3
R673 plus.n8 plus.n7 56.2338
R674 plus.n28 plus.n27 56.2338
R675 plus.n59 plus.n58 56.2338
R676 plus.n39 plus.n38 56.2338
R677 plus.n11 plus.n5 51.852
R678 plus.n26 plus.n25 51.852
R679 plus.n57 plus.n56 51.852
R680 plus.n42 plus.n36 51.852
R681 plus.n13 plus.n12 47.4702
R682 plus.n22 plus.n1 47.4702
R683 plus.n53 plus.n32 47.4702
R684 plus.n44 plus.n43 47.4702
R685 plus.n15 plus.n14 43.0884
R686 plus.n21 plus.n20 43.0884
R687 plus.n52 plus.n51 43.0884
R688 plus.n46 plus.n45 43.0884
R689 plus.n18 plus.n3 38.7066
R690 plus.n19 plus.n18 38.7066
R691 plus.n50 plus.n49 38.7066
R692 plus.n49 plus.n34 38.7066
R693 plus.n15 plus.n3 34.3247
R694 plus.n20 plus.n19 34.3247
R695 plus.n51 plus.n50 34.3247
R696 plus.n46 plus.n34 34.3247
R697 plus.n14 plus.n13 29.9429
R698 plus.n22 plus.n21 29.9429
R699 plus.n53 plus.n52 29.9429
R700 plus.n45 plus.n44 29.9429
R701 plus plus.n61 28.6505
R702 plus.n12 plus.n11 25.5611
R703 plus.n25 plus.n1 25.5611
R704 plus.n56 plus.n32 25.5611
R705 plus.n43 plus.n42 25.5611
R706 plus.n8 plus.n5 21.1793
R707 plus.n27 plus.n26 21.1793
R708 plus.n58 plus.n57 21.1793
R709 plus.n39 plus.n36 21.1793
R710 plus.n7 plus.n6 16.7975
R711 plus.n29 plus.n28 16.7975
R712 plus.n60 plus.n59 16.7975
R713 plus.n38 plus.n37 16.7975
R714 plus plus.n30 9.86035
R715 plus.n10 plus.n9 0.189894
R716 plus.n10 plus.n4 0.189894
R717 plus.n16 plus.n4 0.189894
R718 plus.n17 plus.n16 0.189894
R719 plus.n17 plus.n2 0.189894
R720 plus.n23 plus.n2 0.189894
R721 plus.n24 plus.n23 0.189894
R722 plus.n24 plus.n0 0.189894
R723 plus.n30 plus.n0 0.189894
R724 plus.n61 plus.n31 0.189894
R725 plus.n55 plus.n31 0.189894
R726 plus.n55 plus.n54 0.189894
R727 plus.n54 plus.n33 0.189894
R728 plus.n48 plus.n33 0.189894
R729 plus.n48 plus.n47 0.189894
R730 plus.n47 plus.n35 0.189894
R731 plus.n41 plus.n35 0.189894
R732 plus.n41 plus.n40 0.189894
R733 drain_left.n13 drain_left.n11 67.6477
R734 drain_left.n7 drain_left.n5 67.6476
R735 drain_left.n2 drain_left.n0 67.6476
R736 drain_left.n19 drain_left.n18 67.1908
R737 drain_left.n17 drain_left.n16 67.1908
R738 drain_left.n15 drain_left.n14 67.1908
R739 drain_left.n13 drain_left.n12 67.1908
R740 drain_left.n21 drain_left.n20 67.1907
R741 drain_left.n7 drain_left.n6 67.1907
R742 drain_left.n9 drain_left.n8 67.1907
R743 drain_left.n4 drain_left.n3 67.1907
R744 drain_left.n2 drain_left.n1 67.1907
R745 drain_left drain_left.n10 27.1621
R746 drain_left drain_left.n21 6.11011
R747 drain_left.n5 drain_left.t6 3.3005
R748 drain_left.n5 drain_left.t7 3.3005
R749 drain_left.n6 drain_left.t15 3.3005
R750 drain_left.n6 drain_left.t9 3.3005
R751 drain_left.n8 drain_left.t16 3.3005
R752 drain_left.n8 drain_left.t8 3.3005
R753 drain_left.n3 drain_left.t18 3.3005
R754 drain_left.n3 drain_left.t12 3.3005
R755 drain_left.n1 drain_left.t23 3.3005
R756 drain_left.n1 drain_left.t21 3.3005
R757 drain_left.n0 drain_left.t13 3.3005
R758 drain_left.n0 drain_left.t17 3.3005
R759 drain_left.n20 drain_left.t22 3.3005
R760 drain_left.n20 drain_left.t2 3.3005
R761 drain_left.n18 drain_left.t5 3.3005
R762 drain_left.n18 drain_left.t14 3.3005
R763 drain_left.n16 drain_left.t20 3.3005
R764 drain_left.n16 drain_left.t1 3.3005
R765 drain_left.n14 drain_left.t4 3.3005
R766 drain_left.n14 drain_left.t11 3.3005
R767 drain_left.n12 drain_left.t0 3.3005
R768 drain_left.n12 drain_left.t3 3.3005
R769 drain_left.n11 drain_left.t10 3.3005
R770 drain_left.n11 drain_left.t19 3.3005
R771 drain_left.n9 drain_left.n7 0.457397
R772 drain_left.n4 drain_left.n2 0.457397
R773 drain_left.n15 drain_left.n13 0.457397
R774 drain_left.n17 drain_left.n15 0.457397
R775 drain_left.n19 drain_left.n17 0.457397
R776 drain_left.n21 drain_left.n19 0.457397
R777 drain_left.n10 drain_left.n9 0.173602
R778 drain_left.n10 drain_left.n4 0.173602
C0 plus minus 4.655f
C1 drain_right source 28.693699f
C2 drain_right minus 3.43471f
C3 drain_right plus 0.359911f
C4 drain_left source 28.693499f
C5 drain_left minus 0.171754f
C6 minus source 3.42992f
C7 drain_left plus 3.63986f
C8 drain_right drain_left 1.11966f
C9 plus source 3.44394f
C10 drain_right a_n2094_n2088# 5.99983f
C11 drain_left a_n2094_n2088# 6.32922f
C12 source a_n2094_n2088# 5.413197f
C13 minus a_n2094_n2088# 7.67265f
C14 plus a_n2094_n2088# 9.37445f
C15 drain_left.t13 a_n2094_n2088# 0.181597f
C16 drain_left.t17 a_n2094_n2088# 0.181597f
C17 drain_left.n0 a_n2094_n2088# 1.51748f
C18 drain_left.t23 a_n2094_n2088# 0.181597f
C19 drain_left.t21 a_n2094_n2088# 0.181597f
C20 drain_left.n1 a_n2094_n2088# 1.51452f
C21 drain_left.n2 a_n2094_n2088# 0.859726f
C22 drain_left.t18 a_n2094_n2088# 0.181597f
C23 drain_left.t12 a_n2094_n2088# 0.181597f
C24 drain_left.n3 a_n2094_n2088# 1.51452f
C25 drain_left.n4 a_n2094_n2088# 0.393739f
C26 drain_left.t6 a_n2094_n2088# 0.181597f
C27 drain_left.t7 a_n2094_n2088# 0.181597f
C28 drain_left.n5 a_n2094_n2088# 1.51748f
C29 drain_left.t15 a_n2094_n2088# 0.181597f
C30 drain_left.t9 a_n2094_n2088# 0.181597f
C31 drain_left.n6 a_n2094_n2088# 1.51452f
C32 drain_left.n7 a_n2094_n2088# 0.859726f
C33 drain_left.t16 a_n2094_n2088# 0.181597f
C34 drain_left.t8 a_n2094_n2088# 0.181597f
C35 drain_left.n8 a_n2094_n2088# 1.51452f
C36 drain_left.n9 a_n2094_n2088# 0.393739f
C37 drain_left.n10 a_n2094_n2088# 1.46318f
C38 drain_left.t10 a_n2094_n2088# 0.181597f
C39 drain_left.t19 a_n2094_n2088# 0.181597f
C40 drain_left.n11 a_n2094_n2088# 1.51749f
C41 drain_left.t0 a_n2094_n2088# 0.181597f
C42 drain_left.t3 a_n2094_n2088# 0.181597f
C43 drain_left.n12 a_n2094_n2088# 1.51452f
C44 drain_left.n13 a_n2094_n2088# 0.859712f
C45 drain_left.t4 a_n2094_n2088# 0.181597f
C46 drain_left.t11 a_n2094_n2088# 0.181597f
C47 drain_left.n14 a_n2094_n2088# 1.51452f
C48 drain_left.n15 a_n2094_n2088# 0.423626f
C49 drain_left.t20 a_n2094_n2088# 0.181597f
C50 drain_left.t1 a_n2094_n2088# 0.181597f
C51 drain_left.n16 a_n2094_n2088# 1.51452f
C52 drain_left.n17 a_n2094_n2088# 0.423626f
C53 drain_left.t5 a_n2094_n2088# 0.181597f
C54 drain_left.t14 a_n2094_n2088# 0.181597f
C55 drain_left.n18 a_n2094_n2088# 1.51452f
C56 drain_left.n19 a_n2094_n2088# 0.423626f
C57 drain_left.t22 a_n2094_n2088# 0.181597f
C58 drain_left.t2 a_n2094_n2088# 0.181597f
C59 drain_left.n20 a_n2094_n2088# 1.51452f
C60 drain_left.n21 a_n2094_n2088# 0.737085f
C61 plus.n0 a_n2094_n2088# 0.052655f
C62 plus.t1 a_n2094_n2088# 0.180028f
C63 plus.t9 a_n2094_n2088# 0.180028f
C64 plus.t18 a_n2094_n2088# 0.180028f
C65 plus.n1 a_n2094_n2088# 0.088046f
C66 plus.n2 a_n2094_n2088# 0.052655f
C67 plus.t22 a_n2094_n2088# 0.180028f
C68 plus.t3 a_n2094_n2088# 0.180028f
C69 plus.t12 a_n2094_n2088# 0.180028f
C70 plus.n3 a_n2094_n2088# 0.088046f
C71 plus.n4 a_n2094_n2088# 0.052655f
C72 plus.t19 a_n2094_n2088# 0.180028f
C73 plus.t20 a_n2094_n2088# 0.180028f
C74 plus.t23 a_n2094_n2088# 0.180028f
C75 plus.n5 a_n2094_n2088# 0.088046f
C76 plus.t13 a_n2094_n2088# 0.185944f
C77 plus.n6 a_n2094_n2088# 0.104386f
C78 plus.t4 a_n2094_n2088# 0.180028f
C79 plus.n7 a_n2094_n2088# 0.088046f
C80 plus.n8 a_n2094_n2088# 0.018441f
C81 plus.n9 a_n2094_n2088# 0.122434f
C82 plus.n10 a_n2094_n2088# 0.052655f
C83 plus.n11 a_n2094_n2088# 0.018441f
C84 plus.n12 a_n2094_n2088# 0.088046f
C85 plus.n13 a_n2094_n2088# 0.018441f
C86 plus.n14 a_n2094_n2088# 0.088046f
C87 plus.n15 a_n2094_n2088# 0.018441f
C88 plus.n16 a_n2094_n2088# 0.052655f
C89 plus.n17 a_n2094_n2088# 0.052655f
C90 plus.n18 a_n2094_n2088# 0.018441f
C91 plus.n19 a_n2094_n2088# 0.088046f
C92 plus.n20 a_n2094_n2088# 0.018441f
C93 plus.n21 a_n2094_n2088# 0.088046f
C94 plus.n22 a_n2094_n2088# 0.018441f
C95 plus.n23 a_n2094_n2088# 0.052655f
C96 plus.n24 a_n2094_n2088# 0.052655f
C97 plus.n25 a_n2094_n2088# 0.018441f
C98 plus.n26 a_n2094_n2088# 0.088046f
C99 plus.n27 a_n2094_n2088# 0.018441f
C100 plus.n28 a_n2094_n2088# 0.088046f
C101 plus.t21 a_n2094_n2088# 0.185944f
C102 plus.n29 a_n2094_n2088# 0.104304f
C103 plus.n30 a_n2094_n2088# 0.44979f
C104 plus.n31 a_n2094_n2088# 0.052655f
C105 plus.t10 a_n2094_n2088# 0.185944f
C106 plus.t6 a_n2094_n2088# 0.180028f
C107 plus.t0 a_n2094_n2088# 0.180028f
C108 plus.t2 a_n2094_n2088# 0.180028f
C109 plus.n32 a_n2094_n2088# 0.088046f
C110 plus.n33 a_n2094_n2088# 0.052655f
C111 plus.t5 a_n2094_n2088# 0.180028f
C112 plus.t11 a_n2094_n2088# 0.180028f
C113 plus.t7 a_n2094_n2088# 0.180028f
C114 plus.n34 a_n2094_n2088# 0.088046f
C115 plus.n35 a_n2094_n2088# 0.052655f
C116 plus.t15 a_n2094_n2088# 0.180028f
C117 plus.t8 a_n2094_n2088# 0.180028f
C118 plus.t14 a_n2094_n2088# 0.180028f
C119 plus.n36 a_n2094_n2088# 0.088046f
C120 plus.t16 a_n2094_n2088# 0.185944f
C121 plus.n37 a_n2094_n2088# 0.104386f
C122 plus.t17 a_n2094_n2088# 0.180028f
C123 plus.n38 a_n2094_n2088# 0.088046f
C124 plus.n39 a_n2094_n2088# 0.018441f
C125 plus.n40 a_n2094_n2088# 0.122434f
C126 plus.n41 a_n2094_n2088# 0.052655f
C127 plus.n42 a_n2094_n2088# 0.018441f
C128 plus.n43 a_n2094_n2088# 0.088046f
C129 plus.n44 a_n2094_n2088# 0.018441f
C130 plus.n45 a_n2094_n2088# 0.088046f
C131 plus.n46 a_n2094_n2088# 0.018441f
C132 plus.n47 a_n2094_n2088# 0.052655f
C133 plus.n48 a_n2094_n2088# 0.052655f
C134 plus.n49 a_n2094_n2088# 0.018441f
C135 plus.n50 a_n2094_n2088# 0.088046f
C136 plus.n51 a_n2094_n2088# 0.018441f
C137 plus.n52 a_n2094_n2088# 0.088046f
C138 plus.n53 a_n2094_n2088# 0.018441f
C139 plus.n54 a_n2094_n2088# 0.052655f
C140 plus.n55 a_n2094_n2088# 0.052655f
C141 plus.n56 a_n2094_n2088# 0.018441f
C142 plus.n57 a_n2094_n2088# 0.088046f
C143 plus.n58 a_n2094_n2088# 0.018441f
C144 plus.n59 a_n2094_n2088# 0.088046f
C145 plus.n60 a_n2094_n2088# 0.104304f
C146 plus.n61 a_n2094_n2088# 1.41422f
C147 source.n0 a_n2094_n2088# 0.04998f
C148 source.n1 a_n2094_n2088# 0.035558f
C149 source.n2 a_n2094_n2088# 0.019108f
C150 source.n3 a_n2094_n2088# 0.045163f
C151 source.n4 a_n2094_n2088# 0.020232f
C152 source.n5 a_n2094_n2088# 0.035558f
C153 source.n6 a_n2094_n2088# 0.019108f
C154 source.n7 a_n2094_n2088# 0.045163f
C155 source.n8 a_n2094_n2088# 0.020232f
C156 source.n9 a_n2094_n2088# 0.152165f
C157 source.t9 a_n2094_n2088# 0.07361f
C158 source.n10 a_n2094_n2088# 0.033872f
C159 source.n11 a_n2094_n2088# 0.026678f
C160 source.n12 a_n2094_n2088# 0.019108f
C161 source.n13 a_n2094_n2088# 0.846075f
C162 source.n14 a_n2094_n2088# 0.035558f
C163 source.n15 a_n2094_n2088# 0.019108f
C164 source.n16 a_n2094_n2088# 0.020232f
C165 source.n17 a_n2094_n2088# 0.045163f
C166 source.n18 a_n2094_n2088# 0.045163f
C167 source.n19 a_n2094_n2088# 0.020232f
C168 source.n20 a_n2094_n2088# 0.019108f
C169 source.n21 a_n2094_n2088# 0.035558f
C170 source.n22 a_n2094_n2088# 0.035558f
C171 source.n23 a_n2094_n2088# 0.019108f
C172 source.n24 a_n2094_n2088# 0.020232f
C173 source.n25 a_n2094_n2088# 0.045163f
C174 source.n26 a_n2094_n2088# 0.097771f
C175 source.n27 a_n2094_n2088# 0.020232f
C176 source.n28 a_n2094_n2088# 0.019108f
C177 source.n29 a_n2094_n2088# 0.082191f
C178 source.n30 a_n2094_n2088# 0.054706f
C179 source.n31 a_n2094_n2088# 0.84435f
C180 source.t1 a_n2094_n2088# 0.168595f
C181 source.t21 a_n2094_n2088# 0.168595f
C182 source.n32 a_n2094_n2088# 1.31304f
C183 source.n33 a_n2094_n2088# 0.438024f
C184 source.t14 a_n2094_n2088# 0.168595f
C185 source.t12 a_n2094_n2088# 0.168595f
C186 source.n34 a_n2094_n2088# 1.31304f
C187 source.n35 a_n2094_n2088# 0.438024f
C188 source.t10 a_n2094_n2088# 0.168595f
C189 source.t15 a_n2094_n2088# 0.168595f
C190 source.n36 a_n2094_n2088# 1.31304f
C191 source.n37 a_n2094_n2088# 0.438024f
C192 source.t3 a_n2094_n2088# 0.168595f
C193 source.t2 a_n2094_n2088# 0.168595f
C194 source.n38 a_n2094_n2088# 1.31304f
C195 source.n39 a_n2094_n2088# 0.438024f
C196 source.t20 a_n2094_n2088# 0.168595f
C197 source.t19 a_n2094_n2088# 0.168595f
C198 source.n40 a_n2094_n2088# 1.31304f
C199 source.n41 a_n2094_n2088# 0.438024f
C200 source.n42 a_n2094_n2088# 0.04998f
C201 source.n43 a_n2094_n2088# 0.035558f
C202 source.n44 a_n2094_n2088# 0.019108f
C203 source.n45 a_n2094_n2088# 0.045163f
C204 source.n46 a_n2094_n2088# 0.020232f
C205 source.n47 a_n2094_n2088# 0.035558f
C206 source.n48 a_n2094_n2088# 0.019108f
C207 source.n49 a_n2094_n2088# 0.045163f
C208 source.n50 a_n2094_n2088# 0.020232f
C209 source.n51 a_n2094_n2088# 0.152165f
C210 source.t5 a_n2094_n2088# 0.07361f
C211 source.n52 a_n2094_n2088# 0.033872f
C212 source.n53 a_n2094_n2088# 0.026678f
C213 source.n54 a_n2094_n2088# 0.019108f
C214 source.n55 a_n2094_n2088# 0.846075f
C215 source.n56 a_n2094_n2088# 0.035558f
C216 source.n57 a_n2094_n2088# 0.019108f
C217 source.n58 a_n2094_n2088# 0.020232f
C218 source.n59 a_n2094_n2088# 0.045163f
C219 source.n60 a_n2094_n2088# 0.045163f
C220 source.n61 a_n2094_n2088# 0.020232f
C221 source.n62 a_n2094_n2088# 0.019108f
C222 source.n63 a_n2094_n2088# 0.035558f
C223 source.n64 a_n2094_n2088# 0.035558f
C224 source.n65 a_n2094_n2088# 0.019108f
C225 source.n66 a_n2094_n2088# 0.020232f
C226 source.n67 a_n2094_n2088# 0.045163f
C227 source.n68 a_n2094_n2088# 0.097771f
C228 source.n69 a_n2094_n2088# 0.020232f
C229 source.n70 a_n2094_n2088# 0.019108f
C230 source.n71 a_n2094_n2088# 0.082191f
C231 source.n72 a_n2094_n2088# 0.054706f
C232 source.n73 a_n2094_n2088# 0.13655f
C233 source.n74 a_n2094_n2088# 0.04998f
C234 source.n75 a_n2094_n2088# 0.035558f
C235 source.n76 a_n2094_n2088# 0.019108f
C236 source.n77 a_n2094_n2088# 0.045163f
C237 source.n78 a_n2094_n2088# 0.020232f
C238 source.n79 a_n2094_n2088# 0.035558f
C239 source.n80 a_n2094_n2088# 0.019108f
C240 source.n81 a_n2094_n2088# 0.045163f
C241 source.n82 a_n2094_n2088# 0.020232f
C242 source.n83 a_n2094_n2088# 0.152165f
C243 source.t36 a_n2094_n2088# 0.07361f
C244 source.n84 a_n2094_n2088# 0.033872f
C245 source.n85 a_n2094_n2088# 0.026678f
C246 source.n86 a_n2094_n2088# 0.019108f
C247 source.n87 a_n2094_n2088# 0.846075f
C248 source.n88 a_n2094_n2088# 0.035558f
C249 source.n89 a_n2094_n2088# 0.019108f
C250 source.n90 a_n2094_n2088# 0.020232f
C251 source.n91 a_n2094_n2088# 0.045163f
C252 source.n92 a_n2094_n2088# 0.045163f
C253 source.n93 a_n2094_n2088# 0.020232f
C254 source.n94 a_n2094_n2088# 0.019108f
C255 source.n95 a_n2094_n2088# 0.035558f
C256 source.n96 a_n2094_n2088# 0.035558f
C257 source.n97 a_n2094_n2088# 0.019108f
C258 source.n98 a_n2094_n2088# 0.020232f
C259 source.n99 a_n2094_n2088# 0.045163f
C260 source.n100 a_n2094_n2088# 0.097771f
C261 source.n101 a_n2094_n2088# 0.020232f
C262 source.n102 a_n2094_n2088# 0.019108f
C263 source.n103 a_n2094_n2088# 0.082191f
C264 source.n104 a_n2094_n2088# 0.054706f
C265 source.n105 a_n2094_n2088# 0.13655f
C266 source.t45 a_n2094_n2088# 0.168595f
C267 source.t40 a_n2094_n2088# 0.168595f
C268 source.n106 a_n2094_n2088# 1.31304f
C269 source.n107 a_n2094_n2088# 0.438024f
C270 source.t35 a_n2094_n2088# 0.168595f
C271 source.t31 a_n2094_n2088# 0.168595f
C272 source.n108 a_n2094_n2088# 1.31304f
C273 source.n109 a_n2094_n2088# 0.438024f
C274 source.t44 a_n2094_n2088# 0.168595f
C275 source.t41 a_n2094_n2088# 0.168595f
C276 source.n110 a_n2094_n2088# 1.31304f
C277 source.n111 a_n2094_n2088# 0.438024f
C278 source.t37 a_n2094_n2088# 0.168595f
C279 source.t30 a_n2094_n2088# 0.168595f
C280 source.n112 a_n2094_n2088# 1.31304f
C281 source.n113 a_n2094_n2088# 0.438024f
C282 source.t38 a_n2094_n2088# 0.168595f
C283 source.t39 a_n2094_n2088# 0.168595f
C284 source.n114 a_n2094_n2088# 1.31304f
C285 source.n115 a_n2094_n2088# 0.438024f
C286 source.n116 a_n2094_n2088# 0.04998f
C287 source.n117 a_n2094_n2088# 0.035558f
C288 source.n118 a_n2094_n2088# 0.019108f
C289 source.n119 a_n2094_n2088# 0.045163f
C290 source.n120 a_n2094_n2088# 0.020232f
C291 source.n121 a_n2094_n2088# 0.035558f
C292 source.n122 a_n2094_n2088# 0.019108f
C293 source.n123 a_n2094_n2088# 0.045163f
C294 source.n124 a_n2094_n2088# 0.020232f
C295 source.n125 a_n2094_n2088# 0.152165f
C296 source.t42 a_n2094_n2088# 0.07361f
C297 source.n126 a_n2094_n2088# 0.033872f
C298 source.n127 a_n2094_n2088# 0.026678f
C299 source.n128 a_n2094_n2088# 0.019108f
C300 source.n129 a_n2094_n2088# 0.846075f
C301 source.n130 a_n2094_n2088# 0.035558f
C302 source.n131 a_n2094_n2088# 0.019108f
C303 source.n132 a_n2094_n2088# 0.020232f
C304 source.n133 a_n2094_n2088# 0.045163f
C305 source.n134 a_n2094_n2088# 0.045163f
C306 source.n135 a_n2094_n2088# 0.020232f
C307 source.n136 a_n2094_n2088# 0.019108f
C308 source.n137 a_n2094_n2088# 0.035558f
C309 source.n138 a_n2094_n2088# 0.035558f
C310 source.n139 a_n2094_n2088# 0.019108f
C311 source.n140 a_n2094_n2088# 0.020232f
C312 source.n141 a_n2094_n2088# 0.045163f
C313 source.n142 a_n2094_n2088# 0.097771f
C314 source.n143 a_n2094_n2088# 0.020232f
C315 source.n144 a_n2094_n2088# 0.019108f
C316 source.n145 a_n2094_n2088# 0.082191f
C317 source.n146 a_n2094_n2088# 0.054706f
C318 source.n147 a_n2094_n2088# 1.29931f
C319 source.n148 a_n2094_n2088# 0.04998f
C320 source.n149 a_n2094_n2088# 0.035558f
C321 source.n150 a_n2094_n2088# 0.019108f
C322 source.n151 a_n2094_n2088# 0.045163f
C323 source.n152 a_n2094_n2088# 0.020232f
C324 source.n153 a_n2094_n2088# 0.035558f
C325 source.n154 a_n2094_n2088# 0.019108f
C326 source.n155 a_n2094_n2088# 0.045163f
C327 source.n156 a_n2094_n2088# 0.020232f
C328 source.n157 a_n2094_n2088# 0.152165f
C329 source.t4 a_n2094_n2088# 0.07361f
C330 source.n158 a_n2094_n2088# 0.033872f
C331 source.n159 a_n2094_n2088# 0.026678f
C332 source.n160 a_n2094_n2088# 0.019108f
C333 source.n161 a_n2094_n2088# 0.846075f
C334 source.n162 a_n2094_n2088# 0.035558f
C335 source.n163 a_n2094_n2088# 0.019108f
C336 source.n164 a_n2094_n2088# 0.020232f
C337 source.n165 a_n2094_n2088# 0.045163f
C338 source.n166 a_n2094_n2088# 0.045163f
C339 source.n167 a_n2094_n2088# 0.020232f
C340 source.n168 a_n2094_n2088# 0.019108f
C341 source.n169 a_n2094_n2088# 0.035558f
C342 source.n170 a_n2094_n2088# 0.035558f
C343 source.n171 a_n2094_n2088# 0.019108f
C344 source.n172 a_n2094_n2088# 0.020232f
C345 source.n173 a_n2094_n2088# 0.045163f
C346 source.n174 a_n2094_n2088# 0.097771f
C347 source.n175 a_n2094_n2088# 0.020232f
C348 source.n176 a_n2094_n2088# 0.019108f
C349 source.n177 a_n2094_n2088# 0.082191f
C350 source.n178 a_n2094_n2088# 0.054706f
C351 source.n179 a_n2094_n2088# 1.29931f
C352 source.t8 a_n2094_n2088# 0.168595f
C353 source.t22 a_n2094_n2088# 0.168595f
C354 source.n180 a_n2094_n2088# 1.31303f
C355 source.n181 a_n2094_n2088# 0.438033f
C356 source.t16 a_n2094_n2088# 0.168595f
C357 source.t17 a_n2094_n2088# 0.168595f
C358 source.n182 a_n2094_n2088# 1.31303f
C359 source.n183 a_n2094_n2088# 0.438033f
C360 source.t7 a_n2094_n2088# 0.168595f
C361 source.t11 a_n2094_n2088# 0.168595f
C362 source.n184 a_n2094_n2088# 1.31303f
C363 source.n185 a_n2094_n2088# 0.438033f
C364 source.t6 a_n2094_n2088# 0.168595f
C365 source.t0 a_n2094_n2088# 0.168595f
C366 source.n186 a_n2094_n2088# 1.31303f
C367 source.n187 a_n2094_n2088# 0.438033f
C368 source.t13 a_n2094_n2088# 0.168595f
C369 source.t23 a_n2094_n2088# 0.168595f
C370 source.n188 a_n2094_n2088# 1.31303f
C371 source.n189 a_n2094_n2088# 0.438033f
C372 source.n190 a_n2094_n2088# 0.04998f
C373 source.n191 a_n2094_n2088# 0.035558f
C374 source.n192 a_n2094_n2088# 0.019108f
C375 source.n193 a_n2094_n2088# 0.045163f
C376 source.n194 a_n2094_n2088# 0.020232f
C377 source.n195 a_n2094_n2088# 0.035558f
C378 source.n196 a_n2094_n2088# 0.019108f
C379 source.n197 a_n2094_n2088# 0.045163f
C380 source.n198 a_n2094_n2088# 0.020232f
C381 source.n199 a_n2094_n2088# 0.152165f
C382 source.t18 a_n2094_n2088# 0.07361f
C383 source.n200 a_n2094_n2088# 0.033872f
C384 source.n201 a_n2094_n2088# 0.026678f
C385 source.n202 a_n2094_n2088# 0.019108f
C386 source.n203 a_n2094_n2088# 0.846075f
C387 source.n204 a_n2094_n2088# 0.035558f
C388 source.n205 a_n2094_n2088# 0.019108f
C389 source.n206 a_n2094_n2088# 0.020232f
C390 source.n207 a_n2094_n2088# 0.045163f
C391 source.n208 a_n2094_n2088# 0.045163f
C392 source.n209 a_n2094_n2088# 0.020232f
C393 source.n210 a_n2094_n2088# 0.019108f
C394 source.n211 a_n2094_n2088# 0.035558f
C395 source.n212 a_n2094_n2088# 0.035558f
C396 source.n213 a_n2094_n2088# 0.019108f
C397 source.n214 a_n2094_n2088# 0.020232f
C398 source.n215 a_n2094_n2088# 0.045163f
C399 source.n216 a_n2094_n2088# 0.097771f
C400 source.n217 a_n2094_n2088# 0.020232f
C401 source.n218 a_n2094_n2088# 0.019108f
C402 source.n219 a_n2094_n2088# 0.082191f
C403 source.n220 a_n2094_n2088# 0.054706f
C404 source.n221 a_n2094_n2088# 0.13655f
C405 source.n222 a_n2094_n2088# 0.04998f
C406 source.n223 a_n2094_n2088# 0.035558f
C407 source.n224 a_n2094_n2088# 0.019108f
C408 source.n225 a_n2094_n2088# 0.045163f
C409 source.n226 a_n2094_n2088# 0.020232f
C410 source.n227 a_n2094_n2088# 0.035558f
C411 source.n228 a_n2094_n2088# 0.019108f
C412 source.n229 a_n2094_n2088# 0.045163f
C413 source.n230 a_n2094_n2088# 0.020232f
C414 source.n231 a_n2094_n2088# 0.152165f
C415 source.t32 a_n2094_n2088# 0.07361f
C416 source.n232 a_n2094_n2088# 0.033872f
C417 source.n233 a_n2094_n2088# 0.026678f
C418 source.n234 a_n2094_n2088# 0.019108f
C419 source.n235 a_n2094_n2088# 0.846075f
C420 source.n236 a_n2094_n2088# 0.035558f
C421 source.n237 a_n2094_n2088# 0.019108f
C422 source.n238 a_n2094_n2088# 0.020232f
C423 source.n239 a_n2094_n2088# 0.045163f
C424 source.n240 a_n2094_n2088# 0.045163f
C425 source.n241 a_n2094_n2088# 0.020232f
C426 source.n242 a_n2094_n2088# 0.019108f
C427 source.n243 a_n2094_n2088# 0.035558f
C428 source.n244 a_n2094_n2088# 0.035558f
C429 source.n245 a_n2094_n2088# 0.019108f
C430 source.n246 a_n2094_n2088# 0.020232f
C431 source.n247 a_n2094_n2088# 0.045163f
C432 source.n248 a_n2094_n2088# 0.097771f
C433 source.n249 a_n2094_n2088# 0.020232f
C434 source.n250 a_n2094_n2088# 0.019108f
C435 source.n251 a_n2094_n2088# 0.082191f
C436 source.n252 a_n2094_n2088# 0.054706f
C437 source.n253 a_n2094_n2088# 0.13655f
C438 source.t26 a_n2094_n2088# 0.168595f
C439 source.t33 a_n2094_n2088# 0.168595f
C440 source.n254 a_n2094_n2088# 1.31303f
C441 source.n255 a_n2094_n2088# 0.438033f
C442 source.t27 a_n2094_n2088# 0.168595f
C443 source.t43 a_n2094_n2088# 0.168595f
C444 source.n256 a_n2094_n2088# 1.31303f
C445 source.n257 a_n2094_n2088# 0.438033f
C446 source.t24 a_n2094_n2088# 0.168595f
C447 source.t46 a_n2094_n2088# 0.168595f
C448 source.n258 a_n2094_n2088# 1.31303f
C449 source.n259 a_n2094_n2088# 0.438033f
C450 source.t25 a_n2094_n2088# 0.168595f
C451 source.t47 a_n2094_n2088# 0.168595f
C452 source.n260 a_n2094_n2088# 1.31303f
C453 source.n261 a_n2094_n2088# 0.438033f
C454 source.t28 a_n2094_n2088# 0.168595f
C455 source.t34 a_n2094_n2088# 0.168595f
C456 source.n262 a_n2094_n2088# 1.31303f
C457 source.n263 a_n2094_n2088# 0.438033f
C458 source.n264 a_n2094_n2088# 0.04998f
C459 source.n265 a_n2094_n2088# 0.035558f
C460 source.n266 a_n2094_n2088# 0.019108f
C461 source.n267 a_n2094_n2088# 0.045163f
C462 source.n268 a_n2094_n2088# 0.020232f
C463 source.n269 a_n2094_n2088# 0.035558f
C464 source.n270 a_n2094_n2088# 0.019108f
C465 source.n271 a_n2094_n2088# 0.045163f
C466 source.n272 a_n2094_n2088# 0.020232f
C467 source.n273 a_n2094_n2088# 0.152165f
C468 source.t29 a_n2094_n2088# 0.07361f
C469 source.n274 a_n2094_n2088# 0.033872f
C470 source.n275 a_n2094_n2088# 0.026678f
C471 source.n276 a_n2094_n2088# 0.019108f
C472 source.n277 a_n2094_n2088# 0.846075f
C473 source.n278 a_n2094_n2088# 0.035558f
C474 source.n279 a_n2094_n2088# 0.019108f
C475 source.n280 a_n2094_n2088# 0.020232f
C476 source.n281 a_n2094_n2088# 0.045163f
C477 source.n282 a_n2094_n2088# 0.045163f
C478 source.n283 a_n2094_n2088# 0.020232f
C479 source.n284 a_n2094_n2088# 0.019108f
C480 source.n285 a_n2094_n2088# 0.035558f
C481 source.n286 a_n2094_n2088# 0.035558f
C482 source.n287 a_n2094_n2088# 0.019108f
C483 source.n288 a_n2094_n2088# 0.020232f
C484 source.n289 a_n2094_n2088# 0.045163f
C485 source.n290 a_n2094_n2088# 0.097771f
C486 source.n291 a_n2094_n2088# 0.020232f
C487 source.n292 a_n2094_n2088# 0.019108f
C488 source.n293 a_n2094_n2088# 0.082191f
C489 source.n294 a_n2094_n2088# 0.054706f
C490 source.n295 a_n2094_n2088# 0.329359f
C491 source.n296 a_n2094_n2088# 1.45021f
C492 drain_right.t2 a_n2094_n2088# 0.181313f
C493 drain_right.t10 a_n2094_n2088# 0.181313f
C494 drain_right.n0 a_n2094_n2088# 1.51511f
C495 drain_right.t9 a_n2094_n2088# 0.181313f
C496 drain_right.t7 a_n2094_n2088# 0.181313f
C497 drain_right.n1 a_n2094_n2088# 1.51215f
C498 drain_right.n2 a_n2094_n2088# 0.858385f
C499 drain_right.t20 a_n2094_n2088# 0.181313f
C500 drain_right.t3 a_n2094_n2088# 0.181313f
C501 drain_right.n3 a_n2094_n2088# 1.51215f
C502 drain_right.n4 a_n2094_n2088# 0.393124f
C503 drain_right.t6 a_n2094_n2088# 0.181313f
C504 drain_right.t21 a_n2094_n2088# 0.181313f
C505 drain_right.n5 a_n2094_n2088# 1.51511f
C506 drain_right.t0 a_n2094_n2088# 0.181313f
C507 drain_right.t18 a_n2094_n2088# 0.181313f
C508 drain_right.n6 a_n2094_n2088# 1.51215f
C509 drain_right.n7 a_n2094_n2088# 0.858385f
C510 drain_right.t1 a_n2094_n2088# 0.181313f
C511 drain_right.t4 a_n2094_n2088# 0.181313f
C512 drain_right.n8 a_n2094_n2088# 1.51215f
C513 drain_right.n9 a_n2094_n2088# 0.393124f
C514 drain_right.n10 a_n2094_n2088# 1.38361f
C515 drain_right.t14 a_n2094_n2088# 0.181313f
C516 drain_right.t11 a_n2094_n2088# 0.181313f
C517 drain_right.n11 a_n2094_n2088# 1.51511f
C518 drain_right.t16 a_n2094_n2088# 0.181313f
C519 drain_right.t15 a_n2094_n2088# 0.181313f
C520 drain_right.n12 a_n2094_n2088# 1.51216f
C521 drain_right.n13 a_n2094_n2088# 0.858378f
C522 drain_right.t13 a_n2094_n2088# 0.181313f
C523 drain_right.t17 a_n2094_n2088# 0.181313f
C524 drain_right.n14 a_n2094_n2088# 1.51216f
C525 drain_right.n15 a_n2094_n2088# 0.422965f
C526 drain_right.t12 a_n2094_n2088# 0.181313f
C527 drain_right.t22 a_n2094_n2088# 0.181313f
C528 drain_right.n16 a_n2094_n2088# 1.51216f
C529 drain_right.n17 a_n2094_n2088# 0.422965f
C530 drain_right.t23 a_n2094_n2088# 0.181313f
C531 drain_right.t8 a_n2094_n2088# 0.181313f
C532 drain_right.n18 a_n2094_n2088# 1.51216f
C533 drain_right.n19 a_n2094_n2088# 0.422965f
C534 drain_right.t19 a_n2094_n2088# 0.181313f
C535 drain_right.t5 a_n2094_n2088# 0.181313f
C536 drain_right.n20 a_n2094_n2088# 1.51216f
C537 drain_right.n21 a_n2094_n2088# 0.735928f
C538 minus.n0 a_n2094_n2088# 0.051288f
C539 minus.t5 a_n2094_n2088# 0.181117f
C540 minus.t9 a_n2094_n2088# 0.175354f
C541 minus.t8 a_n2094_n2088# 0.175354f
C542 minus.t10 a_n2094_n2088# 0.175354f
C543 minus.n1 a_n2094_n2088# 0.085761f
C544 minus.n2 a_n2094_n2088# 0.051288f
C545 minus.t17 a_n2094_n2088# 0.175354f
C546 minus.t3 a_n2094_n2088# 0.175354f
C547 minus.t6 a_n2094_n2088# 0.175354f
C548 minus.n3 a_n2094_n2088# 0.085761f
C549 minus.n4 a_n2094_n2088# 0.051288f
C550 minus.t12 a_n2094_n2088# 0.175354f
C551 minus.t16 a_n2094_n2088# 0.175354f
C552 minus.t2 a_n2094_n2088# 0.175354f
C553 minus.n5 a_n2094_n2088# 0.085761f
C554 minus.t11 a_n2094_n2088# 0.181117f
C555 minus.n6 a_n2094_n2088# 0.101676f
C556 minus.t7 a_n2094_n2088# 0.175354f
C557 minus.n7 a_n2094_n2088# 0.085761f
C558 minus.n8 a_n2094_n2088# 0.017963f
C559 minus.n9 a_n2094_n2088# 0.119255f
C560 minus.n10 a_n2094_n2088# 0.051288f
C561 minus.n11 a_n2094_n2088# 0.017963f
C562 minus.n12 a_n2094_n2088# 0.085761f
C563 minus.n13 a_n2094_n2088# 0.017963f
C564 minus.n14 a_n2094_n2088# 0.085761f
C565 minus.n15 a_n2094_n2088# 0.017963f
C566 minus.n16 a_n2094_n2088# 0.051288f
C567 minus.n17 a_n2094_n2088# 0.051288f
C568 minus.n18 a_n2094_n2088# 0.017963f
C569 minus.n19 a_n2094_n2088# 0.085761f
C570 minus.n20 a_n2094_n2088# 0.017963f
C571 minus.n21 a_n2094_n2088# 0.085761f
C572 minus.n22 a_n2094_n2088# 0.017963f
C573 minus.n23 a_n2094_n2088# 0.051288f
C574 minus.n24 a_n2094_n2088# 0.051288f
C575 minus.n25 a_n2094_n2088# 0.017963f
C576 minus.n26 a_n2094_n2088# 0.085761f
C577 minus.n27 a_n2094_n2088# 0.017963f
C578 minus.n28 a_n2094_n2088# 0.085761f
C579 minus.n29 a_n2094_n2088# 0.101597f
C580 minus.n30 a_n2094_n2088# 1.52479f
C581 minus.n31 a_n2094_n2088# 0.051288f
C582 minus.t13 a_n2094_n2088# 0.175354f
C583 minus.t19 a_n2094_n2088# 0.175354f
C584 minus.t0 a_n2094_n2088# 0.175354f
C585 minus.n32 a_n2094_n2088# 0.085761f
C586 minus.n33 a_n2094_n2088# 0.051288f
C587 minus.t22 a_n2094_n2088# 0.175354f
C588 minus.t1 a_n2094_n2088# 0.175354f
C589 minus.t23 a_n2094_n2088# 0.175354f
C590 minus.n34 a_n2094_n2088# 0.085761f
C591 minus.n35 a_n2094_n2088# 0.051288f
C592 minus.t4 a_n2094_n2088# 0.175354f
C593 minus.t20 a_n2094_n2088# 0.175354f
C594 minus.t14 a_n2094_n2088# 0.175354f
C595 minus.n36 a_n2094_n2088# 0.085761f
C596 minus.t15 a_n2094_n2088# 0.181117f
C597 minus.n37 a_n2094_n2088# 0.101676f
C598 minus.t21 a_n2094_n2088# 0.175354f
C599 minus.n38 a_n2094_n2088# 0.085761f
C600 minus.n39 a_n2094_n2088# 0.017963f
C601 minus.n40 a_n2094_n2088# 0.119255f
C602 minus.n41 a_n2094_n2088# 0.051288f
C603 minus.n42 a_n2094_n2088# 0.017963f
C604 minus.n43 a_n2094_n2088# 0.085761f
C605 minus.n44 a_n2094_n2088# 0.017963f
C606 minus.n45 a_n2094_n2088# 0.085761f
C607 minus.n46 a_n2094_n2088# 0.017963f
C608 minus.n47 a_n2094_n2088# 0.051288f
C609 minus.n48 a_n2094_n2088# 0.051288f
C610 minus.n49 a_n2094_n2088# 0.017963f
C611 minus.n50 a_n2094_n2088# 0.085761f
C612 minus.n51 a_n2094_n2088# 0.017963f
C613 minus.n52 a_n2094_n2088# 0.085761f
C614 minus.n53 a_n2094_n2088# 0.017963f
C615 minus.n54 a_n2094_n2088# 0.051288f
C616 minus.n55 a_n2094_n2088# 0.051288f
C617 minus.n56 a_n2094_n2088# 0.017963f
C618 minus.n57 a_n2094_n2088# 0.085761f
C619 minus.n58 a_n2094_n2088# 0.017963f
C620 minus.n59 a_n2094_n2088# 0.085761f
C621 minus.t18 a_n2094_n2088# 0.181117f
C622 minus.n60 a_n2094_n2088# 0.101597f
C623 minus.n61 a_n2094_n2088# 0.333994f
C624 minus.n62 a_n2094_n2088# 1.87178f
.ends

