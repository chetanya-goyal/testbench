* NGSPICE file created from diffpair243.ext - technology: sky130A

.subckt diffpair243 minus drain_right drain_left source plus
X0 source plus drain_left a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X1 a_n1366_n2088# a_n1366_n2088# a_n1366_n2088# a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=22.8 ps=103.6 w=6 l=0.15
X2 a_n1366_n2088# a_n1366_n2088# a_n1366_n2088# a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X3 drain_left plus source a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X4 a_n1366_n2088# a_n1366_n2088# a_n1366_n2088# a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X5 drain_right minus source a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X6 source plus drain_left a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X7 source minus drain_right a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X8 a_n1366_n2088# a_n1366_n2088# a_n1366_n2088# a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X9 source minus drain_right a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X10 drain_right minus source a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X11 drain_right minus source a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X12 source minus drain_right a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X13 source plus drain_left a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X14 drain_right minus source a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X15 source minus drain_right a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=2.85 pd=12.95 as=1.5 ps=6.5 w=6 l=0.15
X16 drain_left plus source a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=2.85 ps=12.95 w=6 l=0.15
X17 source plus drain_left a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X18 drain_left plus source a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
X19 drain_left plus source a_n1366_n2088# sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.15
.ends

