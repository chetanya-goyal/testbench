* NGSPICE file created from diffpair563.ext - technology: sky130A

.subckt diffpair563 minus drain_right drain_left source plus
X0 a_n1366_n4888# a_n1366_n4888# a_n1366_n4888# a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=76 ps=327.6 w=20 l=0.15
X1 drain_right.t7 minus.t0 source.t6 a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X2 source.t5 minus.t1 drain_right.t6 a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X3 drain_left.t7 plus.t0 source.t15 a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X4 a_n1366_n4888# a_n1366_n4888# a_n1366_n4888# a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X5 source.t10 minus.t2 drain_right.t5 a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X6 a_n1366_n4888# a_n1366_n4888# a_n1366_n4888# a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X7 source.t2 plus.t1 drain_left.t6 a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X8 drain_right.t4 minus.t3 source.t7 a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X9 source.t9 minus.t4 drain_right.t3 a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X10 a_n1366_n4888# a_n1366_n4888# a_n1366_n4888# a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=0 ps=0 w=20 l=0.15
X11 drain_left.t5 plus.t2 source.t1 a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X12 source.t4 plus.t3 drain_left.t4 a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=9.5 pd=40.95 as=5 ps=20.5 w=20 l=0.15
X13 drain_right.t2 minus.t5 source.t8 a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X14 drain_right.t1 minus.t6 source.t11 a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X15 drain_left.t3 plus.t4 source.t0 a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=9.5 ps=40.95 w=20 l=0.15
X16 source.t14 plus.t5 drain_left.t2 a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X17 source.t3 plus.t6 drain_left.t1 a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X18 drain_left.t0 plus.t7 source.t13 a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
X19 source.t12 minus.t7 drain_right.t0 a_n1366_n4888# sky130_fd_pr__nfet_01v8 ad=5 pd=20.5 as=5 ps=20.5 w=20 l=0.15
R0 minus.n5 minus.t4 3491.58
R1 minus.n1 minus.t3 3491.58
R2 minus.n12 minus.t0 3491.58
R3 minus.n8 minus.t1 3491.58
R4 minus.n4 minus.t5 3422.2
R5 minus.n2 minus.t2 3422.2
R6 minus.n11 minus.t7 3422.2
R7 minus.n9 minus.t6 3422.2
R8 minus.n1 minus.n0 161.489
R9 minus.n8 minus.n7 161.489
R10 minus.n6 minus.n5 161.3
R11 minus.n3 minus.n0 161.3
R12 minus.n13 minus.n12 161.3
R13 minus.n10 minus.n7 161.3
R14 minus.n4 minus.n3 47.4702
R15 minus.n3 minus.n2 47.4702
R16 minus.n10 minus.n9 47.4702
R17 minus.n11 minus.n10 47.4702
R18 minus.n14 minus.n6 40.4361
R19 minus.n5 minus.n4 25.5611
R20 minus.n2 minus.n1 25.5611
R21 minus.n9 minus.n8 25.5611
R22 minus.n12 minus.n11 25.5611
R23 minus.n14 minus.n13 6.58005
R24 minus.n6 minus.n0 0.189894
R25 minus.n13 minus.n7 0.189894
R26 minus minus.n14 0.188
R27 source.n0 source.t0 44.6397
R28 source.n3 source.t4 44.6396
R29 source.n4 source.t7 44.6396
R30 source.n7 source.t9 44.6396
R31 source.n15 source.t6 44.6395
R32 source.n12 source.t5 44.6395
R33 source.n11 source.t1 44.6395
R34 source.n8 source.t2 44.6395
R35 source.n2 source.n1 43.1397
R36 source.n6 source.n5 43.1397
R37 source.n14 source.n13 43.1396
R38 source.n10 source.n9 43.1396
R39 source.n8 source.n7 27.9087
R40 source.n16 source.n0 22.3656
R41 source.n16 source.n15 5.5436
R42 source.n13 source.t11 1.5005
R43 source.n13 source.t12 1.5005
R44 source.n9 source.t15 1.5005
R45 source.n9 source.t3 1.5005
R46 source.n1 source.t13 1.5005
R47 source.n1 source.t14 1.5005
R48 source.n5 source.t8 1.5005
R49 source.n5 source.t10 1.5005
R50 source.n7 source.n6 0.560845
R51 source.n6 source.n4 0.560845
R52 source.n3 source.n2 0.560845
R53 source.n2 source.n0 0.560845
R54 source.n10 source.n8 0.560845
R55 source.n11 source.n10 0.560845
R56 source.n14 source.n12 0.560845
R57 source.n15 source.n14 0.560845
R58 source.n4 source.n3 0.470328
R59 source.n12 source.n11 0.470328
R60 source source.n16 0.188
R61 drain_right.n5 drain_right.n3 60.3788
R62 drain_right.n2 drain_right.n1 60.0432
R63 drain_right.n2 drain_right.n0 60.0432
R64 drain_right.n5 drain_right.n4 59.8185
R65 drain_right drain_right.n2 34.8357
R66 drain_right drain_right.n5 6.21356
R67 drain_right.n1 drain_right.t0 1.5005
R68 drain_right.n1 drain_right.t7 1.5005
R69 drain_right.n0 drain_right.t6 1.5005
R70 drain_right.n0 drain_right.t1 1.5005
R71 drain_right.n3 drain_right.t5 1.5005
R72 drain_right.n3 drain_right.t4 1.5005
R73 drain_right.n4 drain_right.t3 1.5005
R74 drain_right.n4 drain_right.t2 1.5005
R75 plus.n1 plus.t3 3491.58
R76 plus.n5 plus.t4 3491.58
R77 plus.n8 plus.t2 3491.58
R78 plus.n12 plus.t1 3491.58
R79 plus.n2 plus.t7 3422.2
R80 plus.n4 plus.t5 3422.2
R81 plus.n9 plus.t6 3422.2
R82 plus.n11 plus.t0 3422.2
R83 plus.n1 plus.n0 161.489
R84 plus.n8 plus.n7 161.489
R85 plus.n3 plus.n0 161.3
R86 plus.n6 plus.n5 161.3
R87 plus.n10 plus.n7 161.3
R88 plus.n13 plus.n12 161.3
R89 plus.n3 plus.n2 47.4702
R90 plus.n4 plus.n3 47.4702
R91 plus.n11 plus.n10 47.4702
R92 plus.n10 plus.n9 47.4702
R93 plus plus.n13 31.2869
R94 plus.n2 plus.n1 25.5611
R95 plus.n5 plus.n4 25.5611
R96 plus.n12 plus.n11 25.5611
R97 plus.n9 plus.n8 25.5611
R98 plus plus.n6 15.2543
R99 plus.n6 plus.n0 0.189894
R100 plus.n13 plus.n7 0.189894
R101 drain_left.n5 drain_left.n3 60.3788
R102 drain_left.n2 drain_left.n1 60.0432
R103 drain_left.n2 drain_left.n0 60.0432
R104 drain_left.n5 drain_left.n4 59.8185
R105 drain_left drain_left.n2 35.3889
R106 drain_left drain_left.n5 6.21356
R107 drain_left.n1 drain_left.t1 1.5005
R108 drain_left.n1 drain_left.t5 1.5005
R109 drain_left.n0 drain_left.t6 1.5005
R110 drain_left.n0 drain_left.t7 1.5005
R111 drain_left.n4 drain_left.t2 1.5005
R112 drain_left.n4 drain_left.t3 1.5005
R113 drain_left.n3 drain_left.t4 1.5005
R114 drain_left.n3 drain_left.t0 1.5005
C0 drain_left minus 0.170499f
C1 source plus 2.46827f
C2 source minus 2.45423f
C3 minus plus 6.31655f
C4 drain_right drain_left 0.640281f
C5 drain_right source 26.9295f
C6 drain_right plus 0.282599f
C7 drain_right minus 3.39574f
C8 source drain_left 26.930199f
C9 drain_left plus 3.52513f
C10 drain_right a_n1366_n4888# 6.84971f
C11 drain_left a_n1366_n4888# 7.04335f
C12 source a_n1366_n4888# 12.931394f
C13 minus a_n1366_n4888# 5.533225f
C14 plus a_n1366_n4888# 8.396939f
C15 drain_left.t6 a_n1366_n4888# 0.674884f
C16 drain_left.t7 a_n1366_n4888# 0.674884f
C17 drain_left.n0 a_n1366_n4888# 4.53229f
C18 drain_left.t1 a_n1366_n4888# 0.674884f
C19 drain_left.t5 a_n1366_n4888# 0.674884f
C20 drain_left.n1 a_n1366_n4888# 4.53229f
C21 drain_left.n2 a_n1366_n4888# 2.4394f
C22 drain_left.t4 a_n1366_n4888# 0.674884f
C23 drain_left.t0 a_n1366_n4888# 0.674884f
C24 drain_left.n3 a_n1366_n4888# 4.53433f
C25 drain_left.t2 a_n1366_n4888# 0.674884f
C26 drain_left.t3 a_n1366_n4888# 0.674884f
C27 drain_left.n4 a_n1366_n4888# 4.53107f
C28 drain_left.n5 a_n1366_n4888# 0.92266f
C29 plus.n0 a_n1366_n4888# 0.14635f
C30 plus.t5 a_n1366_n4888# 0.522133f
C31 plus.t7 a_n1366_n4888# 0.522133f
C32 plus.t3 a_n1366_n4888# 0.52627f
C33 plus.n1 a_n1366_n4888# 0.230423f
C34 plus.n2 a_n1366_n4888# 0.203484f
C35 plus.n3 a_n1366_n4888# 0.026214f
C36 plus.n4 a_n1366_n4888# 0.203484f
C37 plus.t4 a_n1366_n4888# 0.52627f
C38 plus.n5 a_n1366_n4888# 0.230323f
C39 plus.n6 a_n1366_n4888# 0.949674f
C40 plus.n7 a_n1366_n4888# 0.14635f
C41 plus.t1 a_n1366_n4888# 0.52627f
C42 plus.t0 a_n1366_n4888# 0.522133f
C43 plus.t6 a_n1366_n4888# 0.522133f
C44 plus.t2 a_n1366_n4888# 0.52627f
C45 plus.n8 a_n1366_n4888# 0.230423f
C46 plus.n9 a_n1366_n4888# 0.203484f
C47 plus.n10 a_n1366_n4888# 0.026214f
C48 plus.n11 a_n1366_n4888# 0.203484f
C49 plus.n12 a_n1366_n4888# 0.230323f
C50 plus.n13 a_n1366_n4888# 2.0373f
C51 drain_right.t6 a_n1366_n4888# 0.675112f
C52 drain_right.t1 a_n1366_n4888# 0.675112f
C53 drain_right.n0 a_n1366_n4888# 4.53382f
C54 drain_right.t0 a_n1366_n4888# 0.675112f
C55 drain_right.t7 a_n1366_n4888# 0.675112f
C56 drain_right.n1 a_n1366_n4888# 4.53382f
C57 drain_right.n2 a_n1366_n4888# 2.3811f
C58 drain_right.t5 a_n1366_n4888# 0.675112f
C59 drain_right.t4 a_n1366_n4888# 0.675112f
C60 drain_right.n3 a_n1366_n4888# 4.53586f
C61 drain_right.t3 a_n1366_n4888# 0.675112f
C62 drain_right.t2 a_n1366_n4888# 0.675112f
C63 drain_right.n4 a_n1366_n4888# 4.532609f
C64 drain_right.n5 a_n1366_n4888# 0.922972f
C65 source.t0 a_n1366_n4888# 3.94438f
C66 source.n0 a_n1366_n4888# 1.60143f
C67 source.t13 a_n1366_n4888# 0.485004f
C68 source.t14 a_n1366_n4888# 0.485004f
C69 source.n1 a_n1366_n4888# 3.19166f
C70 source.n2 a_n1366_n4888# 0.281117f
C71 source.t4 a_n1366_n4888# 3.94439f
C72 source.n3 a_n1366_n4888# 0.395488f
C73 source.t7 a_n1366_n4888# 3.94439f
C74 source.n4 a_n1366_n4888# 0.395488f
C75 source.t8 a_n1366_n4888# 0.485004f
C76 source.t10 a_n1366_n4888# 0.485004f
C77 source.n5 a_n1366_n4888# 3.19166f
C78 source.n6 a_n1366_n4888# 0.281117f
C79 source.t9 a_n1366_n4888# 3.94439f
C80 source.n7 a_n1366_n4888# 1.96083f
C81 source.t2 a_n1366_n4888# 3.94437f
C82 source.n8 a_n1366_n4888# 1.96085f
C83 source.t15 a_n1366_n4888# 0.485004f
C84 source.t3 a_n1366_n4888# 0.485004f
C85 source.n9 a_n1366_n4888# 3.19166f
C86 source.n10 a_n1366_n4888# 0.281111f
C87 source.t1 a_n1366_n4888# 3.94437f
C88 source.n11 a_n1366_n4888# 0.395508f
C89 source.t5 a_n1366_n4888# 3.94437f
C90 source.n12 a_n1366_n4888# 0.395508f
C91 source.t11 a_n1366_n4888# 0.485004f
C92 source.t12 a_n1366_n4888# 0.485004f
C93 source.n13 a_n1366_n4888# 3.19166f
C94 source.n14 a_n1366_n4888# 0.281111f
C95 source.t6 a_n1366_n4888# 3.94437f
C96 source.n15 a_n1366_n4888# 0.51074f
C97 source.n16 a_n1366_n4888# 1.82392f
C98 minus.n0 a_n1366_n4888# 0.1437f
C99 minus.t4 a_n1366_n4888# 0.516742f
C100 minus.t5 a_n1366_n4888# 0.512679f
C101 minus.t2 a_n1366_n4888# 0.512679f
C102 minus.t3 a_n1366_n4888# 0.516742f
C103 minus.n1 a_n1366_n4888# 0.226251f
C104 minus.n2 a_n1366_n4888# 0.1998f
C105 minus.n3 a_n1366_n4888# 0.02574f
C106 minus.n4 a_n1366_n4888# 0.1998f
C107 minus.n5 a_n1366_n4888# 0.226153f
C108 minus.n6 a_n1366_n4888# 2.54342f
C109 minus.n7 a_n1366_n4888# 0.1437f
C110 minus.t7 a_n1366_n4888# 0.512679f
C111 minus.t6 a_n1366_n4888# 0.512679f
C112 minus.t1 a_n1366_n4888# 0.516742f
C113 minus.n8 a_n1366_n4888# 0.226251f
C114 minus.n9 a_n1366_n4888# 0.1998f
C115 minus.n10 a_n1366_n4888# 0.02574f
C116 minus.n11 a_n1366_n4888# 0.1998f
C117 minus.t0 a_n1366_n4888# 0.516742f
C118 minus.n12 a_n1366_n4888# 0.226153f
C119 minus.n13 a_n1366_n4888# 0.408084f
C120 minus.n14 a_n1366_n4888# 3.04808f
.ends

