* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t18 minus.t0 drain_right.t1 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X1 a_n2072_n1288# a_n2072_n1288# a_n2072_n1288# a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.8
X2 source.t17 minus.t1 drain_right.t6 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X3 source.t19 plus.t0 drain_left.t9 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X4 source.t3 plus.t1 drain_left.t8 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X5 a_n2072_n1288# a_n2072_n1288# a_n2072_n1288# a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X6 a_n2072_n1288# a_n2072_n1288# a_n2072_n1288# a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X7 drain_right.t7 minus.t2 source.t16 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X8 source.t15 minus.t3 drain_right.t3 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X9 drain_right.t2 minus.t4 source.t14 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X10 drain_right.t4 minus.t5 source.t13 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X11 drain_left.t7 plus.t2 source.t2 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X12 source.t12 minus.t6 drain_right.t0 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X13 drain_right.t8 minus.t7 source.t11 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X14 a_n2072_n1288# a_n2072_n1288# a_n2072_n1288# a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.8
X15 source.t8 plus.t3 drain_left.t6 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X16 drain_right.t9 minus.t8 source.t10 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X17 drain_left.t5 plus.t4 source.t4 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X18 drain_right.t5 minus.t9 source.t9 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X19 drain_left.t4 plus.t5 source.t7 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X20 source.t5 plus.t6 drain_left.t3 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
X21 drain_left.t2 plus.t7 source.t6 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.8
X22 drain_left.t1 plus.t8 source.t0 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.8
X23 drain_left.t0 plus.t9 source.t1 a_n2072_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.8
R0 minus.n9 minus.n8 161.3
R1 minus.n7 minus.n0 161.3
R2 minus.n19 minus.n18 161.3
R3 minus.n17 minus.n10 161.3
R4 minus.n3 minus.t4 132.55
R5 minus.n13 minus.t8 132.55
R6 minus.n2 minus.t3 109.355
R7 minus.n1 minus.t2 109.355
R8 minus.n6 minus.t6 109.355
R9 minus.n8 minus.t7 109.355
R10 minus.n12 minus.t0 109.355
R11 minus.n11 minus.t9 109.355
R12 minus.n16 minus.t1 109.355
R13 minus.n18 minus.t5 109.355
R14 minus.n6 minus.n5 80.6037
R15 minus.n4 minus.n1 80.6037
R16 minus.n16 minus.n15 80.6037
R17 minus.n14 minus.n11 80.6037
R18 minus.n2 minus.n1 48.2005
R19 minus.n6 minus.n1 48.2005
R20 minus.n12 minus.n11 48.2005
R21 minus.n16 minus.n11 48.2005
R22 minus.n7 minus.n6 32.1338
R23 minus.n17 minus.n16 32.1338
R24 minus.n4 minus.n3 31.8629
R25 minus.n14 minus.n13 31.8629
R26 minus.n20 minus.n9 29.5706
R27 minus.n3 minus.n2 16.2333
R28 minus.n13 minus.n12 16.2333
R29 minus.n8 minus.n7 16.0672
R30 minus.n18 minus.n17 16.0672
R31 minus.n20 minus.n19 6.67664
R32 minus.n5 minus.n4 0.380177
R33 minus.n15 minus.n14 0.380177
R34 minus.n5 minus.n0 0.285035
R35 minus.n15 minus.n10 0.285035
R36 minus.n9 minus.n0 0.189894
R37 minus.n19 minus.n10 0.189894
R38 minus minus.n20 0.188
R39 drain_right.n2 drain_right.n0 289.615
R40 drain_right.n16 drain_right.n14 289.615
R41 drain_right.n3 drain_right.n2 185
R42 drain_right.n17 drain_right.n16 185
R43 drain_right.t9 drain_right.n1 167.117
R44 drain_right.t8 drain_right.n15 167.117
R45 drain_right.n13 drain_right.n11 101.769
R46 drain_right.n10 drain_right.n9 101.471
R47 drain_right.n13 drain_right.n12 100.796
R48 drain_right.n8 drain_right.n7 100.796
R49 drain_right.n2 drain_right.t9 52.3082
R50 drain_right.n16 drain_right.t8 52.3082
R51 drain_right.n8 drain_right.n6 49.0625
R52 drain_right.n21 drain_right.n20 48.0884
R53 drain_right drain_right.n10 23.3782
R54 drain_right.n9 drain_right.t6 9.9005
R55 drain_right.n9 drain_right.t4 9.9005
R56 drain_right.n7 drain_right.t1 9.9005
R57 drain_right.n7 drain_right.t5 9.9005
R58 drain_right.n11 drain_right.t3 9.9005
R59 drain_right.n11 drain_right.t2 9.9005
R60 drain_right.n12 drain_right.t0 9.9005
R61 drain_right.n12 drain_right.t7 9.9005
R62 drain_right.n3 drain_right.n1 9.71174
R63 drain_right.n17 drain_right.n15 9.71174
R64 drain_right.n6 drain_right.n5 9.45567
R65 drain_right.n20 drain_right.n19 9.45567
R66 drain_right.n5 drain_right.n4 9.3005
R67 drain_right.n19 drain_right.n18 9.3005
R68 drain_right.n6 drain_right.n0 8.14595
R69 drain_right.n20 drain_right.n14 8.14595
R70 drain_right.n4 drain_right.n3 7.3702
R71 drain_right.n18 drain_right.n17 7.3702
R72 drain_right drain_right.n21 6.14028
R73 drain_right.n4 drain_right.n0 5.81868
R74 drain_right.n18 drain_right.n14 5.81868
R75 drain_right.n5 drain_right.n1 3.44771
R76 drain_right.n19 drain_right.n15 3.44771
R77 drain_right.n21 drain_right.n13 0.974638
R78 drain_right.n10 drain_right.n8 0.188688
R79 source.n42 source.n40 289.615
R80 source.n30 source.n28 289.615
R81 source.n2 source.n0 289.615
R82 source.n14 source.n12 289.615
R83 source.n43 source.n42 185
R84 source.n31 source.n30 185
R85 source.n3 source.n2 185
R86 source.n15 source.n14 185
R87 source.t13 source.n41 167.117
R88 source.t6 source.n29 167.117
R89 source.t7 source.n1 167.117
R90 source.t14 source.n13 167.117
R91 source.n9 source.n8 84.1169
R92 source.n11 source.n10 84.1169
R93 source.n21 source.n20 84.1169
R94 source.n23 source.n22 84.1169
R95 source.n39 source.n38 84.1168
R96 source.n37 source.n36 84.1168
R97 source.n27 source.n26 84.1168
R98 source.n25 source.n24 84.1168
R99 source.n42 source.t13 52.3082
R100 source.n30 source.t6 52.3082
R101 source.n2 source.t7 52.3082
R102 source.n14 source.t14 52.3082
R103 source.n47 source.n46 31.4096
R104 source.n35 source.n34 31.4096
R105 source.n7 source.n6 31.4096
R106 source.n19 source.n18 31.4096
R107 source.n25 source.n23 15.6602
R108 source.n38 source.t9 9.9005
R109 source.n38 source.t17 9.9005
R110 source.n36 source.t10 9.9005
R111 source.n36 source.t18 9.9005
R112 source.n26 source.t1 9.9005
R113 source.n26 source.t19 9.9005
R114 source.n24 source.t2 9.9005
R115 source.n24 source.t3 9.9005
R116 source.n8 source.t4 9.9005
R117 source.n8 source.t8 9.9005
R118 source.n10 source.t0 9.9005
R119 source.n10 source.t5 9.9005
R120 source.n20 source.t16 9.9005
R121 source.n20 source.t15 9.9005
R122 source.n22 source.t11 9.9005
R123 source.n22 source.t12 9.9005
R124 source.n43 source.n41 9.71174
R125 source.n31 source.n29 9.71174
R126 source.n3 source.n1 9.71174
R127 source.n15 source.n13 9.71174
R128 source.n46 source.n45 9.45567
R129 source.n34 source.n33 9.45567
R130 source.n6 source.n5 9.45567
R131 source.n18 source.n17 9.45567
R132 source.n45 source.n44 9.3005
R133 source.n33 source.n32 9.3005
R134 source.n5 source.n4 9.3005
R135 source.n17 source.n16 9.3005
R136 source.n48 source.n7 8.93611
R137 source.n46 source.n40 8.14595
R138 source.n34 source.n28 8.14595
R139 source.n6 source.n0 8.14595
R140 source.n18 source.n12 8.14595
R141 source.n44 source.n43 7.3702
R142 source.n32 source.n31 7.3702
R143 source.n4 source.n3 7.3702
R144 source.n16 source.n15 7.3702
R145 source.n44 source.n40 5.81868
R146 source.n32 source.n28 5.81868
R147 source.n4 source.n0 5.81868
R148 source.n16 source.n12 5.81868
R149 source.n48 source.n47 5.7505
R150 source.n45 source.n41 3.44771
R151 source.n33 source.n29 3.44771
R152 source.n5 source.n1 3.44771
R153 source.n17 source.n13 3.44771
R154 source.n23 source.n21 0.974638
R155 source.n21 source.n19 0.974638
R156 source.n11 source.n9 0.974638
R157 source.n9 source.n7 0.974638
R158 source.n27 source.n25 0.974638
R159 source.n35 source.n27 0.974638
R160 source.n39 source.n37 0.974638
R161 source.n47 source.n39 0.974638
R162 source.n19 source.n11 0.957397
R163 source.n37 source.n35 0.957397
R164 source source.n48 0.188
R165 plus.n7 plus.n0 161.3
R166 plus.n9 plus.n8 161.3
R167 plus.n17 plus.n10 161.3
R168 plus.n19 plus.n18 161.3
R169 plus.n3 plus.t8 132.55
R170 plus.n13 plus.t7 132.55
R171 plus.n8 plus.t5 109.355
R172 plus.n6 plus.t3 109.355
R173 plus.n5 plus.t4 109.355
R174 plus.n4 plus.t6 109.355
R175 plus.n18 plus.t2 109.355
R176 plus.n16 plus.t1 109.355
R177 plus.n15 plus.t9 109.355
R178 plus.n14 plus.t0 109.355
R179 plus.n5 plus.n2 80.6037
R180 plus.n6 plus.n1 80.6037
R181 plus.n15 plus.n12 80.6037
R182 plus.n16 plus.n11 80.6037
R183 plus.n6 plus.n5 48.2005
R184 plus.n5 plus.n4 48.2005
R185 plus.n16 plus.n15 48.2005
R186 plus.n15 plus.n14 48.2005
R187 plus.n7 plus.n6 32.1338
R188 plus.n17 plus.n16 32.1338
R189 plus.n3 plus.n2 31.8629
R190 plus.n13 plus.n12 31.8629
R191 plus plus.n19 27.2396
R192 plus.n4 plus.n3 16.2333
R193 plus.n14 plus.n13 16.2333
R194 plus.n8 plus.n7 16.0672
R195 plus.n18 plus.n17 16.0672
R196 plus plus.n9 8.5327
R197 plus.n2 plus.n1 0.380177
R198 plus.n12 plus.n11 0.380177
R199 plus.n1 plus.n0 0.285035
R200 plus.n11 plus.n10 0.285035
R201 plus.n9 plus.n0 0.189894
R202 plus.n19 plus.n10 0.189894
R203 drain_left.n2 drain_left.n0 289.615
R204 drain_left.n13 drain_left.n11 289.615
R205 drain_left.n3 drain_left.n2 185
R206 drain_left.n14 drain_left.n13 185
R207 drain_left.t7 drain_left.n1 167.117
R208 drain_left.t1 drain_left.n12 167.117
R209 drain_left.n10 drain_left.n9 101.471
R210 drain_left.n21 drain_left.n20 100.796
R211 drain_left.n19 drain_left.n18 100.796
R212 drain_left.n8 drain_left.n7 100.796
R213 drain_left.n2 drain_left.t7 52.3082
R214 drain_left.n13 drain_left.t1 52.3082
R215 drain_left.n8 drain_left.n6 49.0625
R216 drain_left.n19 drain_left.n17 49.0625
R217 drain_left drain_left.n10 23.9314
R218 drain_left.n9 drain_left.t9 9.9005
R219 drain_left.n9 drain_left.t2 9.9005
R220 drain_left.n7 drain_left.t8 9.9005
R221 drain_left.n7 drain_left.t0 9.9005
R222 drain_left.n20 drain_left.t6 9.9005
R223 drain_left.n20 drain_left.t4 9.9005
R224 drain_left.n18 drain_left.t3 9.9005
R225 drain_left.n18 drain_left.t5 9.9005
R226 drain_left.n3 drain_left.n1 9.71174
R227 drain_left.n14 drain_left.n12 9.71174
R228 drain_left.n6 drain_left.n5 9.45567
R229 drain_left.n17 drain_left.n16 9.45567
R230 drain_left.n5 drain_left.n4 9.3005
R231 drain_left.n16 drain_left.n15 9.3005
R232 drain_left.n6 drain_left.n0 8.14595
R233 drain_left.n17 drain_left.n11 8.14595
R234 drain_left.n4 drain_left.n3 7.3702
R235 drain_left.n15 drain_left.n14 7.3702
R236 drain_left drain_left.n21 6.62735
R237 drain_left.n4 drain_left.n0 5.81868
R238 drain_left.n15 drain_left.n11 5.81868
R239 drain_left.n5 drain_left.n1 3.44771
R240 drain_left.n16 drain_left.n12 3.44771
R241 drain_left.n21 drain_left.n19 0.974638
R242 drain_left.n10 drain_left.n8 0.188688
C0 source drain_left 4.50249f
C1 plus drain_right 0.365907f
C2 minus drain_left 0.178807f
C3 minus source 1.98352f
C4 plus drain_left 1.77003f
C5 plus source 1.99756f
C6 drain_right drain_left 1.03091f
C7 drain_right source 4.50291f
C8 plus minus 3.88023f
C9 drain_right minus 1.56775f
C10 drain_right a_n2072_n1288# 3.884497f
C11 drain_left a_n2072_n1288# 4.155849f
C12 source a_n2072_n1288# 2.671324f
C13 minus a_n2072_n1288# 7.288625f
C14 plus a_n2072_n1288# 7.807425f
C15 drain_left.n0 a_n2072_n1288# 0.025704f
C16 drain_left.n1 a_n2072_n1288# 0.056872f
C17 drain_left.t7 a_n2072_n1288# 0.04268f
C18 drain_left.n2 a_n2072_n1288# 0.04451f
C19 drain_left.n3 a_n2072_n1288# 0.014348f
C20 drain_left.n4 a_n2072_n1288# 0.009463f
C21 drain_left.n5 a_n2072_n1288# 0.12536f
C22 drain_left.n6 a_n2072_n1288# 0.042104f
C23 drain_left.t8 a_n2072_n1288# 0.027833f
C24 drain_left.t0 a_n2072_n1288# 0.027833f
C25 drain_left.n7 a_n2072_n1288# 0.174852f
C26 drain_left.n8 a_n2072_n1288# 0.28979f
C27 drain_left.t9 a_n2072_n1288# 0.027833f
C28 drain_left.t2 a_n2072_n1288# 0.027833f
C29 drain_left.n9 a_n2072_n1288# 0.176423f
C30 drain_left.n10 a_n2072_n1288# 0.795828f
C31 drain_left.n11 a_n2072_n1288# 0.025704f
C32 drain_left.n12 a_n2072_n1288# 0.056872f
C33 drain_left.t1 a_n2072_n1288# 0.04268f
C34 drain_left.n13 a_n2072_n1288# 0.04451f
C35 drain_left.n14 a_n2072_n1288# 0.014348f
C36 drain_left.n15 a_n2072_n1288# 0.009463f
C37 drain_left.n16 a_n2072_n1288# 0.12536f
C38 drain_left.n17 a_n2072_n1288# 0.042104f
C39 drain_left.t3 a_n2072_n1288# 0.027833f
C40 drain_left.t5 a_n2072_n1288# 0.027833f
C41 drain_left.n18 a_n2072_n1288# 0.174853f
C42 drain_left.n19 a_n2072_n1288# 0.332218f
C43 drain_left.t6 a_n2072_n1288# 0.027833f
C44 drain_left.t4 a_n2072_n1288# 0.027833f
C45 drain_left.n20 a_n2072_n1288# 0.174853f
C46 drain_left.n21 a_n2072_n1288# 0.403253f
C47 plus.n0 a_n2072_n1288# 0.031315f
C48 plus.t5 a_n2072_n1288# 0.116278f
C49 plus.t3 a_n2072_n1288# 0.116278f
C50 plus.n1 a_n2072_n1288# 0.039089f
C51 plus.t4 a_n2072_n1288# 0.116278f
C52 plus.n2 a_n2072_n1288# 0.144015f
C53 plus.t6 a_n2072_n1288# 0.116278f
C54 plus.t8 a_n2072_n1288# 0.130356f
C55 plus.n3 a_n2072_n1288# 0.069028f
C56 plus.n4 a_n2072_n1288# 0.085322f
C57 plus.n5 a_n2072_n1288# 0.08589f
C58 plus.n6 a_n2072_n1288# 0.084298f
C59 plus.n7 a_n2072_n1288# 0.005325f
C60 plus.n8 a_n2072_n1288# 0.077381f
C61 plus.n9 a_n2072_n1288# 0.177988f
C62 plus.n10 a_n2072_n1288# 0.031315f
C63 plus.t2 a_n2072_n1288# 0.116278f
C64 plus.n11 a_n2072_n1288# 0.039089f
C65 plus.t1 a_n2072_n1288# 0.116278f
C66 plus.n12 a_n2072_n1288# 0.144015f
C67 plus.t9 a_n2072_n1288# 0.116278f
C68 plus.t7 a_n2072_n1288# 0.130356f
C69 plus.n13 a_n2072_n1288# 0.069028f
C70 plus.t0 a_n2072_n1288# 0.116278f
C71 plus.n14 a_n2072_n1288# 0.085322f
C72 plus.n15 a_n2072_n1288# 0.08589f
C73 plus.n16 a_n2072_n1288# 0.084298f
C74 plus.n17 a_n2072_n1288# 0.005325f
C75 plus.n18 a_n2072_n1288# 0.077381f
C76 plus.n19 a_n2072_n1288# 0.57176f
C77 source.n0 a_n2072_n1288# 0.032727f
C78 source.n1 a_n2072_n1288# 0.072411f
C79 source.t7 a_n2072_n1288# 0.054341f
C80 source.n2 a_n2072_n1288# 0.056672f
C81 source.n3 a_n2072_n1288# 0.018269f
C82 source.n4 a_n2072_n1288# 0.012049f
C83 source.n5 a_n2072_n1288# 0.159613f
C84 source.n6 a_n2072_n1288# 0.035876f
C85 source.n7 a_n2072_n1288# 0.393673f
C86 source.t4 a_n2072_n1288# 0.035437f
C87 source.t8 a_n2072_n1288# 0.035437f
C88 source.n8 a_n2072_n1288# 0.189447f
C89 source.n9 a_n2072_n1288# 0.315083f
C90 source.t0 a_n2072_n1288# 0.035437f
C91 source.t5 a_n2072_n1288# 0.035437f
C92 source.n10 a_n2072_n1288# 0.189447f
C93 source.n11 a_n2072_n1288# 0.313838f
C94 source.n12 a_n2072_n1288# 0.032727f
C95 source.n13 a_n2072_n1288# 0.072411f
C96 source.t14 a_n2072_n1288# 0.054341f
C97 source.n14 a_n2072_n1288# 0.056672f
C98 source.n15 a_n2072_n1288# 0.018269f
C99 source.n16 a_n2072_n1288# 0.012049f
C100 source.n17 a_n2072_n1288# 0.159613f
C101 source.n18 a_n2072_n1288# 0.035876f
C102 source.n19 a_n2072_n1288# 0.157975f
C103 source.t16 a_n2072_n1288# 0.035437f
C104 source.t15 a_n2072_n1288# 0.035437f
C105 source.n20 a_n2072_n1288# 0.189447f
C106 source.n21 a_n2072_n1288# 0.315083f
C107 source.t11 a_n2072_n1288# 0.035437f
C108 source.t12 a_n2072_n1288# 0.035437f
C109 source.n22 a_n2072_n1288# 0.189447f
C110 source.n23 a_n2072_n1288# 0.836108f
C111 source.t2 a_n2072_n1288# 0.035437f
C112 source.t3 a_n2072_n1288# 0.035437f
C113 source.n24 a_n2072_n1288# 0.189446f
C114 source.n25 a_n2072_n1288# 0.836109f
C115 source.t1 a_n2072_n1288# 0.035437f
C116 source.t19 a_n2072_n1288# 0.035437f
C117 source.n26 a_n2072_n1288# 0.189446f
C118 source.n27 a_n2072_n1288# 0.315085f
C119 source.n28 a_n2072_n1288# 0.032727f
C120 source.n29 a_n2072_n1288# 0.072411f
C121 source.t6 a_n2072_n1288# 0.054341f
C122 source.n30 a_n2072_n1288# 0.056672f
C123 source.n31 a_n2072_n1288# 0.018269f
C124 source.n32 a_n2072_n1288# 0.012049f
C125 source.n33 a_n2072_n1288# 0.159613f
C126 source.n34 a_n2072_n1288# 0.035876f
C127 source.n35 a_n2072_n1288# 0.157975f
C128 source.t10 a_n2072_n1288# 0.035437f
C129 source.t18 a_n2072_n1288# 0.035437f
C130 source.n36 a_n2072_n1288# 0.189446f
C131 source.n37 a_n2072_n1288# 0.313839f
C132 source.t9 a_n2072_n1288# 0.035437f
C133 source.t17 a_n2072_n1288# 0.035437f
C134 source.n38 a_n2072_n1288# 0.189446f
C135 source.n39 a_n2072_n1288# 0.315085f
C136 source.n40 a_n2072_n1288# 0.032727f
C137 source.n41 a_n2072_n1288# 0.072411f
C138 source.t13 a_n2072_n1288# 0.054341f
C139 source.n42 a_n2072_n1288# 0.056672f
C140 source.n43 a_n2072_n1288# 0.018269f
C141 source.n44 a_n2072_n1288# 0.012049f
C142 source.n45 a_n2072_n1288# 0.159613f
C143 source.n46 a_n2072_n1288# 0.035876f
C144 source.n47 a_n2072_n1288# 0.273899f
C145 source.n48 a_n2072_n1288# 0.568106f
C146 drain_right.n0 a_n2072_n1288# 0.026103f
C147 drain_right.n1 a_n2072_n1288# 0.057756f
C148 drain_right.t9 a_n2072_n1288# 0.043343f
C149 drain_right.n2 a_n2072_n1288# 0.045202f
C150 drain_right.n3 a_n2072_n1288# 0.014571f
C151 drain_right.n4 a_n2072_n1288# 0.00961f
C152 drain_right.n5 a_n2072_n1288# 0.127309f
C153 drain_right.n6 a_n2072_n1288# 0.042759f
C154 drain_right.t1 a_n2072_n1288# 0.028265f
C155 drain_right.t5 a_n2072_n1288# 0.028265f
C156 drain_right.n7 a_n2072_n1288# 0.177571f
C157 drain_right.n8 a_n2072_n1288# 0.294295f
C158 drain_right.t6 a_n2072_n1288# 0.028265f
C159 drain_right.t4 a_n2072_n1288# 0.028265f
C160 drain_right.n9 a_n2072_n1288# 0.179166f
C161 drain_right.n10 a_n2072_n1288# 0.773234f
C162 drain_right.t3 a_n2072_n1288# 0.028265f
C163 drain_right.t2 a_n2072_n1288# 0.028265f
C164 drain_right.n11 a_n2072_n1288# 0.180025f
C165 drain_right.t0 a_n2072_n1288# 0.028265f
C166 drain_right.t7 a_n2072_n1288# 0.028265f
C167 drain_right.n12 a_n2072_n1288# 0.177572f
C168 drain_right.n13 a_n2072_n1288# 0.503061f
C169 drain_right.n14 a_n2072_n1288# 0.026103f
C170 drain_right.n15 a_n2072_n1288# 0.057756f
C171 drain_right.t8 a_n2072_n1288# 0.043343f
C172 drain_right.n16 a_n2072_n1288# 0.045202f
C173 drain_right.n17 a_n2072_n1288# 0.014571f
C174 drain_right.n18 a_n2072_n1288# 0.00961f
C175 drain_right.n19 a_n2072_n1288# 0.127309f
C176 drain_right.n20 a_n2072_n1288# 0.040972f
C177 drain_right.n21 a_n2072_n1288# 0.258126f
C178 minus.n0 a_n2072_n1288# 0.030939f
C179 minus.t2 a_n2072_n1288# 0.11488f
C180 minus.n1 a_n2072_n1288# 0.084857f
C181 minus.t6 a_n2072_n1288# 0.11488f
C182 minus.t4 a_n2072_n1288# 0.128788f
C183 minus.t3 a_n2072_n1288# 0.11488f
C184 minus.n2 a_n2072_n1288# 0.084296f
C185 minus.n3 a_n2072_n1288# 0.068198f
C186 minus.n4 a_n2072_n1288# 0.142284f
C187 minus.n5 a_n2072_n1288# 0.038619f
C188 minus.n6 a_n2072_n1288# 0.083285f
C189 minus.n7 a_n2072_n1288# 0.005261f
C190 minus.t7 a_n2072_n1288# 0.11488f
C191 minus.n8 a_n2072_n1288# 0.076451f
C192 minus.n9 a_n2072_n1288# 0.592307f
C193 minus.n10 a_n2072_n1288# 0.030939f
C194 minus.t9 a_n2072_n1288# 0.11488f
C195 minus.n11 a_n2072_n1288# 0.084857f
C196 minus.t8 a_n2072_n1288# 0.128788f
C197 minus.t0 a_n2072_n1288# 0.11488f
C198 minus.n12 a_n2072_n1288# 0.084296f
C199 minus.n13 a_n2072_n1288# 0.068198f
C200 minus.n14 a_n2072_n1288# 0.142284f
C201 minus.n15 a_n2072_n1288# 0.038619f
C202 minus.t1 a_n2072_n1288# 0.11488f
C203 minus.n16 a_n2072_n1288# 0.083285f
C204 minus.n17 a_n2072_n1288# 0.005261f
C205 minus.t5 a_n2072_n1288# 0.11488f
C206 minus.n18 a_n2072_n1288# 0.076451f
C207 minus.n19 a_n2072_n1288# 0.161153f
C208 minus.n20 a_n2072_n1288# 0.726315f
.ends

