* NGSPICE file created from diffpair145.ext - technology: sky130A

.subckt diffpair145 minus drain_right drain_left source plus
X0 source.t21 plus.t0 drain_left.t7 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X1 source.t1 minus.t0 drain_right.t11 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X2 drain_right.t10 minus.t1 source.t23 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X3 drain_left.t3 plus.t1 source.t20 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X4 source.t19 plus.t2 drain_left.t9 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X5 source.t18 plus.t3 drain_left.t11 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X6 drain_left.t10 plus.t4 source.t17 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X7 source.t16 plus.t5 drain_left.t5 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X8 drain_right.t9 minus.t2 source.t5 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X9 a_n2158_n1288# a_n2158_n1288# a_n2158_n1288# a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.7
X10 drain_right.t8 minus.t3 source.t4 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X11 drain_left.t6 plus.t6 source.t15 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X12 source.t14 plus.t7 drain_left.t8 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X13 drain_left.t4 plus.t8 source.t13 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X14 drain_right.t7 minus.t4 source.t22 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X15 a_n2158_n1288# a_n2158_n1288# a_n2158_n1288# a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X16 drain_right.t6 minus.t5 source.t9 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X17 source.t7 minus.t6 drain_right.t5 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X18 drain_left.t1 plus.t9 source.t12 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X19 drain_right.t4 minus.t7 source.t6 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X20 source.t3 minus.t8 drain_right.t3 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X21 source.t0 minus.t9 drain_right.t2 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X22 source.t11 plus.t10 drain_left.t0 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X23 drain_left.t2 plus.t11 source.t10 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.7
X24 source.t8 minus.t10 drain_right.t1 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.7
X25 source.t2 minus.t11 drain_right.t0 a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.7
X26 a_n2158_n1288# a_n2158_n1288# a_n2158_n1288# a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
X27 a_n2158_n1288# a_n2158_n1288# a_n2158_n1288# a_n2158_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.7
R0 plus.n7 plus.n6 161.3
R1 plus.n8 plus.n3 161.3
R2 plus.n10 plus.n9 161.3
R3 plus.n11 plus.n2 161.3
R4 plus.n13 plus.n12 161.3
R5 plus.n14 plus.n1 161.3
R6 plus.n15 plus.n0 161.3
R7 plus.n17 plus.n16 161.3
R8 plus.n25 plus.n24 161.3
R9 plus.n26 plus.n21 161.3
R10 plus.n28 plus.n27 161.3
R11 plus.n29 plus.n20 161.3
R12 plus.n31 plus.n30 161.3
R13 plus.n32 plus.n19 161.3
R14 plus.n33 plus.n18 161.3
R15 plus.n35 plus.n34 161.3
R16 plus.n5 plus.t3 148.28
R17 plus.n23 plus.t11 148.28
R18 plus.n16 plus.t8 124.977
R19 plus.n14 plus.t2 124.977
R20 plus.n2 plus.t6 124.977
R21 plus.n8 plus.t0 124.977
R22 plus.n4 plus.t9 124.977
R23 plus.n34 plus.t7 124.977
R24 plus.n32 plus.t4 124.977
R25 plus.n20 plus.t5 124.977
R26 plus.n26 plus.t1 124.977
R27 plus.n22 plus.t10 124.977
R28 plus.n6 plus.n5 44.8907
R29 plus.n24 plus.n23 44.8907
R30 plus.n16 plus.n15 32.8641
R31 plus.n34 plus.n33 32.8641
R32 plus.n14 plus.n13 28.4823
R33 plus.n7 plus.n4 28.4823
R34 plus.n32 plus.n31 28.4823
R35 plus.n25 plus.n22 28.4823
R36 plus plus.n35 27.5331
R37 plus.n9 plus.n8 24.1005
R38 plus.n9 plus.n2 24.1005
R39 plus.n27 plus.n20 24.1005
R40 plus.n27 plus.n26 24.1005
R41 plus.n13 plus.n2 19.7187
R42 plus.n8 plus.n7 19.7187
R43 plus.n31 plus.n20 19.7187
R44 plus.n26 plus.n25 19.7187
R45 plus.n5 plus.n4 18.4104
R46 plus.n23 plus.n22 18.4104
R47 plus.n15 plus.n14 15.3369
R48 plus.n33 plus.n32 15.3369
R49 plus plus.n17 8.5005
R50 plus.n6 plus.n3 0.189894
R51 plus.n10 plus.n3 0.189894
R52 plus.n11 plus.n10 0.189894
R53 plus.n12 plus.n11 0.189894
R54 plus.n12 plus.n1 0.189894
R55 plus.n1 plus.n0 0.189894
R56 plus.n17 plus.n0 0.189894
R57 plus.n35 plus.n18 0.189894
R58 plus.n19 plus.n18 0.189894
R59 plus.n30 plus.n19 0.189894
R60 plus.n30 plus.n29 0.189894
R61 plus.n29 plus.n28 0.189894
R62 plus.n28 plus.n21 0.189894
R63 plus.n24 plus.n21 0.189894
R64 drain_left.n6 drain_left.n4 101.683
R65 drain_left.n3 drain_left.n2 101.629
R66 drain_left.n3 drain_left.n0 101.629
R67 drain_left.n8 drain_left.n7 100.796
R68 drain_left.n6 drain_left.n5 100.796
R69 drain_left.n3 drain_left.n1 100.796
R70 drain_left drain_left.n3 24.231
R71 drain_left.n1 drain_left.t5 9.9005
R72 drain_left.n1 drain_left.t3 9.9005
R73 drain_left.n2 drain_left.t0 9.9005
R74 drain_left.n2 drain_left.t2 9.9005
R75 drain_left.n0 drain_left.t8 9.9005
R76 drain_left.n0 drain_left.t10 9.9005
R77 drain_left.n7 drain_left.t9 9.9005
R78 drain_left.n7 drain_left.t4 9.9005
R79 drain_left.n5 drain_left.t7 9.9005
R80 drain_left.n5 drain_left.t6 9.9005
R81 drain_left.n4 drain_left.t11 9.9005
R82 drain_left.n4 drain_left.t1 9.9005
R83 drain_left drain_left.n8 6.54115
R84 drain_left.n8 drain_left.n6 0.888431
R85 source.n74 source.n72 289.615
R86 source.n62 source.n60 289.615
R87 source.n54 source.n52 289.615
R88 source.n42 source.n40 289.615
R89 source.n2 source.n0 289.615
R90 source.n14 source.n12 289.615
R91 source.n22 source.n20 289.615
R92 source.n34 source.n32 289.615
R93 source.n75 source.n74 185
R94 source.n63 source.n62 185
R95 source.n55 source.n54 185
R96 source.n43 source.n42 185
R97 source.n3 source.n2 185
R98 source.n15 source.n14 185
R99 source.n23 source.n22 185
R100 source.n35 source.n34 185
R101 source.t23 source.n73 167.117
R102 source.t7 source.n61 167.117
R103 source.t10 source.n53 167.117
R104 source.t14 source.n41 167.117
R105 source.t13 source.n1 167.117
R106 source.t18 source.n13 167.117
R107 source.t9 source.n21 167.117
R108 source.t2 source.n33 167.117
R109 source.n9 source.n8 84.1169
R110 source.n11 source.n10 84.1169
R111 source.n29 source.n28 84.1169
R112 source.n31 source.n30 84.1169
R113 source.n71 source.n70 84.1168
R114 source.n69 source.n68 84.1168
R115 source.n51 source.n50 84.1168
R116 source.n49 source.n48 84.1168
R117 source.n74 source.t23 52.3082
R118 source.n62 source.t7 52.3082
R119 source.n54 source.t10 52.3082
R120 source.n42 source.t14 52.3082
R121 source.n2 source.t13 52.3082
R122 source.n14 source.t18 52.3082
R123 source.n22 source.t9 52.3082
R124 source.n34 source.t2 52.3082
R125 source.n79 source.n78 31.4096
R126 source.n67 source.n66 31.4096
R127 source.n59 source.n58 31.4096
R128 source.n47 source.n46 31.4096
R129 source.n7 source.n6 31.4096
R130 source.n19 source.n18 31.4096
R131 source.n27 source.n26 31.4096
R132 source.n39 source.n38 31.4096
R133 source.n47 source.n39 14.5999
R134 source.n70 source.t6 9.9005
R135 source.n70 source.t0 9.9005
R136 source.n68 source.t22 9.9005
R137 source.n68 source.t3 9.9005
R138 source.n50 source.t20 9.9005
R139 source.n50 source.t11 9.9005
R140 source.n48 source.t17 9.9005
R141 source.n48 source.t16 9.9005
R142 source.n8 source.t15 9.9005
R143 source.n8 source.t19 9.9005
R144 source.n10 source.t12 9.9005
R145 source.n10 source.t21 9.9005
R146 source.n28 source.t4 9.9005
R147 source.n28 source.t1 9.9005
R148 source.n30 source.t5 9.9005
R149 source.n30 source.t8 9.9005
R150 source.n75 source.n73 9.71174
R151 source.n63 source.n61 9.71174
R152 source.n55 source.n53 9.71174
R153 source.n43 source.n41 9.71174
R154 source.n3 source.n1 9.71174
R155 source.n15 source.n13 9.71174
R156 source.n23 source.n21 9.71174
R157 source.n35 source.n33 9.71174
R158 source.n78 source.n77 9.45567
R159 source.n66 source.n65 9.45567
R160 source.n58 source.n57 9.45567
R161 source.n46 source.n45 9.45567
R162 source.n6 source.n5 9.45567
R163 source.n18 source.n17 9.45567
R164 source.n26 source.n25 9.45567
R165 source.n38 source.n37 9.45567
R166 source.n77 source.n76 9.3005
R167 source.n65 source.n64 9.3005
R168 source.n57 source.n56 9.3005
R169 source.n45 source.n44 9.3005
R170 source.n5 source.n4 9.3005
R171 source.n17 source.n16 9.3005
R172 source.n25 source.n24 9.3005
R173 source.n37 source.n36 9.3005
R174 source.n80 source.n7 8.893
R175 source.n78 source.n72 8.14595
R176 source.n66 source.n60 8.14595
R177 source.n58 source.n52 8.14595
R178 source.n46 source.n40 8.14595
R179 source.n6 source.n0 8.14595
R180 source.n18 source.n12 8.14595
R181 source.n26 source.n20 8.14595
R182 source.n38 source.n32 8.14595
R183 source.n76 source.n75 7.3702
R184 source.n64 source.n63 7.3702
R185 source.n56 source.n55 7.3702
R186 source.n44 source.n43 7.3702
R187 source.n4 source.n3 7.3702
R188 source.n16 source.n15 7.3702
R189 source.n24 source.n23 7.3702
R190 source.n36 source.n35 7.3702
R191 source.n76 source.n72 5.81868
R192 source.n64 source.n60 5.81868
R193 source.n56 source.n52 5.81868
R194 source.n44 source.n40 5.81868
R195 source.n4 source.n0 5.81868
R196 source.n16 source.n12 5.81868
R197 source.n24 source.n20 5.81868
R198 source.n36 source.n32 5.81868
R199 source.n80 source.n79 5.7074
R200 source.n77 source.n73 3.44771
R201 source.n65 source.n61 3.44771
R202 source.n57 source.n53 3.44771
R203 source.n45 source.n41 3.44771
R204 source.n5 source.n1 3.44771
R205 source.n17 source.n13 3.44771
R206 source.n25 source.n21 3.44771
R207 source.n37 source.n33 3.44771
R208 source.n39 source.n31 0.888431
R209 source.n31 source.n29 0.888431
R210 source.n29 source.n27 0.888431
R211 source.n19 source.n11 0.888431
R212 source.n11 source.n9 0.888431
R213 source.n9 source.n7 0.888431
R214 source.n49 source.n47 0.888431
R215 source.n51 source.n49 0.888431
R216 source.n59 source.n51 0.888431
R217 source.n69 source.n67 0.888431
R218 source.n71 source.n69 0.888431
R219 source.n79 source.n71 0.888431
R220 source.n27 source.n19 0.470328
R221 source.n67 source.n59 0.470328
R222 source source.n80 0.188
R223 minus.n17 minus.n16 161.3
R224 minus.n15 minus.n0 161.3
R225 minus.n14 minus.n13 161.3
R226 minus.n12 minus.n1 161.3
R227 minus.n11 minus.n10 161.3
R228 minus.n9 minus.n2 161.3
R229 minus.n8 minus.n7 161.3
R230 minus.n6 minus.n3 161.3
R231 minus.n35 minus.n34 161.3
R232 minus.n33 minus.n18 161.3
R233 minus.n32 minus.n31 161.3
R234 minus.n30 minus.n19 161.3
R235 minus.n29 minus.n28 161.3
R236 minus.n27 minus.n20 161.3
R237 minus.n26 minus.n25 161.3
R238 minus.n24 minus.n21 161.3
R239 minus.n5 minus.t5 148.28
R240 minus.n23 minus.t6 148.28
R241 minus.n4 minus.t0 124.977
R242 minus.n8 minus.t3 124.977
R243 minus.n10 minus.t10 124.977
R244 minus.n14 minus.t2 124.977
R245 minus.n16 minus.t11 124.977
R246 minus.n22 minus.t4 124.977
R247 minus.n26 minus.t8 124.977
R248 minus.n28 minus.t7 124.977
R249 minus.n32 minus.t9 124.977
R250 minus.n34 minus.t1 124.977
R251 minus.n6 minus.n5 44.8907
R252 minus.n24 minus.n23 44.8907
R253 minus.n16 minus.n15 32.8641
R254 minus.n34 minus.n33 32.8641
R255 minus.n36 minus.n17 29.8641
R256 minus.n4 minus.n3 28.4823
R257 minus.n14 minus.n1 28.4823
R258 minus.n22 minus.n21 28.4823
R259 minus.n32 minus.n19 28.4823
R260 minus.n10 minus.n9 24.1005
R261 minus.n9 minus.n8 24.1005
R262 minus.n27 minus.n26 24.1005
R263 minus.n28 minus.n27 24.1005
R264 minus.n8 minus.n3 19.7187
R265 minus.n10 minus.n1 19.7187
R266 minus.n26 minus.n21 19.7187
R267 minus.n28 minus.n19 19.7187
R268 minus.n5 minus.n4 18.4104
R269 minus.n23 minus.n22 18.4104
R270 minus.n15 minus.n14 15.3369
R271 minus.n33 minus.n32 15.3369
R272 minus.n36 minus.n35 6.64444
R273 minus.n17 minus.n0 0.189894
R274 minus.n13 minus.n0 0.189894
R275 minus.n13 minus.n12 0.189894
R276 minus.n12 minus.n11 0.189894
R277 minus.n11 minus.n2 0.189894
R278 minus.n7 minus.n2 0.189894
R279 minus.n7 minus.n6 0.189894
R280 minus.n25 minus.n24 0.189894
R281 minus.n25 minus.n20 0.189894
R282 minus.n29 minus.n20 0.189894
R283 minus.n30 minus.n29 0.189894
R284 minus.n31 minus.n30 0.189894
R285 minus.n31 minus.n18 0.189894
R286 minus.n35 minus.n18 0.189894
R287 minus minus.n36 0.188
R288 drain_right.n6 drain_right.n4 101.683
R289 drain_right.n3 drain_right.n2 101.629
R290 drain_right.n3 drain_right.n0 101.629
R291 drain_right.n6 drain_right.n5 100.796
R292 drain_right.n8 drain_right.n7 100.796
R293 drain_right.n3 drain_right.n1 100.796
R294 drain_right drain_right.n3 23.6777
R295 drain_right.n1 drain_right.t3 9.9005
R296 drain_right.n1 drain_right.t4 9.9005
R297 drain_right.n2 drain_right.t2 9.9005
R298 drain_right.n2 drain_right.t10 9.9005
R299 drain_right.n0 drain_right.t5 9.9005
R300 drain_right.n0 drain_right.t7 9.9005
R301 drain_right.n4 drain_right.t11 9.9005
R302 drain_right.n4 drain_right.t6 9.9005
R303 drain_right.n5 drain_right.t1 9.9005
R304 drain_right.n5 drain_right.t8 9.9005
R305 drain_right.n7 drain_right.t0 9.9005
R306 drain_right.n7 drain_right.t9 9.9005
R307 drain_right drain_right.n8 6.54115
R308 drain_right.n8 drain_right.n6 0.888431
C0 plus drain_right 0.373454f
C1 source drain_left 4.92681f
C2 drain_left minus 0.177688f
C3 source plus 2.16734f
C4 plus minus 3.99068f
C5 source drain_right 4.92885f
C6 drain_right minus 1.72949f
C7 source minus 2.15338f
C8 plus drain_left 1.94117f
C9 drain_left drain_right 1.08515f
C10 drain_right a_n2158_n1288# 3.81703f
C11 drain_left a_n2158_n1288# 4.08709f
C12 source a_n2158_n1288# 3.215412f
C13 minus a_n2158_n1288# 7.686388f
C14 plus a_n2158_n1288# 8.5856f
C15 drain_right.t5 a_n2158_n1288# 0.030499f
C16 drain_right.t7 a_n2158_n1288# 0.030499f
C17 drain_right.n0 a_n2158_n1288# 0.193759f
C18 drain_right.t3 a_n2158_n1288# 0.030499f
C19 drain_right.t4 a_n2158_n1288# 0.030499f
C20 drain_right.n1 a_n2158_n1288# 0.191605f
C21 drain_right.t2 a_n2158_n1288# 0.030499f
C22 drain_right.t10 a_n2158_n1288# 0.030499f
C23 drain_right.n2 a_n2158_n1288# 0.193759f
C24 drain_right.n3 a_n2158_n1288# 1.31625f
C25 drain_right.t11 a_n2158_n1288# 0.030499f
C26 drain_right.t6 a_n2158_n1288# 0.030499f
C27 drain_right.n4 a_n2158_n1288# 0.193927f
C28 drain_right.t1 a_n2158_n1288# 0.030499f
C29 drain_right.t8 a_n2158_n1288# 0.030499f
C30 drain_right.n5 a_n2158_n1288# 0.191605f
C31 drain_right.n6 a_n2158_n1288# 0.521704f
C32 drain_right.t0 a_n2158_n1288# 0.030499f
C33 drain_right.t9 a_n2158_n1288# 0.030499f
C34 drain_right.n7 a_n2158_n1288# 0.191605f
C35 drain_right.n8 a_n2158_n1288# 0.428815f
C36 minus.n0 a_n2158_n1288# 0.03522f
C37 minus.n1 a_n2158_n1288# 0.007992f
C38 minus.t2 a_n2158_n1288# 0.152695f
C39 minus.n2 a_n2158_n1288# 0.03522f
C40 minus.n3 a_n2158_n1288# 0.007992f
C41 minus.t3 a_n2158_n1288# 0.152695f
C42 minus.t5 a_n2158_n1288# 0.169369f
C43 minus.t0 a_n2158_n1288# 0.152695f
C44 minus.n4 a_n2158_n1288# 0.110082f
C45 minus.n5 a_n2158_n1288# 0.092622f
C46 minus.n6 a_n2158_n1288# 0.147753f
C47 minus.n7 a_n2158_n1288# 0.03522f
C48 minus.n8 a_n2158_n1288# 0.106143f
C49 minus.n9 a_n2158_n1288# 0.007992f
C50 minus.t10 a_n2158_n1288# 0.152695f
C51 minus.n10 a_n2158_n1288# 0.106143f
C52 minus.n11 a_n2158_n1288# 0.03522f
C53 minus.n12 a_n2158_n1288# 0.03522f
C54 minus.n13 a_n2158_n1288# 0.03522f
C55 minus.n14 a_n2158_n1288# 0.106143f
C56 minus.n15 a_n2158_n1288# 0.007992f
C57 minus.t11 a_n2158_n1288# 0.152695f
C58 minus.n16 a_n2158_n1288# 0.104515f
C59 minus.n17 a_n2158_n1288# 0.913901f
C60 minus.n18 a_n2158_n1288# 0.03522f
C61 minus.n19 a_n2158_n1288# 0.007992f
C62 minus.n20 a_n2158_n1288# 0.03522f
C63 minus.n21 a_n2158_n1288# 0.007992f
C64 minus.t6 a_n2158_n1288# 0.169369f
C65 minus.t4 a_n2158_n1288# 0.152695f
C66 minus.n22 a_n2158_n1288# 0.110082f
C67 minus.n23 a_n2158_n1288# 0.092622f
C68 minus.n24 a_n2158_n1288# 0.147753f
C69 minus.n25 a_n2158_n1288# 0.03522f
C70 minus.t8 a_n2158_n1288# 0.152695f
C71 minus.n26 a_n2158_n1288# 0.106143f
C72 minus.n27 a_n2158_n1288# 0.007992f
C73 minus.t7 a_n2158_n1288# 0.152695f
C74 minus.n28 a_n2158_n1288# 0.106143f
C75 minus.n29 a_n2158_n1288# 0.03522f
C76 minus.n30 a_n2158_n1288# 0.03522f
C77 minus.n31 a_n2158_n1288# 0.03522f
C78 minus.t9 a_n2158_n1288# 0.152695f
C79 minus.n32 a_n2158_n1288# 0.106143f
C80 minus.n33 a_n2158_n1288# 0.007992f
C81 minus.t1 a_n2158_n1288# 0.152695f
C82 minus.n34 a_n2158_n1288# 0.104515f
C83 minus.n35 a_n2158_n1288# 0.242165f
C84 minus.n36 a_n2158_n1288# 1.12174f
C85 source.n0 a_n2158_n1288# 0.042445f
C86 source.n1 a_n2158_n1288# 0.093914f
C87 source.t13 a_n2158_n1288# 0.070478f
C88 source.n2 a_n2158_n1288# 0.073501f
C89 source.n3 a_n2158_n1288# 0.023694f
C90 source.n4 a_n2158_n1288# 0.015627f
C91 source.n5 a_n2158_n1288# 0.207009f
C92 source.n6 a_n2158_n1288# 0.046529f
C93 source.n7 a_n2158_n1288# 0.496314f
C94 source.t15 a_n2158_n1288# 0.04596f
C95 source.t19 a_n2158_n1288# 0.04596f
C96 source.n8 a_n2158_n1288# 0.245703f
C97 source.n9 a_n2158_n1288# 0.392491f
C98 source.t12 a_n2158_n1288# 0.04596f
C99 source.t21 a_n2158_n1288# 0.04596f
C100 source.n10 a_n2158_n1288# 0.245703f
C101 source.n11 a_n2158_n1288# 0.392491f
C102 source.n12 a_n2158_n1288# 0.042445f
C103 source.n13 a_n2158_n1288# 0.093914f
C104 source.t18 a_n2158_n1288# 0.070478f
C105 source.n14 a_n2158_n1288# 0.073501f
C106 source.n15 a_n2158_n1288# 0.023694f
C107 source.n16 a_n2158_n1288# 0.015627f
C108 source.n17 a_n2158_n1288# 0.207009f
C109 source.n18 a_n2158_n1288# 0.046529f
C110 source.n19 a_n2158_n1288# 0.151167f
C111 source.n20 a_n2158_n1288# 0.042445f
C112 source.n21 a_n2158_n1288# 0.093914f
C113 source.t9 a_n2158_n1288# 0.070478f
C114 source.n22 a_n2158_n1288# 0.073501f
C115 source.n23 a_n2158_n1288# 0.023694f
C116 source.n24 a_n2158_n1288# 0.015627f
C117 source.n25 a_n2158_n1288# 0.207009f
C118 source.n26 a_n2158_n1288# 0.046529f
C119 source.n27 a_n2158_n1288# 0.151167f
C120 source.t4 a_n2158_n1288# 0.04596f
C121 source.t1 a_n2158_n1288# 0.04596f
C122 source.n28 a_n2158_n1288# 0.245703f
C123 source.n29 a_n2158_n1288# 0.392491f
C124 source.t5 a_n2158_n1288# 0.04596f
C125 source.t8 a_n2158_n1288# 0.04596f
C126 source.n30 a_n2158_n1288# 0.245703f
C127 source.n31 a_n2158_n1288# 0.392491f
C128 source.n32 a_n2158_n1288# 0.042445f
C129 source.n33 a_n2158_n1288# 0.093914f
C130 source.t2 a_n2158_n1288# 0.070478f
C131 source.n34 a_n2158_n1288# 0.073501f
C132 source.n35 a_n2158_n1288# 0.023694f
C133 source.n36 a_n2158_n1288# 0.015627f
C134 source.n37 a_n2158_n1288# 0.207009f
C135 source.n38 a_n2158_n1288# 0.046529f
C136 source.n39 a_n2158_n1288# 0.774806f
C137 source.n40 a_n2158_n1288# 0.042445f
C138 source.n41 a_n2158_n1288# 0.093914f
C139 source.t14 a_n2158_n1288# 0.070478f
C140 source.n42 a_n2158_n1288# 0.073501f
C141 source.n43 a_n2158_n1288# 0.023694f
C142 source.n44 a_n2158_n1288# 0.015627f
C143 source.n45 a_n2158_n1288# 0.207009f
C144 source.n46 a_n2158_n1288# 0.046529f
C145 source.n47 a_n2158_n1288# 0.774806f
C146 source.t17 a_n2158_n1288# 0.04596f
C147 source.t16 a_n2158_n1288# 0.04596f
C148 source.n48 a_n2158_n1288# 0.245701f
C149 source.n49 a_n2158_n1288# 0.392492f
C150 source.t20 a_n2158_n1288# 0.04596f
C151 source.t11 a_n2158_n1288# 0.04596f
C152 source.n50 a_n2158_n1288# 0.245701f
C153 source.n51 a_n2158_n1288# 0.392492f
C154 source.n52 a_n2158_n1288# 0.042445f
C155 source.n53 a_n2158_n1288# 0.093914f
C156 source.t10 a_n2158_n1288# 0.070478f
C157 source.n54 a_n2158_n1288# 0.073501f
C158 source.n55 a_n2158_n1288# 0.023694f
C159 source.n56 a_n2158_n1288# 0.015627f
C160 source.n57 a_n2158_n1288# 0.207009f
C161 source.n58 a_n2158_n1288# 0.046529f
C162 source.n59 a_n2158_n1288# 0.151167f
C163 source.n60 a_n2158_n1288# 0.042445f
C164 source.n61 a_n2158_n1288# 0.093914f
C165 source.t7 a_n2158_n1288# 0.070478f
C166 source.n62 a_n2158_n1288# 0.073501f
C167 source.n63 a_n2158_n1288# 0.023694f
C168 source.n64 a_n2158_n1288# 0.015627f
C169 source.n65 a_n2158_n1288# 0.207009f
C170 source.n66 a_n2158_n1288# 0.046529f
C171 source.n67 a_n2158_n1288# 0.151167f
C172 source.t22 a_n2158_n1288# 0.04596f
C173 source.t3 a_n2158_n1288# 0.04596f
C174 source.n68 a_n2158_n1288# 0.245701f
C175 source.n69 a_n2158_n1288# 0.392492f
C176 source.t6 a_n2158_n1288# 0.04596f
C177 source.t0 a_n2158_n1288# 0.04596f
C178 source.n70 a_n2158_n1288# 0.245701f
C179 source.n71 a_n2158_n1288# 0.392492f
C180 source.n72 a_n2158_n1288# 0.042445f
C181 source.n73 a_n2158_n1288# 0.093914f
C182 source.t23 a_n2158_n1288# 0.070478f
C183 source.n74 a_n2158_n1288# 0.073501f
C184 source.n75 a_n2158_n1288# 0.023694f
C185 source.n76 a_n2158_n1288# 0.015627f
C186 source.n77 a_n2158_n1288# 0.207009f
C187 source.n78 a_n2158_n1288# 0.046529f
C188 source.n79 a_n2158_n1288# 0.340859f
C189 source.n80 a_n2158_n1288# 0.733124f
C190 drain_left.t8 a_n2158_n1288# 0.030036f
C191 drain_left.t10 a_n2158_n1288# 0.030036f
C192 drain_left.n0 a_n2158_n1288# 0.190819f
C193 drain_left.t5 a_n2158_n1288# 0.030036f
C194 drain_left.t3 a_n2158_n1288# 0.030036f
C195 drain_left.n1 a_n2158_n1288# 0.188698f
C196 drain_left.t0 a_n2158_n1288# 0.030036f
C197 drain_left.t2 a_n2158_n1288# 0.030036f
C198 drain_left.n2 a_n2158_n1288# 0.190819f
C199 drain_left.n3 a_n2158_n1288# 1.3334f
C200 drain_left.t11 a_n2158_n1288# 0.030036f
C201 drain_left.t1 a_n2158_n1288# 0.030036f
C202 drain_left.n4 a_n2158_n1288# 0.190985f
C203 drain_left.t7 a_n2158_n1288# 0.030036f
C204 drain_left.t6 a_n2158_n1288# 0.030036f
C205 drain_left.n5 a_n2158_n1288# 0.188698f
C206 drain_left.n6 a_n2158_n1288# 0.513788f
C207 drain_left.t9 a_n2158_n1288# 0.030036f
C208 drain_left.t4 a_n2158_n1288# 0.030036f
C209 drain_left.n7 a_n2158_n1288# 0.188698f
C210 drain_left.n8 a_n2158_n1288# 0.422309f
C211 plus.n0 a_n2158_n1288# 0.03563f
C212 plus.t8 a_n2158_n1288# 0.154469f
C213 plus.t2 a_n2158_n1288# 0.154469f
C214 plus.n1 a_n2158_n1288# 0.03563f
C215 plus.t6 a_n2158_n1288# 0.154469f
C216 plus.n2 a_n2158_n1288# 0.107377f
C217 plus.n3 a_n2158_n1288# 0.03563f
C218 plus.t0 a_n2158_n1288# 0.154469f
C219 plus.t9 a_n2158_n1288# 0.154469f
C220 plus.n4 a_n2158_n1288# 0.111362f
C221 plus.t3 a_n2158_n1288# 0.171337f
C222 plus.n5 a_n2158_n1288# 0.093698f
C223 plus.n6 a_n2158_n1288# 0.14947f
C224 plus.n7 a_n2158_n1288# 0.008085f
C225 plus.n8 a_n2158_n1288# 0.107377f
C226 plus.n9 a_n2158_n1288# 0.008085f
C227 plus.n10 a_n2158_n1288# 0.03563f
C228 plus.n11 a_n2158_n1288# 0.03563f
C229 plus.n12 a_n2158_n1288# 0.03563f
C230 plus.n13 a_n2158_n1288# 0.008085f
C231 plus.n14 a_n2158_n1288# 0.107377f
C232 plus.n15 a_n2158_n1288# 0.008085f
C233 plus.n16 a_n2158_n1288# 0.105729f
C234 plus.n17 a_n2158_n1288# 0.267414f
C235 plus.n18 a_n2158_n1288# 0.03563f
C236 plus.t7 a_n2158_n1288# 0.154469f
C237 plus.n19 a_n2158_n1288# 0.03563f
C238 plus.t4 a_n2158_n1288# 0.154469f
C239 plus.t5 a_n2158_n1288# 0.154469f
C240 plus.n20 a_n2158_n1288# 0.107377f
C241 plus.n21 a_n2158_n1288# 0.03563f
C242 plus.t1 a_n2158_n1288# 0.154469f
C243 plus.t10 a_n2158_n1288# 0.154469f
C244 plus.n22 a_n2158_n1288# 0.111362f
C245 plus.t11 a_n2158_n1288# 0.171337f
C246 plus.n23 a_n2158_n1288# 0.093698f
C247 plus.n24 a_n2158_n1288# 0.14947f
C248 plus.n25 a_n2158_n1288# 0.008085f
C249 plus.n26 a_n2158_n1288# 0.107377f
C250 plus.n27 a_n2158_n1288# 0.008085f
C251 plus.n28 a_n2158_n1288# 0.03563f
C252 plus.n29 a_n2158_n1288# 0.03563f
C253 plus.n30 a_n2158_n1288# 0.03563f
C254 plus.n31 a_n2158_n1288# 0.008085f
C255 plus.n32 a_n2158_n1288# 0.107377f
C256 plus.n33 a_n2158_n1288# 0.008085f
C257 plus.n34 a_n2158_n1288# 0.105729f
C258 plus.n35 a_n2158_n1288# 0.881164f
.ends

