* NGSPICE file created from diffpair113.ext - technology: sky130A

.subckt diffpair113 minus drain_right drain_left source plus
X0 source.t14 minus.t0 drain_right.t0 a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X1 source.t15 plus.t0 drain_left.t7 a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X2 drain_right.t4 minus.t1 source.t13 a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X3 a_n1346_n1288# a_n1346_n1288# a_n1346_n1288# a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=6.24 ps=38.24 w=2 l=0.3
X4 drain_right.t5 minus.t2 source.t12 a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X5 source.t0 plus.t1 drain_left.t6 a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X6 a_n1346_n1288# a_n1346_n1288# a_n1346_n1288# a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X7 a_n1346_n1288# a_n1346_n1288# a_n1346_n1288# a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X8 drain_left.t5 plus.t2 source.t1 a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X9 drain_left.t4 plus.t3 source.t6 a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X10 source.t11 minus.t3 drain_right.t1 a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X11 source.t5 plus.t4 drain_left.t3 a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X12 source.t10 minus.t4 drain_right.t6 a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.3
X13 drain_right.t7 minus.t5 source.t9 a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X14 drain_right.t2 minus.t6 source.t8 a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X15 source.t2 plus.t5 drain_left.t2 a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X16 source.t7 minus.t7 drain_right.t3 a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.3
X17 drain_left.t1 plus.t6 source.t4 a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
X18 a_n1346_n1288# a_n1346_n1288# a_n1346_n1288# a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.3
X19 drain_left.t0 plus.t7 source.t3 a_n1346_n1288# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.3
R0 minus.n7 minus.t4 293.582
R1 minus.n2 minus.t5 293.582
R2 minus.n16 minus.t2 293.582
R3 minus.n11 minus.t0 293.582
R4 minus.n6 minus.t1 265.101
R5 minus.n1 minus.t7 265.101
R6 minus.n15 minus.t3 265.101
R7 minus.n10 minus.t6 265.101
R8 minus.n3 minus.n2 161.489
R9 minus.n12 minus.n11 161.489
R10 minus.n8 minus.n7 161.3
R11 minus.n5 minus.n0 161.3
R12 minus.n4 minus.n3 161.3
R13 minus.n17 minus.n16 161.3
R14 minus.n14 minus.n9 161.3
R15 minus.n13 minus.n12 161.3
R16 minus.n5 minus.n4 73.0308
R17 minus.n14 minus.n13 73.0308
R18 minus.n7 minus.n6 63.5369
R19 minus.n2 minus.n1 63.5369
R20 minus.n11 minus.n10 63.5369
R21 minus.n16 minus.n15 63.5369
R22 minus.n18 minus.n8 26.6066
R23 minus.n6 minus.n5 9.49444
R24 minus.n4 minus.n1 9.49444
R25 minus.n13 minus.n10 9.49444
R26 minus.n15 minus.n14 9.49444
R27 minus.n18 minus.n17 6.46262
R28 minus.n8 minus.n0 0.189894
R29 minus.n3 minus.n0 0.189894
R30 minus.n12 minus.n9 0.189894
R31 minus.n17 minus.n9 0.189894
R32 minus minus.n18 0.188
R33 drain_right.n5 drain_right.n3 101.338
R34 drain_right.n2 drain_right.n1 101.011
R35 drain_right.n2 drain_right.n0 101.011
R36 drain_right.n5 drain_right.n4 100.796
R37 drain_right drain_right.n2 21.1389
R38 drain_right.n1 drain_right.t1 9.9005
R39 drain_right.n1 drain_right.t5 9.9005
R40 drain_right.n0 drain_right.t0 9.9005
R41 drain_right.n0 drain_right.t2 9.9005
R42 drain_right.n3 drain_right.t3 9.9005
R43 drain_right.n3 drain_right.t7 9.9005
R44 drain_right.n4 drain_right.t6 9.9005
R45 drain_right.n4 drain_right.t4 9.9005
R46 drain_right drain_right.n5 6.19632
R47 source.n66 source.n64 289.615
R48 source.n56 source.n54 289.615
R49 source.n48 source.n46 289.615
R50 source.n38 source.n36 289.615
R51 source.n2 source.n0 289.615
R52 source.n12 source.n10 289.615
R53 source.n20 source.n18 289.615
R54 source.n30 source.n28 289.615
R55 source.n67 source.n66 185
R56 source.n57 source.n56 185
R57 source.n49 source.n48 185
R58 source.n39 source.n38 185
R59 source.n3 source.n2 185
R60 source.n13 source.n12 185
R61 source.n21 source.n20 185
R62 source.n31 source.n30 185
R63 source.t12 source.n65 167.117
R64 source.t14 source.n55 167.117
R65 source.t4 source.n47 167.117
R66 source.t15 source.n37 167.117
R67 source.t3 source.n1 167.117
R68 source.t0 source.n11 167.117
R69 source.t9 source.n19 167.117
R70 source.t10 source.n29 167.117
R71 source.n9 source.n8 84.1169
R72 source.n27 source.n26 84.1169
R73 source.n63 source.n62 84.1168
R74 source.n45 source.n44 84.1168
R75 source.n66 source.t12 52.3082
R76 source.n56 source.t14 52.3082
R77 source.n48 source.t4 52.3082
R78 source.n38 source.t15 52.3082
R79 source.n2 source.t3 52.3082
R80 source.n12 source.t0 52.3082
R81 source.n20 source.t9 52.3082
R82 source.n30 source.t10 52.3082
R83 source.n71 source.n70 31.4096
R84 source.n61 source.n60 31.4096
R85 source.n53 source.n52 31.4096
R86 source.n43 source.n42 31.4096
R87 source.n7 source.n6 31.4096
R88 source.n17 source.n16 31.4096
R89 source.n25 source.n24 31.4096
R90 source.n35 source.n34 31.4096
R91 source.n43 source.n35 14.2551
R92 source.n62 source.t8 9.9005
R93 source.n62 source.t11 9.9005
R94 source.n44 source.t1 9.9005
R95 source.n44 source.t5 9.9005
R96 source.n8 source.t6 9.9005
R97 source.n8 source.t2 9.9005
R98 source.n26 source.t13 9.9005
R99 source.n26 source.t7 9.9005
R100 source.n67 source.n65 9.71174
R101 source.n57 source.n55 9.71174
R102 source.n49 source.n47 9.71174
R103 source.n39 source.n37 9.71174
R104 source.n3 source.n1 9.71174
R105 source.n13 source.n11 9.71174
R106 source.n21 source.n19 9.71174
R107 source.n31 source.n29 9.71174
R108 source.n70 source.n69 9.45567
R109 source.n60 source.n59 9.45567
R110 source.n52 source.n51 9.45567
R111 source.n42 source.n41 9.45567
R112 source.n6 source.n5 9.45567
R113 source.n16 source.n15 9.45567
R114 source.n24 source.n23 9.45567
R115 source.n34 source.n33 9.45567
R116 source.n69 source.n68 9.3005
R117 source.n59 source.n58 9.3005
R118 source.n51 source.n50 9.3005
R119 source.n41 source.n40 9.3005
R120 source.n5 source.n4 9.3005
R121 source.n15 source.n14 9.3005
R122 source.n23 source.n22 9.3005
R123 source.n33 source.n32 9.3005
R124 source.n72 source.n7 8.72059
R125 source.n70 source.n64 8.14595
R126 source.n60 source.n54 8.14595
R127 source.n52 source.n46 8.14595
R128 source.n42 source.n36 8.14595
R129 source.n6 source.n0 8.14595
R130 source.n16 source.n10 8.14595
R131 source.n24 source.n18 8.14595
R132 source.n34 source.n28 8.14595
R133 source.n68 source.n67 7.3702
R134 source.n58 source.n57 7.3702
R135 source.n50 source.n49 7.3702
R136 source.n40 source.n39 7.3702
R137 source.n4 source.n3 7.3702
R138 source.n14 source.n13 7.3702
R139 source.n22 source.n21 7.3702
R140 source.n32 source.n31 7.3702
R141 source.n68 source.n64 5.81868
R142 source.n58 source.n54 5.81868
R143 source.n50 source.n46 5.81868
R144 source.n40 source.n36 5.81868
R145 source.n4 source.n0 5.81868
R146 source.n14 source.n10 5.81868
R147 source.n22 source.n18 5.81868
R148 source.n32 source.n28 5.81868
R149 source.n72 source.n71 5.53498
R150 source.n69 source.n65 3.44771
R151 source.n59 source.n55 3.44771
R152 source.n51 source.n47 3.44771
R153 source.n41 source.n37 3.44771
R154 source.n5 source.n1 3.44771
R155 source.n15 source.n11 3.44771
R156 source.n23 source.n19 3.44771
R157 source.n33 source.n29 3.44771
R158 source.n35 source.n27 0.543603
R159 source.n27 source.n25 0.543603
R160 source.n17 source.n9 0.543603
R161 source.n9 source.n7 0.543603
R162 source.n45 source.n43 0.543603
R163 source.n53 source.n45 0.543603
R164 source.n63 source.n61 0.543603
R165 source.n71 source.n63 0.543603
R166 source.n25 source.n17 0.470328
R167 source.n61 source.n53 0.470328
R168 source source.n72 0.188
R169 plus.n2 plus.t1 293.582
R170 plus.n7 plus.t7 293.582
R171 plus.n11 plus.t6 293.582
R172 plus.n16 plus.t0 293.582
R173 plus.n1 plus.t3 265.101
R174 plus.n6 plus.t5 265.101
R175 plus.n10 plus.t4 265.101
R176 plus.n15 plus.t2 265.101
R177 plus.n3 plus.n2 161.489
R178 plus.n12 plus.n11 161.489
R179 plus.n4 plus.n3 161.3
R180 plus.n5 plus.n0 161.3
R181 plus.n8 plus.n7 161.3
R182 plus.n13 plus.n12 161.3
R183 plus.n14 plus.n9 161.3
R184 plus.n17 plus.n16 161.3
R185 plus.n5 plus.n4 73.0308
R186 plus.n14 plus.n13 73.0308
R187 plus.n2 plus.n1 63.5369
R188 plus.n7 plus.n6 63.5369
R189 plus.n16 plus.n15 63.5369
R190 plus.n11 plus.n10 63.5369
R191 plus plus.n17 24.2755
R192 plus.n4 plus.n1 9.49444
R193 plus.n6 plus.n5 9.49444
R194 plus.n15 plus.n14 9.49444
R195 plus.n13 plus.n10 9.49444
R196 plus plus.n8 8.31868
R197 plus.n3 plus.n0 0.189894
R198 plus.n8 plus.n0 0.189894
R199 plus.n17 plus.n9 0.189894
R200 plus.n12 plus.n9 0.189894
R201 drain_left.n5 drain_left.n3 101.338
R202 drain_left.n2 drain_left.n1 101.011
R203 drain_left.n2 drain_left.n0 101.011
R204 drain_left.n5 drain_left.n4 100.796
R205 drain_left drain_left.n2 21.6922
R206 drain_left.n1 drain_left.t3 9.9005
R207 drain_left.n1 drain_left.t1 9.9005
R208 drain_left.n0 drain_left.t7 9.9005
R209 drain_left.n0 drain_left.t5 9.9005
R210 drain_left.n4 drain_left.t2 9.9005
R211 drain_left.n4 drain_left.t0 9.9005
R212 drain_left.n3 drain_left.t6 9.9005
R213 drain_left.n3 drain_left.t4 9.9005
R214 drain_left drain_left.n5 6.19632
C0 drain_left drain_right 0.630082f
C1 plus drain_right 0.28718f
C2 drain_left minus 0.176448f
C3 plus minus 2.98791f
C4 source drain_right 4.2789f
C5 plus drain_left 0.982145f
C6 source minus 0.931207f
C7 minus drain_right 0.854965f
C8 source drain_left 4.2797f
C9 source plus 0.94517f
C10 drain_right a_n1346_n1288# 3.11901f
C11 drain_left a_n1346_n1288# 3.28181f
C12 source a_n1346_n1288# 2.885341f
C13 minus a_n1346_n1288# 4.39489f
C14 plus a_n1346_n1288# 5.086843f
C15 drain_left.t7 a_n1346_n1288# 0.038065f
C16 drain_left.t5 a_n1346_n1288# 0.038065f
C17 drain_left.n0 a_n1346_n1288# 0.239683f
C18 drain_left.t3 a_n1346_n1288# 0.038065f
C19 drain_left.t1 a_n1346_n1288# 0.038065f
C20 drain_left.n1 a_n1346_n1288# 0.239683f
C21 drain_left.n2 a_n1346_n1288# 1.07934f
C22 drain_left.t6 a_n1346_n1288# 0.038065f
C23 drain_left.t4 a_n1346_n1288# 0.038065f
C24 drain_left.n3 a_n1346_n1288# 0.240628f
C25 drain_left.t2 a_n1346_n1288# 0.038065f
C26 drain_left.t0 a_n1346_n1288# 0.038065f
C27 drain_left.n4 a_n1346_n1288# 0.239137f
C28 drain_left.n5 a_n1346_n1288# 0.745957f
C29 plus.n0 a_n1346_n1288# 0.035105f
C30 plus.t5 a_n1346_n1288# 0.06198f
C31 plus.t3 a_n1346_n1288# 0.06198f
C32 plus.n1 a_n1346_n1288# 0.043288f
C33 plus.t1 a_n1346_n1288# 0.06617f
C34 plus.n2 a_n1346_n1288# 0.053496f
C35 plus.n3 a_n1346_n1288# 0.074277f
C36 plus.n4 a_n1346_n1288# 0.013052f
C37 plus.n5 a_n1346_n1288# 0.013052f
C38 plus.n6 a_n1346_n1288# 0.043288f
C39 plus.t7 a_n1346_n1288# 0.06617f
C40 plus.n7 a_n1346_n1288# 0.05345f
C41 plus.n8 a_n1346_n1288# 0.247702f
C42 plus.n9 a_n1346_n1288# 0.035105f
C43 plus.t0 a_n1346_n1288# 0.06617f
C44 plus.t2 a_n1346_n1288# 0.06198f
C45 plus.t4 a_n1346_n1288# 0.06198f
C46 plus.n10 a_n1346_n1288# 0.043288f
C47 plus.t6 a_n1346_n1288# 0.06617f
C48 plus.n11 a_n1346_n1288# 0.053496f
C49 plus.n12 a_n1346_n1288# 0.074277f
C50 plus.n13 a_n1346_n1288# 0.013052f
C51 plus.n14 a_n1346_n1288# 0.013052f
C52 plus.n15 a_n1346_n1288# 0.043288f
C53 plus.n16 a_n1346_n1288# 0.05345f
C54 plus.n17 a_n1346_n1288# 0.708366f
C55 source.n0 a_n1346_n1288# 0.034328f
C56 source.n1 a_n1346_n1288# 0.075955f
C57 source.t3 a_n1346_n1288# 0.057001f
C58 source.n2 a_n1346_n1288# 0.059446f
C59 source.n3 a_n1346_n1288# 0.019163f
C60 source.n4 a_n1346_n1288# 0.012638f
C61 source.n5 a_n1346_n1288# 0.167425f
C62 source.n6 a_n1346_n1288# 0.037632f
C63 source.n7 a_n1346_n1288# 0.355107f
C64 source.t6 a_n1346_n1288# 0.037172f
C65 source.t2 a_n1346_n1288# 0.037172f
C66 source.n8 a_n1346_n1288# 0.198719f
C67 source.n9 a_n1346_n1288# 0.265172f
C68 source.n10 a_n1346_n1288# 0.034328f
C69 source.n11 a_n1346_n1288# 0.075955f
C70 source.t0 a_n1346_n1288# 0.057001f
C71 source.n12 a_n1346_n1288# 0.059446f
C72 source.n13 a_n1346_n1288# 0.019163f
C73 source.n14 a_n1346_n1288# 0.012638f
C74 source.n15 a_n1346_n1288# 0.167425f
C75 source.n16 a_n1346_n1288# 0.037632f
C76 source.n17 a_n1346_n1288# 0.096128f
C77 source.n18 a_n1346_n1288# 0.034328f
C78 source.n19 a_n1346_n1288# 0.075955f
C79 source.t9 a_n1346_n1288# 0.057001f
C80 source.n20 a_n1346_n1288# 0.059446f
C81 source.n21 a_n1346_n1288# 0.019163f
C82 source.n22 a_n1346_n1288# 0.012638f
C83 source.n23 a_n1346_n1288# 0.167425f
C84 source.n24 a_n1346_n1288# 0.037632f
C85 source.n25 a_n1346_n1288# 0.096128f
C86 source.t13 a_n1346_n1288# 0.037172f
C87 source.t7 a_n1346_n1288# 0.037172f
C88 source.n26 a_n1346_n1288# 0.198719f
C89 source.n27 a_n1346_n1288# 0.265172f
C90 source.n28 a_n1346_n1288# 0.034328f
C91 source.n29 a_n1346_n1288# 0.075955f
C92 source.t10 a_n1346_n1288# 0.057001f
C93 source.n30 a_n1346_n1288# 0.059446f
C94 source.n31 a_n1346_n1288# 0.019163f
C95 source.n32 a_n1346_n1288# 0.012638f
C96 source.n33 a_n1346_n1288# 0.167425f
C97 source.n34 a_n1346_n1288# 0.037632f
C98 source.n35 a_n1346_n1288# 0.574381f
C99 source.n36 a_n1346_n1288# 0.034328f
C100 source.n37 a_n1346_n1288# 0.075955f
C101 source.t15 a_n1346_n1288# 0.057001f
C102 source.n38 a_n1346_n1288# 0.059446f
C103 source.n39 a_n1346_n1288# 0.019163f
C104 source.n40 a_n1346_n1288# 0.012638f
C105 source.n41 a_n1346_n1288# 0.167425f
C106 source.n42 a_n1346_n1288# 0.037632f
C107 source.n43 a_n1346_n1288# 0.574381f
C108 source.t1 a_n1346_n1288# 0.037172f
C109 source.t5 a_n1346_n1288# 0.037172f
C110 source.n44 a_n1346_n1288# 0.198718f
C111 source.n45 a_n1346_n1288# 0.265174f
C112 source.n46 a_n1346_n1288# 0.034328f
C113 source.n47 a_n1346_n1288# 0.075955f
C114 source.t4 a_n1346_n1288# 0.057001f
C115 source.n48 a_n1346_n1288# 0.059446f
C116 source.n49 a_n1346_n1288# 0.019163f
C117 source.n50 a_n1346_n1288# 0.012638f
C118 source.n51 a_n1346_n1288# 0.167425f
C119 source.n52 a_n1346_n1288# 0.037632f
C120 source.n53 a_n1346_n1288# 0.096128f
C121 source.n54 a_n1346_n1288# 0.034328f
C122 source.n55 a_n1346_n1288# 0.075955f
C123 source.t14 a_n1346_n1288# 0.057001f
C124 source.n56 a_n1346_n1288# 0.059446f
C125 source.n57 a_n1346_n1288# 0.019163f
C126 source.n58 a_n1346_n1288# 0.012638f
C127 source.n59 a_n1346_n1288# 0.167425f
C128 source.n60 a_n1346_n1288# 0.037632f
C129 source.n61 a_n1346_n1288# 0.096128f
C130 source.t8 a_n1346_n1288# 0.037172f
C131 source.t11 a_n1346_n1288# 0.037172f
C132 source.n62 a_n1346_n1288# 0.198718f
C133 source.n63 a_n1346_n1288# 0.265174f
C134 source.n64 a_n1346_n1288# 0.034328f
C135 source.n65 a_n1346_n1288# 0.075955f
C136 source.t12 a_n1346_n1288# 0.057001f
C137 source.n66 a_n1346_n1288# 0.059446f
C138 source.n67 a_n1346_n1288# 0.019163f
C139 source.n68 a_n1346_n1288# 0.012638f
C140 source.n69 a_n1346_n1288# 0.167425f
C141 source.n70 a_n1346_n1288# 0.037632f
C142 source.n71 a_n1346_n1288# 0.228895f
C143 source.n72 a_n1346_n1288# 0.581488f
C144 drain_right.t0 a_n1346_n1288# 0.038918f
C145 drain_right.t2 a_n1346_n1288# 0.038918f
C146 drain_right.n0 a_n1346_n1288# 0.245052f
C147 drain_right.t1 a_n1346_n1288# 0.038918f
C148 drain_right.t5 a_n1346_n1288# 0.038918f
C149 drain_right.n1 a_n1346_n1288# 0.245052f
C150 drain_right.n2 a_n1346_n1288# 1.05503f
C151 drain_right.t3 a_n1346_n1288# 0.038918f
C152 drain_right.t7 a_n1346_n1288# 0.038918f
C153 drain_right.n3 a_n1346_n1288# 0.246019f
C154 drain_right.t6 a_n1346_n1288# 0.038918f
C155 drain_right.t4 a_n1346_n1288# 0.038918f
C156 drain_right.n4 a_n1346_n1288# 0.244494f
C157 drain_right.n5 a_n1346_n1288# 0.762667f
C158 minus.n0 a_n1346_n1288# 0.034294f
C159 minus.t4 a_n1346_n1288# 0.06464f
C160 minus.t1 a_n1346_n1288# 0.060548f
C161 minus.t7 a_n1346_n1288# 0.060548f
C162 minus.n1 a_n1346_n1288# 0.042287f
C163 minus.t5 a_n1346_n1288# 0.06464f
C164 minus.n2 a_n1346_n1288# 0.052259f
C165 minus.n3 a_n1346_n1288# 0.07256f
C166 minus.n4 a_n1346_n1288# 0.012751f
C167 minus.n5 a_n1346_n1288# 0.012751f
C168 minus.n6 a_n1346_n1288# 0.042287f
C169 minus.n7 a_n1346_n1288# 0.052214f
C170 minus.n8 a_n1346_n1288# 0.72065f
C171 minus.n9 a_n1346_n1288# 0.034294f
C172 minus.t3 a_n1346_n1288# 0.060548f
C173 minus.t6 a_n1346_n1288# 0.060548f
C174 minus.n10 a_n1346_n1288# 0.042287f
C175 minus.t0 a_n1346_n1288# 0.06464f
C176 minus.n11 a_n1346_n1288# 0.052259f
C177 minus.n12 a_n1346_n1288# 0.07256f
C178 minus.n13 a_n1346_n1288# 0.012751f
C179 minus.n14 a_n1346_n1288# 0.012751f
C180 minus.n15 a_n1346_n1288# 0.042287f
C181 minus.t2 a_n1346_n1288# 0.06464f
C182 minus.n16 a_n1346_n1288# 0.052214f
C183 minus.n17 a_n1346_n1288# 0.221179f
C184 minus.n18 a_n1346_n1288# 0.892093f
.ends

