* NGSPICE file created from diffpair696.ext - technology: sky130A

.subckt diffpair696 minus drain_right drain_left source plus
X0 source.t27 plus.t0 drain_left.t5 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X1 drain_left.t4 plus.t1 source.t26 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.6
X2 source.t10 minus.t0 drain_right.t13 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X3 source.t25 plus.t2 drain_left.t1 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X4 drain_right.t12 minus.t1 source.t0 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X5 source.t9 minus.t2 drain_right.t11 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X6 drain_left.t0 plus.t3 source.t24 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X7 drain_right.t10 minus.t3 source.t12 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X8 drain_right.t9 minus.t4 source.t1 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.6
X9 source.t2 minus.t5 drain_right.t8 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X10 source.t23 plus.t4 drain_left.t3 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X11 drain_left.t2 plus.t5 source.t22 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X12 drain_right.t7 minus.t6 source.t3 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X13 source.t8 minus.t7 drain_right.t6 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X14 source.t21 plus.t6 drain_left.t7 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X15 drain_right.t5 minus.t8 source.t11 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X16 source.t20 plus.t7 drain_left.t6 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X17 source.t4 minus.t9 drain_right.t4 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X18 a_n2204_n5888# a_n2204_n5888# a_n2204_n5888# a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.6
X19 drain_left.t9 plus.t8 source.t19 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X20 drain_right.t3 minus.t10 source.t7 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.6
X21 drain_right.t2 minus.t11 source.t6 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.6
X22 source.t18 plus.t9 drain_left.t8 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X23 drain_left.t13 plus.t10 source.t17 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.6
X24 a_n2204_n5888# a_n2204_n5888# a_n2204_n5888# a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.6
X25 drain_right.t1 minus.t12 source.t13 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.6
X26 drain_left.t12 plus.t11 source.t16 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X27 drain_left.t11 plus.t12 source.t15 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.6
X28 a_n2204_n5888# a_n2204_n5888# a_n2204_n5888# a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.6
X29 a_n2204_n5888# a_n2204_n5888# a_n2204_n5888# a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.6
X30 source.t5 minus.t13 drain_right.t0 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.6
X31 drain_left.t10 plus.t13 source.t14 a_n2204_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.6
R0 plus.n5 plus.t10 1093.48
R1 plus.n23 plus.t13 1093.48
R2 plus.n16 plus.t1 1069.64
R3 plus.n14 plus.t2 1069.64
R4 plus.n2 plus.t5 1069.64
R5 plus.n9 plus.t7 1069.64
R6 plus.n8 plus.t8 1069.64
R7 plus.n4 plus.t9 1069.64
R8 plus.n34 plus.t12 1069.64
R9 plus.n32 plus.t4 1069.64
R10 plus.n20 plus.t3 1069.64
R11 plus.n27 plus.t0 1069.64
R12 plus.n26 plus.t11 1069.64
R13 plus.n22 plus.t6 1069.64
R14 plus.n7 plus.n6 161.3
R15 plus.n8 plus.n3 161.3
R16 plus.n11 plus.n2 161.3
R17 plus.n13 plus.n12 161.3
R18 plus.n14 plus.n1 161.3
R19 plus.n15 plus.n0 161.3
R20 plus.n17 plus.n16 161.3
R21 plus.n25 plus.n24 161.3
R22 plus.n26 plus.n21 161.3
R23 plus.n29 plus.n20 161.3
R24 plus.n31 plus.n30 161.3
R25 plus.n32 plus.n19 161.3
R26 plus.n33 plus.n18 161.3
R27 plus.n35 plus.n34 161.3
R28 plus.n10 plus.n9 80.6037
R29 plus.n28 plus.n27 80.6037
R30 plus.n9 plus.n2 48.2005
R31 plus.n9 plus.n8 48.2005
R32 plus.n27 plus.n20 48.2005
R33 plus.n27 plus.n26 48.2005
R34 plus.n14 plus.n13 45.2793
R35 plus.n7 plus.n4 45.2793
R36 plus.n32 plus.n31 45.2793
R37 plus.n25 plus.n22 45.2793
R38 plus.n24 plus.n23 44.9119
R39 plus.n6 plus.n5 44.9119
R40 plus plus.n35 36.3494
R41 plus.n16 plus.n15 35.055
R42 plus.n34 plus.n33 35.055
R43 plus.n23 plus.n22 17.739
R44 plus.n5 plus.n4 17.739
R45 plus plus.n17 17.1425
R46 plus.n15 plus.n14 13.146
R47 plus.n33 plus.n32 13.146
R48 plus.n13 plus.n2 2.92171
R49 plus.n8 plus.n7 2.92171
R50 plus.n31 plus.n20 2.92171
R51 plus.n26 plus.n25 2.92171
R52 plus.n10 plus.n3 0.285035
R53 plus.n11 plus.n10 0.285035
R54 plus.n29 plus.n28 0.285035
R55 plus.n28 plus.n21 0.285035
R56 plus.n6 plus.n3 0.189894
R57 plus.n12 plus.n11 0.189894
R58 plus.n12 plus.n1 0.189894
R59 plus.n1 plus.n0 0.189894
R60 plus.n17 plus.n0 0.189894
R61 plus.n35 plus.n18 0.189894
R62 plus.n19 plus.n18 0.189894
R63 plus.n30 plus.n19 0.189894
R64 plus.n30 plus.n29 0.189894
R65 plus.n24 plus.n21 0.189894
R66 drain_left.n134 drain_left.n0 289.615
R67 drain_left.n279 drain_left.n145 289.615
R68 drain_left.n44 drain_left.n43 185
R69 drain_left.n49 drain_left.n48 185
R70 drain_left.n51 drain_left.n50 185
R71 drain_left.n40 drain_left.n39 185
R72 drain_left.n57 drain_left.n56 185
R73 drain_left.n59 drain_left.n58 185
R74 drain_left.n36 drain_left.n35 185
R75 drain_left.n66 drain_left.n65 185
R76 drain_left.n67 drain_left.n34 185
R77 drain_left.n69 drain_left.n68 185
R78 drain_left.n32 drain_left.n31 185
R79 drain_left.n75 drain_left.n74 185
R80 drain_left.n77 drain_left.n76 185
R81 drain_left.n28 drain_left.n27 185
R82 drain_left.n83 drain_left.n82 185
R83 drain_left.n85 drain_left.n84 185
R84 drain_left.n24 drain_left.n23 185
R85 drain_left.n91 drain_left.n90 185
R86 drain_left.n93 drain_left.n92 185
R87 drain_left.n20 drain_left.n19 185
R88 drain_left.n99 drain_left.n98 185
R89 drain_left.n101 drain_left.n100 185
R90 drain_left.n16 drain_left.n15 185
R91 drain_left.n107 drain_left.n106 185
R92 drain_left.n110 drain_left.n109 185
R93 drain_left.n108 drain_left.n12 185
R94 drain_left.n115 drain_left.n11 185
R95 drain_left.n117 drain_left.n116 185
R96 drain_left.n119 drain_left.n118 185
R97 drain_left.n8 drain_left.n7 185
R98 drain_left.n125 drain_left.n124 185
R99 drain_left.n127 drain_left.n126 185
R100 drain_left.n4 drain_left.n3 185
R101 drain_left.n133 drain_left.n132 185
R102 drain_left.n135 drain_left.n134 185
R103 drain_left.n280 drain_left.n279 185
R104 drain_left.n278 drain_left.n277 185
R105 drain_left.n149 drain_left.n148 185
R106 drain_left.n272 drain_left.n271 185
R107 drain_left.n270 drain_left.n269 185
R108 drain_left.n153 drain_left.n152 185
R109 drain_left.n264 drain_left.n263 185
R110 drain_left.n262 drain_left.n261 185
R111 drain_left.n260 drain_left.n156 185
R112 drain_left.n160 drain_left.n157 185
R113 drain_left.n255 drain_left.n254 185
R114 drain_left.n253 drain_left.n252 185
R115 drain_left.n162 drain_left.n161 185
R116 drain_left.n247 drain_left.n246 185
R117 drain_left.n245 drain_left.n244 185
R118 drain_left.n166 drain_left.n165 185
R119 drain_left.n239 drain_left.n238 185
R120 drain_left.n237 drain_left.n236 185
R121 drain_left.n170 drain_left.n169 185
R122 drain_left.n231 drain_left.n230 185
R123 drain_left.n229 drain_left.n228 185
R124 drain_left.n174 drain_left.n173 185
R125 drain_left.n223 drain_left.n222 185
R126 drain_left.n221 drain_left.n220 185
R127 drain_left.n178 drain_left.n177 185
R128 drain_left.n215 drain_left.n214 185
R129 drain_left.n213 drain_left.n180 185
R130 drain_left.n212 drain_left.n211 185
R131 drain_left.n183 drain_left.n181 185
R132 drain_left.n206 drain_left.n205 185
R133 drain_left.n204 drain_left.n203 185
R134 drain_left.n187 drain_left.n186 185
R135 drain_left.n198 drain_left.n197 185
R136 drain_left.n196 drain_left.n195 185
R137 drain_left.n191 drain_left.n190 185
R138 drain_left.n45 drain_left.t11 149.524
R139 drain_left.n192 drain_left.t13 149.524
R140 drain_left.n49 drain_left.n43 104.615
R141 drain_left.n50 drain_left.n49 104.615
R142 drain_left.n50 drain_left.n39 104.615
R143 drain_left.n57 drain_left.n39 104.615
R144 drain_left.n58 drain_left.n57 104.615
R145 drain_left.n58 drain_left.n35 104.615
R146 drain_left.n66 drain_left.n35 104.615
R147 drain_left.n67 drain_left.n66 104.615
R148 drain_left.n68 drain_left.n67 104.615
R149 drain_left.n68 drain_left.n31 104.615
R150 drain_left.n75 drain_left.n31 104.615
R151 drain_left.n76 drain_left.n75 104.615
R152 drain_left.n76 drain_left.n27 104.615
R153 drain_left.n83 drain_left.n27 104.615
R154 drain_left.n84 drain_left.n83 104.615
R155 drain_left.n84 drain_left.n23 104.615
R156 drain_left.n91 drain_left.n23 104.615
R157 drain_left.n92 drain_left.n91 104.615
R158 drain_left.n92 drain_left.n19 104.615
R159 drain_left.n99 drain_left.n19 104.615
R160 drain_left.n100 drain_left.n99 104.615
R161 drain_left.n100 drain_left.n15 104.615
R162 drain_left.n107 drain_left.n15 104.615
R163 drain_left.n109 drain_left.n107 104.615
R164 drain_left.n109 drain_left.n108 104.615
R165 drain_left.n108 drain_left.n11 104.615
R166 drain_left.n117 drain_left.n11 104.615
R167 drain_left.n118 drain_left.n117 104.615
R168 drain_left.n118 drain_left.n7 104.615
R169 drain_left.n125 drain_left.n7 104.615
R170 drain_left.n126 drain_left.n125 104.615
R171 drain_left.n126 drain_left.n3 104.615
R172 drain_left.n133 drain_left.n3 104.615
R173 drain_left.n134 drain_left.n133 104.615
R174 drain_left.n279 drain_left.n278 104.615
R175 drain_left.n278 drain_left.n148 104.615
R176 drain_left.n271 drain_left.n148 104.615
R177 drain_left.n271 drain_left.n270 104.615
R178 drain_left.n270 drain_left.n152 104.615
R179 drain_left.n263 drain_left.n152 104.615
R180 drain_left.n263 drain_left.n262 104.615
R181 drain_left.n262 drain_left.n156 104.615
R182 drain_left.n160 drain_left.n156 104.615
R183 drain_left.n254 drain_left.n160 104.615
R184 drain_left.n254 drain_left.n253 104.615
R185 drain_left.n253 drain_left.n161 104.615
R186 drain_left.n246 drain_left.n161 104.615
R187 drain_left.n246 drain_left.n245 104.615
R188 drain_left.n245 drain_left.n165 104.615
R189 drain_left.n238 drain_left.n165 104.615
R190 drain_left.n238 drain_left.n237 104.615
R191 drain_left.n237 drain_left.n169 104.615
R192 drain_left.n230 drain_left.n169 104.615
R193 drain_left.n230 drain_left.n229 104.615
R194 drain_left.n229 drain_left.n173 104.615
R195 drain_left.n222 drain_left.n173 104.615
R196 drain_left.n222 drain_left.n221 104.615
R197 drain_left.n221 drain_left.n177 104.615
R198 drain_left.n214 drain_left.n177 104.615
R199 drain_left.n214 drain_left.n213 104.615
R200 drain_left.n213 drain_left.n212 104.615
R201 drain_left.n212 drain_left.n181 104.615
R202 drain_left.n205 drain_left.n181 104.615
R203 drain_left.n205 drain_left.n204 104.615
R204 drain_left.n204 drain_left.n186 104.615
R205 drain_left.n197 drain_left.n186 104.615
R206 drain_left.n197 drain_left.n196 104.615
R207 drain_left.n196 drain_left.n190 104.615
R208 drain_left.n143 drain_left.n141 59.5172
R209 drain_left.n143 drain_left.n142 58.7154
R210 drain_left.n140 drain_left.n139 58.7154
R211 drain_left.n287 drain_left.n286 58.7154
R212 drain_left.n285 drain_left.n284 58.7154
R213 drain_left.n289 drain_left.n288 58.7153
R214 drain_left.t11 drain_left.n43 52.3082
R215 drain_left.t13 drain_left.n190 52.3082
R216 drain_left.n140 drain_left.n138 48.1143
R217 drain_left.n285 drain_left.n283 48.1143
R218 drain_left drain_left.n144 41.8255
R219 drain_left.n69 drain_left.n34 13.1884
R220 drain_left.n116 drain_left.n115 13.1884
R221 drain_left.n261 drain_left.n260 13.1884
R222 drain_left.n215 drain_left.n180 13.1884
R223 drain_left.n65 drain_left.n64 12.8005
R224 drain_left.n70 drain_left.n32 12.8005
R225 drain_left.n114 drain_left.n12 12.8005
R226 drain_left.n119 drain_left.n10 12.8005
R227 drain_left.n264 drain_left.n155 12.8005
R228 drain_left.n259 drain_left.n157 12.8005
R229 drain_left.n216 drain_left.n178 12.8005
R230 drain_left.n211 drain_left.n182 12.8005
R231 drain_left.n63 drain_left.n36 12.0247
R232 drain_left.n74 drain_left.n73 12.0247
R233 drain_left.n111 drain_left.n110 12.0247
R234 drain_left.n120 drain_left.n8 12.0247
R235 drain_left.n265 drain_left.n153 12.0247
R236 drain_left.n256 drain_left.n255 12.0247
R237 drain_left.n220 drain_left.n219 12.0247
R238 drain_left.n210 drain_left.n183 12.0247
R239 drain_left.n60 drain_left.n59 11.249
R240 drain_left.n77 drain_left.n30 11.249
R241 drain_left.n106 drain_left.n14 11.249
R242 drain_left.n124 drain_left.n123 11.249
R243 drain_left.n269 drain_left.n268 11.249
R244 drain_left.n252 drain_left.n159 11.249
R245 drain_left.n223 drain_left.n176 11.249
R246 drain_left.n207 drain_left.n206 11.249
R247 drain_left.n56 drain_left.n38 10.4732
R248 drain_left.n78 drain_left.n28 10.4732
R249 drain_left.n105 drain_left.n16 10.4732
R250 drain_left.n127 drain_left.n6 10.4732
R251 drain_left.n272 drain_left.n151 10.4732
R252 drain_left.n251 drain_left.n162 10.4732
R253 drain_left.n224 drain_left.n174 10.4732
R254 drain_left.n203 drain_left.n185 10.4732
R255 drain_left.n45 drain_left.n44 10.2747
R256 drain_left.n192 drain_left.n191 10.2747
R257 drain_left.n55 drain_left.n40 9.69747
R258 drain_left.n82 drain_left.n81 9.69747
R259 drain_left.n102 drain_left.n101 9.69747
R260 drain_left.n128 drain_left.n4 9.69747
R261 drain_left.n273 drain_left.n149 9.69747
R262 drain_left.n248 drain_left.n247 9.69747
R263 drain_left.n228 drain_left.n227 9.69747
R264 drain_left.n202 drain_left.n187 9.69747
R265 drain_left.n138 drain_left.n137 9.45567
R266 drain_left.n283 drain_left.n282 9.45567
R267 drain_left.n2 drain_left.n1 9.3005
R268 drain_left.n131 drain_left.n130 9.3005
R269 drain_left.n129 drain_left.n128 9.3005
R270 drain_left.n6 drain_left.n5 9.3005
R271 drain_left.n123 drain_left.n122 9.3005
R272 drain_left.n121 drain_left.n120 9.3005
R273 drain_left.n10 drain_left.n9 9.3005
R274 drain_left.n89 drain_left.n88 9.3005
R275 drain_left.n87 drain_left.n86 9.3005
R276 drain_left.n26 drain_left.n25 9.3005
R277 drain_left.n81 drain_left.n80 9.3005
R278 drain_left.n79 drain_left.n78 9.3005
R279 drain_left.n30 drain_left.n29 9.3005
R280 drain_left.n73 drain_left.n72 9.3005
R281 drain_left.n71 drain_left.n70 9.3005
R282 drain_left.n47 drain_left.n46 9.3005
R283 drain_left.n42 drain_left.n41 9.3005
R284 drain_left.n53 drain_left.n52 9.3005
R285 drain_left.n55 drain_left.n54 9.3005
R286 drain_left.n38 drain_left.n37 9.3005
R287 drain_left.n61 drain_left.n60 9.3005
R288 drain_left.n63 drain_left.n62 9.3005
R289 drain_left.n64 drain_left.n33 9.3005
R290 drain_left.n22 drain_left.n21 9.3005
R291 drain_left.n95 drain_left.n94 9.3005
R292 drain_left.n97 drain_left.n96 9.3005
R293 drain_left.n18 drain_left.n17 9.3005
R294 drain_left.n103 drain_left.n102 9.3005
R295 drain_left.n105 drain_left.n104 9.3005
R296 drain_left.n14 drain_left.n13 9.3005
R297 drain_left.n112 drain_left.n111 9.3005
R298 drain_left.n114 drain_left.n113 9.3005
R299 drain_left.n137 drain_left.n136 9.3005
R300 drain_left.n194 drain_left.n193 9.3005
R301 drain_left.n189 drain_left.n188 9.3005
R302 drain_left.n200 drain_left.n199 9.3005
R303 drain_left.n202 drain_left.n201 9.3005
R304 drain_left.n185 drain_left.n184 9.3005
R305 drain_left.n208 drain_left.n207 9.3005
R306 drain_left.n210 drain_left.n209 9.3005
R307 drain_left.n182 drain_left.n179 9.3005
R308 drain_left.n241 drain_left.n240 9.3005
R309 drain_left.n243 drain_left.n242 9.3005
R310 drain_left.n164 drain_left.n163 9.3005
R311 drain_left.n249 drain_left.n248 9.3005
R312 drain_left.n251 drain_left.n250 9.3005
R313 drain_left.n159 drain_left.n158 9.3005
R314 drain_left.n257 drain_left.n256 9.3005
R315 drain_left.n259 drain_left.n258 9.3005
R316 drain_left.n282 drain_left.n281 9.3005
R317 drain_left.n147 drain_left.n146 9.3005
R318 drain_left.n276 drain_left.n275 9.3005
R319 drain_left.n274 drain_left.n273 9.3005
R320 drain_left.n151 drain_left.n150 9.3005
R321 drain_left.n268 drain_left.n267 9.3005
R322 drain_left.n266 drain_left.n265 9.3005
R323 drain_left.n155 drain_left.n154 9.3005
R324 drain_left.n168 drain_left.n167 9.3005
R325 drain_left.n235 drain_left.n234 9.3005
R326 drain_left.n233 drain_left.n232 9.3005
R327 drain_left.n172 drain_left.n171 9.3005
R328 drain_left.n227 drain_left.n226 9.3005
R329 drain_left.n225 drain_left.n224 9.3005
R330 drain_left.n176 drain_left.n175 9.3005
R331 drain_left.n219 drain_left.n218 9.3005
R332 drain_left.n217 drain_left.n216 9.3005
R333 drain_left.n52 drain_left.n51 8.92171
R334 drain_left.n85 drain_left.n26 8.92171
R335 drain_left.n98 drain_left.n18 8.92171
R336 drain_left.n132 drain_left.n131 8.92171
R337 drain_left.n277 drain_left.n276 8.92171
R338 drain_left.n244 drain_left.n164 8.92171
R339 drain_left.n231 drain_left.n172 8.92171
R340 drain_left.n199 drain_left.n198 8.92171
R341 drain_left.n48 drain_left.n42 8.14595
R342 drain_left.n86 drain_left.n24 8.14595
R343 drain_left.n97 drain_left.n20 8.14595
R344 drain_left.n135 drain_left.n2 8.14595
R345 drain_left.n280 drain_left.n147 8.14595
R346 drain_left.n243 drain_left.n166 8.14595
R347 drain_left.n232 drain_left.n170 8.14595
R348 drain_left.n195 drain_left.n189 8.14595
R349 drain_left.n47 drain_left.n44 7.3702
R350 drain_left.n90 drain_left.n89 7.3702
R351 drain_left.n94 drain_left.n93 7.3702
R352 drain_left.n136 drain_left.n0 7.3702
R353 drain_left.n281 drain_left.n145 7.3702
R354 drain_left.n240 drain_left.n239 7.3702
R355 drain_left.n236 drain_left.n235 7.3702
R356 drain_left.n194 drain_left.n191 7.3702
R357 drain_left.n90 drain_left.n22 6.59444
R358 drain_left.n93 drain_left.n22 6.59444
R359 drain_left.n138 drain_left.n0 6.59444
R360 drain_left.n283 drain_left.n145 6.59444
R361 drain_left.n239 drain_left.n168 6.59444
R362 drain_left.n236 drain_left.n168 6.59444
R363 drain_left drain_left.n289 6.45494
R364 drain_left.n48 drain_left.n47 5.81868
R365 drain_left.n89 drain_left.n24 5.81868
R366 drain_left.n94 drain_left.n20 5.81868
R367 drain_left.n136 drain_left.n135 5.81868
R368 drain_left.n281 drain_left.n280 5.81868
R369 drain_left.n240 drain_left.n166 5.81868
R370 drain_left.n235 drain_left.n170 5.81868
R371 drain_left.n195 drain_left.n194 5.81868
R372 drain_left.n51 drain_left.n42 5.04292
R373 drain_left.n86 drain_left.n85 5.04292
R374 drain_left.n98 drain_left.n97 5.04292
R375 drain_left.n132 drain_left.n2 5.04292
R376 drain_left.n277 drain_left.n147 5.04292
R377 drain_left.n244 drain_left.n243 5.04292
R378 drain_left.n232 drain_left.n231 5.04292
R379 drain_left.n198 drain_left.n189 5.04292
R380 drain_left.n52 drain_left.n40 4.26717
R381 drain_left.n82 drain_left.n26 4.26717
R382 drain_left.n101 drain_left.n18 4.26717
R383 drain_left.n131 drain_left.n4 4.26717
R384 drain_left.n276 drain_left.n149 4.26717
R385 drain_left.n247 drain_left.n164 4.26717
R386 drain_left.n228 drain_left.n172 4.26717
R387 drain_left.n199 drain_left.n187 4.26717
R388 drain_left.n56 drain_left.n55 3.49141
R389 drain_left.n81 drain_left.n28 3.49141
R390 drain_left.n102 drain_left.n16 3.49141
R391 drain_left.n128 drain_left.n127 3.49141
R392 drain_left.n273 drain_left.n272 3.49141
R393 drain_left.n248 drain_left.n162 3.49141
R394 drain_left.n227 drain_left.n174 3.49141
R395 drain_left.n203 drain_left.n202 3.49141
R396 drain_left.n193 drain_left.n192 2.84303
R397 drain_left.n46 drain_left.n45 2.84303
R398 drain_left.n59 drain_left.n38 2.71565
R399 drain_left.n78 drain_left.n77 2.71565
R400 drain_left.n106 drain_left.n105 2.71565
R401 drain_left.n124 drain_left.n6 2.71565
R402 drain_left.n269 drain_left.n151 2.71565
R403 drain_left.n252 drain_left.n251 2.71565
R404 drain_left.n224 drain_left.n223 2.71565
R405 drain_left.n206 drain_left.n185 2.71565
R406 drain_left.n60 drain_left.n36 1.93989
R407 drain_left.n74 drain_left.n30 1.93989
R408 drain_left.n110 drain_left.n14 1.93989
R409 drain_left.n123 drain_left.n8 1.93989
R410 drain_left.n268 drain_left.n153 1.93989
R411 drain_left.n255 drain_left.n159 1.93989
R412 drain_left.n220 drain_left.n176 1.93989
R413 drain_left.n207 drain_left.n183 1.93989
R414 drain_left.n65 drain_left.n63 1.16414
R415 drain_left.n73 drain_left.n32 1.16414
R416 drain_left.n111 drain_left.n12 1.16414
R417 drain_left.n120 drain_left.n119 1.16414
R418 drain_left.n265 drain_left.n264 1.16414
R419 drain_left.n256 drain_left.n157 1.16414
R420 drain_left.n219 drain_left.n178 1.16414
R421 drain_left.n211 drain_left.n210 1.16414
R422 drain_left.n287 drain_left.n285 0.802224
R423 drain_left.n289 drain_left.n287 0.802224
R424 drain_left.n141 drain_left.t7 0.7925
R425 drain_left.n141 drain_left.t10 0.7925
R426 drain_left.n142 drain_left.t5 0.7925
R427 drain_left.n142 drain_left.t12 0.7925
R428 drain_left.n139 drain_left.t3 0.7925
R429 drain_left.n139 drain_left.t0 0.7925
R430 drain_left.n288 drain_left.t1 0.7925
R431 drain_left.n288 drain_left.t4 0.7925
R432 drain_left.n286 drain_left.t6 0.7925
R433 drain_left.n286 drain_left.t2 0.7925
R434 drain_left.n284 drain_left.t8 0.7925
R435 drain_left.n284 drain_left.t9 0.7925
R436 drain_left.n144 drain_left.n140 0.546447
R437 drain_left.n64 drain_left.n34 0.388379
R438 drain_left.n70 drain_left.n69 0.388379
R439 drain_left.n115 drain_left.n114 0.388379
R440 drain_left.n116 drain_left.n10 0.388379
R441 drain_left.n261 drain_left.n155 0.388379
R442 drain_left.n260 drain_left.n259 0.388379
R443 drain_left.n216 drain_left.n215 0.388379
R444 drain_left.n182 drain_left.n180 0.388379
R445 drain_left.n46 drain_left.n41 0.155672
R446 drain_left.n53 drain_left.n41 0.155672
R447 drain_left.n54 drain_left.n53 0.155672
R448 drain_left.n54 drain_left.n37 0.155672
R449 drain_left.n61 drain_left.n37 0.155672
R450 drain_left.n62 drain_left.n61 0.155672
R451 drain_left.n62 drain_left.n33 0.155672
R452 drain_left.n71 drain_left.n33 0.155672
R453 drain_left.n72 drain_left.n71 0.155672
R454 drain_left.n72 drain_left.n29 0.155672
R455 drain_left.n79 drain_left.n29 0.155672
R456 drain_left.n80 drain_left.n79 0.155672
R457 drain_left.n80 drain_left.n25 0.155672
R458 drain_left.n87 drain_left.n25 0.155672
R459 drain_left.n88 drain_left.n87 0.155672
R460 drain_left.n88 drain_left.n21 0.155672
R461 drain_left.n95 drain_left.n21 0.155672
R462 drain_left.n96 drain_left.n95 0.155672
R463 drain_left.n96 drain_left.n17 0.155672
R464 drain_left.n103 drain_left.n17 0.155672
R465 drain_left.n104 drain_left.n103 0.155672
R466 drain_left.n104 drain_left.n13 0.155672
R467 drain_left.n112 drain_left.n13 0.155672
R468 drain_left.n113 drain_left.n112 0.155672
R469 drain_left.n113 drain_left.n9 0.155672
R470 drain_left.n121 drain_left.n9 0.155672
R471 drain_left.n122 drain_left.n121 0.155672
R472 drain_left.n122 drain_left.n5 0.155672
R473 drain_left.n129 drain_left.n5 0.155672
R474 drain_left.n130 drain_left.n129 0.155672
R475 drain_left.n130 drain_left.n1 0.155672
R476 drain_left.n137 drain_left.n1 0.155672
R477 drain_left.n282 drain_left.n146 0.155672
R478 drain_left.n275 drain_left.n146 0.155672
R479 drain_left.n275 drain_left.n274 0.155672
R480 drain_left.n274 drain_left.n150 0.155672
R481 drain_left.n267 drain_left.n150 0.155672
R482 drain_left.n267 drain_left.n266 0.155672
R483 drain_left.n266 drain_left.n154 0.155672
R484 drain_left.n258 drain_left.n154 0.155672
R485 drain_left.n258 drain_left.n257 0.155672
R486 drain_left.n257 drain_left.n158 0.155672
R487 drain_left.n250 drain_left.n158 0.155672
R488 drain_left.n250 drain_left.n249 0.155672
R489 drain_left.n249 drain_left.n163 0.155672
R490 drain_left.n242 drain_left.n163 0.155672
R491 drain_left.n242 drain_left.n241 0.155672
R492 drain_left.n241 drain_left.n167 0.155672
R493 drain_left.n234 drain_left.n167 0.155672
R494 drain_left.n234 drain_left.n233 0.155672
R495 drain_left.n233 drain_left.n171 0.155672
R496 drain_left.n226 drain_left.n171 0.155672
R497 drain_left.n226 drain_left.n225 0.155672
R498 drain_left.n225 drain_left.n175 0.155672
R499 drain_left.n218 drain_left.n175 0.155672
R500 drain_left.n218 drain_left.n217 0.155672
R501 drain_left.n217 drain_left.n179 0.155672
R502 drain_left.n209 drain_left.n179 0.155672
R503 drain_left.n209 drain_left.n208 0.155672
R504 drain_left.n208 drain_left.n184 0.155672
R505 drain_left.n201 drain_left.n184 0.155672
R506 drain_left.n201 drain_left.n200 0.155672
R507 drain_left.n200 drain_left.n188 0.155672
R508 drain_left.n193 drain_left.n188 0.155672
R509 drain_left.n144 drain_left.n143 0.145585
R510 source.n578 source.n444 289.615
R511 source.n432 source.n298 289.615
R512 source.n134 source.n0 289.615
R513 source.n280 source.n146 289.615
R514 source.n488 source.n487 185
R515 source.n493 source.n492 185
R516 source.n495 source.n494 185
R517 source.n484 source.n483 185
R518 source.n501 source.n500 185
R519 source.n503 source.n502 185
R520 source.n480 source.n479 185
R521 source.n510 source.n509 185
R522 source.n511 source.n478 185
R523 source.n513 source.n512 185
R524 source.n476 source.n475 185
R525 source.n519 source.n518 185
R526 source.n521 source.n520 185
R527 source.n472 source.n471 185
R528 source.n527 source.n526 185
R529 source.n529 source.n528 185
R530 source.n468 source.n467 185
R531 source.n535 source.n534 185
R532 source.n537 source.n536 185
R533 source.n464 source.n463 185
R534 source.n543 source.n542 185
R535 source.n545 source.n544 185
R536 source.n460 source.n459 185
R537 source.n551 source.n550 185
R538 source.n554 source.n553 185
R539 source.n552 source.n456 185
R540 source.n559 source.n455 185
R541 source.n561 source.n560 185
R542 source.n563 source.n562 185
R543 source.n452 source.n451 185
R544 source.n569 source.n568 185
R545 source.n571 source.n570 185
R546 source.n448 source.n447 185
R547 source.n577 source.n576 185
R548 source.n579 source.n578 185
R549 source.n342 source.n341 185
R550 source.n347 source.n346 185
R551 source.n349 source.n348 185
R552 source.n338 source.n337 185
R553 source.n355 source.n354 185
R554 source.n357 source.n356 185
R555 source.n334 source.n333 185
R556 source.n364 source.n363 185
R557 source.n365 source.n332 185
R558 source.n367 source.n366 185
R559 source.n330 source.n329 185
R560 source.n373 source.n372 185
R561 source.n375 source.n374 185
R562 source.n326 source.n325 185
R563 source.n381 source.n380 185
R564 source.n383 source.n382 185
R565 source.n322 source.n321 185
R566 source.n389 source.n388 185
R567 source.n391 source.n390 185
R568 source.n318 source.n317 185
R569 source.n397 source.n396 185
R570 source.n399 source.n398 185
R571 source.n314 source.n313 185
R572 source.n405 source.n404 185
R573 source.n408 source.n407 185
R574 source.n406 source.n310 185
R575 source.n413 source.n309 185
R576 source.n415 source.n414 185
R577 source.n417 source.n416 185
R578 source.n306 source.n305 185
R579 source.n423 source.n422 185
R580 source.n425 source.n424 185
R581 source.n302 source.n301 185
R582 source.n431 source.n430 185
R583 source.n433 source.n432 185
R584 source.n135 source.n134 185
R585 source.n133 source.n132 185
R586 source.n4 source.n3 185
R587 source.n127 source.n126 185
R588 source.n125 source.n124 185
R589 source.n8 source.n7 185
R590 source.n119 source.n118 185
R591 source.n117 source.n116 185
R592 source.n115 source.n11 185
R593 source.n15 source.n12 185
R594 source.n110 source.n109 185
R595 source.n108 source.n107 185
R596 source.n17 source.n16 185
R597 source.n102 source.n101 185
R598 source.n100 source.n99 185
R599 source.n21 source.n20 185
R600 source.n94 source.n93 185
R601 source.n92 source.n91 185
R602 source.n25 source.n24 185
R603 source.n86 source.n85 185
R604 source.n84 source.n83 185
R605 source.n29 source.n28 185
R606 source.n78 source.n77 185
R607 source.n76 source.n75 185
R608 source.n33 source.n32 185
R609 source.n70 source.n69 185
R610 source.n68 source.n35 185
R611 source.n67 source.n66 185
R612 source.n38 source.n36 185
R613 source.n61 source.n60 185
R614 source.n59 source.n58 185
R615 source.n42 source.n41 185
R616 source.n53 source.n52 185
R617 source.n51 source.n50 185
R618 source.n46 source.n45 185
R619 source.n281 source.n280 185
R620 source.n279 source.n278 185
R621 source.n150 source.n149 185
R622 source.n273 source.n272 185
R623 source.n271 source.n270 185
R624 source.n154 source.n153 185
R625 source.n265 source.n264 185
R626 source.n263 source.n262 185
R627 source.n261 source.n157 185
R628 source.n161 source.n158 185
R629 source.n256 source.n255 185
R630 source.n254 source.n253 185
R631 source.n163 source.n162 185
R632 source.n248 source.n247 185
R633 source.n246 source.n245 185
R634 source.n167 source.n166 185
R635 source.n240 source.n239 185
R636 source.n238 source.n237 185
R637 source.n171 source.n170 185
R638 source.n232 source.n231 185
R639 source.n230 source.n229 185
R640 source.n175 source.n174 185
R641 source.n224 source.n223 185
R642 source.n222 source.n221 185
R643 source.n179 source.n178 185
R644 source.n216 source.n215 185
R645 source.n214 source.n181 185
R646 source.n213 source.n212 185
R647 source.n184 source.n182 185
R648 source.n207 source.n206 185
R649 source.n205 source.n204 185
R650 source.n188 source.n187 185
R651 source.n199 source.n198 185
R652 source.n197 source.n196 185
R653 source.n192 source.n191 185
R654 source.n489 source.t6 149.524
R655 source.n343 source.t14 149.524
R656 source.n47 source.t26 149.524
R657 source.n193 source.t7 149.524
R658 source.n493 source.n487 104.615
R659 source.n494 source.n493 104.615
R660 source.n494 source.n483 104.615
R661 source.n501 source.n483 104.615
R662 source.n502 source.n501 104.615
R663 source.n502 source.n479 104.615
R664 source.n510 source.n479 104.615
R665 source.n511 source.n510 104.615
R666 source.n512 source.n511 104.615
R667 source.n512 source.n475 104.615
R668 source.n519 source.n475 104.615
R669 source.n520 source.n519 104.615
R670 source.n520 source.n471 104.615
R671 source.n527 source.n471 104.615
R672 source.n528 source.n527 104.615
R673 source.n528 source.n467 104.615
R674 source.n535 source.n467 104.615
R675 source.n536 source.n535 104.615
R676 source.n536 source.n463 104.615
R677 source.n543 source.n463 104.615
R678 source.n544 source.n543 104.615
R679 source.n544 source.n459 104.615
R680 source.n551 source.n459 104.615
R681 source.n553 source.n551 104.615
R682 source.n553 source.n552 104.615
R683 source.n552 source.n455 104.615
R684 source.n561 source.n455 104.615
R685 source.n562 source.n561 104.615
R686 source.n562 source.n451 104.615
R687 source.n569 source.n451 104.615
R688 source.n570 source.n569 104.615
R689 source.n570 source.n447 104.615
R690 source.n577 source.n447 104.615
R691 source.n578 source.n577 104.615
R692 source.n347 source.n341 104.615
R693 source.n348 source.n347 104.615
R694 source.n348 source.n337 104.615
R695 source.n355 source.n337 104.615
R696 source.n356 source.n355 104.615
R697 source.n356 source.n333 104.615
R698 source.n364 source.n333 104.615
R699 source.n365 source.n364 104.615
R700 source.n366 source.n365 104.615
R701 source.n366 source.n329 104.615
R702 source.n373 source.n329 104.615
R703 source.n374 source.n373 104.615
R704 source.n374 source.n325 104.615
R705 source.n381 source.n325 104.615
R706 source.n382 source.n381 104.615
R707 source.n382 source.n321 104.615
R708 source.n389 source.n321 104.615
R709 source.n390 source.n389 104.615
R710 source.n390 source.n317 104.615
R711 source.n397 source.n317 104.615
R712 source.n398 source.n397 104.615
R713 source.n398 source.n313 104.615
R714 source.n405 source.n313 104.615
R715 source.n407 source.n405 104.615
R716 source.n407 source.n406 104.615
R717 source.n406 source.n309 104.615
R718 source.n415 source.n309 104.615
R719 source.n416 source.n415 104.615
R720 source.n416 source.n305 104.615
R721 source.n423 source.n305 104.615
R722 source.n424 source.n423 104.615
R723 source.n424 source.n301 104.615
R724 source.n431 source.n301 104.615
R725 source.n432 source.n431 104.615
R726 source.n134 source.n133 104.615
R727 source.n133 source.n3 104.615
R728 source.n126 source.n3 104.615
R729 source.n126 source.n125 104.615
R730 source.n125 source.n7 104.615
R731 source.n118 source.n7 104.615
R732 source.n118 source.n117 104.615
R733 source.n117 source.n11 104.615
R734 source.n15 source.n11 104.615
R735 source.n109 source.n15 104.615
R736 source.n109 source.n108 104.615
R737 source.n108 source.n16 104.615
R738 source.n101 source.n16 104.615
R739 source.n101 source.n100 104.615
R740 source.n100 source.n20 104.615
R741 source.n93 source.n20 104.615
R742 source.n93 source.n92 104.615
R743 source.n92 source.n24 104.615
R744 source.n85 source.n24 104.615
R745 source.n85 source.n84 104.615
R746 source.n84 source.n28 104.615
R747 source.n77 source.n28 104.615
R748 source.n77 source.n76 104.615
R749 source.n76 source.n32 104.615
R750 source.n69 source.n32 104.615
R751 source.n69 source.n68 104.615
R752 source.n68 source.n67 104.615
R753 source.n67 source.n36 104.615
R754 source.n60 source.n36 104.615
R755 source.n60 source.n59 104.615
R756 source.n59 source.n41 104.615
R757 source.n52 source.n41 104.615
R758 source.n52 source.n51 104.615
R759 source.n51 source.n45 104.615
R760 source.n280 source.n279 104.615
R761 source.n279 source.n149 104.615
R762 source.n272 source.n149 104.615
R763 source.n272 source.n271 104.615
R764 source.n271 source.n153 104.615
R765 source.n264 source.n153 104.615
R766 source.n264 source.n263 104.615
R767 source.n263 source.n157 104.615
R768 source.n161 source.n157 104.615
R769 source.n255 source.n161 104.615
R770 source.n255 source.n254 104.615
R771 source.n254 source.n162 104.615
R772 source.n247 source.n162 104.615
R773 source.n247 source.n246 104.615
R774 source.n246 source.n166 104.615
R775 source.n239 source.n166 104.615
R776 source.n239 source.n238 104.615
R777 source.n238 source.n170 104.615
R778 source.n231 source.n170 104.615
R779 source.n231 source.n230 104.615
R780 source.n230 source.n174 104.615
R781 source.n223 source.n174 104.615
R782 source.n223 source.n222 104.615
R783 source.n222 source.n178 104.615
R784 source.n215 source.n178 104.615
R785 source.n215 source.n214 104.615
R786 source.n214 source.n213 104.615
R787 source.n213 source.n182 104.615
R788 source.n206 source.n182 104.615
R789 source.n206 source.n205 104.615
R790 source.n205 source.n187 104.615
R791 source.n198 source.n187 104.615
R792 source.n198 source.n197 104.615
R793 source.n197 source.n191 104.615
R794 source.t6 source.n487 52.3082
R795 source.t14 source.n341 52.3082
R796 source.t26 source.n45 52.3082
R797 source.t7 source.n191 52.3082
R798 source.n443 source.n442 42.0366
R799 source.n441 source.n440 42.0366
R800 source.n439 source.n438 42.0366
R801 source.n297 source.n296 42.0366
R802 source.n295 source.n294 42.0366
R803 source.n293 source.n292 42.0366
R804 source.n141 source.n140 42.0366
R805 source.n143 source.n142 42.0366
R806 source.n145 source.n144 42.0366
R807 source.n287 source.n286 42.0366
R808 source.n289 source.n288 42.0366
R809 source.n291 source.n290 42.0366
R810 source.n293 source.n291 32.7397
R811 source.n583 source.n582 30.6338
R812 source.n437 source.n436 30.6338
R813 source.n139 source.n138 30.6338
R814 source.n285 source.n284 30.6338
R815 source.n584 source.n139 26.2741
R816 source.n513 source.n478 13.1884
R817 source.n560 source.n559 13.1884
R818 source.n367 source.n332 13.1884
R819 source.n414 source.n413 13.1884
R820 source.n116 source.n115 13.1884
R821 source.n70 source.n35 13.1884
R822 source.n262 source.n261 13.1884
R823 source.n216 source.n181 13.1884
R824 source.n509 source.n508 12.8005
R825 source.n514 source.n476 12.8005
R826 source.n558 source.n456 12.8005
R827 source.n563 source.n454 12.8005
R828 source.n363 source.n362 12.8005
R829 source.n368 source.n330 12.8005
R830 source.n412 source.n310 12.8005
R831 source.n417 source.n308 12.8005
R832 source.n119 source.n10 12.8005
R833 source.n114 source.n12 12.8005
R834 source.n71 source.n33 12.8005
R835 source.n66 source.n37 12.8005
R836 source.n265 source.n156 12.8005
R837 source.n260 source.n158 12.8005
R838 source.n217 source.n179 12.8005
R839 source.n212 source.n183 12.8005
R840 source.n507 source.n480 12.0247
R841 source.n518 source.n517 12.0247
R842 source.n555 source.n554 12.0247
R843 source.n564 source.n452 12.0247
R844 source.n361 source.n334 12.0247
R845 source.n372 source.n371 12.0247
R846 source.n409 source.n408 12.0247
R847 source.n418 source.n306 12.0247
R848 source.n120 source.n8 12.0247
R849 source.n111 source.n110 12.0247
R850 source.n75 source.n74 12.0247
R851 source.n65 source.n38 12.0247
R852 source.n266 source.n154 12.0247
R853 source.n257 source.n256 12.0247
R854 source.n221 source.n220 12.0247
R855 source.n211 source.n184 12.0247
R856 source.n504 source.n503 11.249
R857 source.n521 source.n474 11.249
R858 source.n550 source.n458 11.249
R859 source.n568 source.n567 11.249
R860 source.n358 source.n357 11.249
R861 source.n375 source.n328 11.249
R862 source.n404 source.n312 11.249
R863 source.n422 source.n421 11.249
R864 source.n124 source.n123 11.249
R865 source.n107 source.n14 11.249
R866 source.n78 source.n31 11.249
R867 source.n62 source.n61 11.249
R868 source.n270 source.n269 11.249
R869 source.n253 source.n160 11.249
R870 source.n224 source.n177 11.249
R871 source.n208 source.n207 11.249
R872 source.n500 source.n482 10.4732
R873 source.n522 source.n472 10.4732
R874 source.n549 source.n460 10.4732
R875 source.n571 source.n450 10.4732
R876 source.n354 source.n336 10.4732
R877 source.n376 source.n326 10.4732
R878 source.n403 source.n314 10.4732
R879 source.n425 source.n304 10.4732
R880 source.n127 source.n6 10.4732
R881 source.n106 source.n17 10.4732
R882 source.n79 source.n29 10.4732
R883 source.n58 source.n40 10.4732
R884 source.n273 source.n152 10.4732
R885 source.n252 source.n163 10.4732
R886 source.n225 source.n175 10.4732
R887 source.n204 source.n186 10.4732
R888 source.n489 source.n488 10.2747
R889 source.n343 source.n342 10.2747
R890 source.n47 source.n46 10.2747
R891 source.n193 source.n192 10.2747
R892 source.n499 source.n484 9.69747
R893 source.n526 source.n525 9.69747
R894 source.n546 source.n545 9.69747
R895 source.n572 source.n448 9.69747
R896 source.n353 source.n338 9.69747
R897 source.n380 source.n379 9.69747
R898 source.n400 source.n399 9.69747
R899 source.n426 source.n302 9.69747
R900 source.n128 source.n4 9.69747
R901 source.n103 source.n102 9.69747
R902 source.n83 source.n82 9.69747
R903 source.n57 source.n42 9.69747
R904 source.n274 source.n150 9.69747
R905 source.n249 source.n248 9.69747
R906 source.n229 source.n228 9.69747
R907 source.n203 source.n188 9.69747
R908 source.n582 source.n581 9.45567
R909 source.n436 source.n435 9.45567
R910 source.n138 source.n137 9.45567
R911 source.n284 source.n283 9.45567
R912 source.n446 source.n445 9.3005
R913 source.n575 source.n574 9.3005
R914 source.n573 source.n572 9.3005
R915 source.n450 source.n449 9.3005
R916 source.n567 source.n566 9.3005
R917 source.n565 source.n564 9.3005
R918 source.n454 source.n453 9.3005
R919 source.n533 source.n532 9.3005
R920 source.n531 source.n530 9.3005
R921 source.n470 source.n469 9.3005
R922 source.n525 source.n524 9.3005
R923 source.n523 source.n522 9.3005
R924 source.n474 source.n473 9.3005
R925 source.n517 source.n516 9.3005
R926 source.n515 source.n514 9.3005
R927 source.n491 source.n490 9.3005
R928 source.n486 source.n485 9.3005
R929 source.n497 source.n496 9.3005
R930 source.n499 source.n498 9.3005
R931 source.n482 source.n481 9.3005
R932 source.n505 source.n504 9.3005
R933 source.n507 source.n506 9.3005
R934 source.n508 source.n477 9.3005
R935 source.n466 source.n465 9.3005
R936 source.n539 source.n538 9.3005
R937 source.n541 source.n540 9.3005
R938 source.n462 source.n461 9.3005
R939 source.n547 source.n546 9.3005
R940 source.n549 source.n548 9.3005
R941 source.n458 source.n457 9.3005
R942 source.n556 source.n555 9.3005
R943 source.n558 source.n557 9.3005
R944 source.n581 source.n580 9.3005
R945 source.n300 source.n299 9.3005
R946 source.n429 source.n428 9.3005
R947 source.n427 source.n426 9.3005
R948 source.n304 source.n303 9.3005
R949 source.n421 source.n420 9.3005
R950 source.n419 source.n418 9.3005
R951 source.n308 source.n307 9.3005
R952 source.n387 source.n386 9.3005
R953 source.n385 source.n384 9.3005
R954 source.n324 source.n323 9.3005
R955 source.n379 source.n378 9.3005
R956 source.n377 source.n376 9.3005
R957 source.n328 source.n327 9.3005
R958 source.n371 source.n370 9.3005
R959 source.n369 source.n368 9.3005
R960 source.n345 source.n344 9.3005
R961 source.n340 source.n339 9.3005
R962 source.n351 source.n350 9.3005
R963 source.n353 source.n352 9.3005
R964 source.n336 source.n335 9.3005
R965 source.n359 source.n358 9.3005
R966 source.n361 source.n360 9.3005
R967 source.n362 source.n331 9.3005
R968 source.n320 source.n319 9.3005
R969 source.n393 source.n392 9.3005
R970 source.n395 source.n394 9.3005
R971 source.n316 source.n315 9.3005
R972 source.n401 source.n400 9.3005
R973 source.n403 source.n402 9.3005
R974 source.n312 source.n311 9.3005
R975 source.n410 source.n409 9.3005
R976 source.n412 source.n411 9.3005
R977 source.n435 source.n434 9.3005
R978 source.n49 source.n48 9.3005
R979 source.n44 source.n43 9.3005
R980 source.n55 source.n54 9.3005
R981 source.n57 source.n56 9.3005
R982 source.n40 source.n39 9.3005
R983 source.n63 source.n62 9.3005
R984 source.n65 source.n64 9.3005
R985 source.n37 source.n34 9.3005
R986 source.n96 source.n95 9.3005
R987 source.n98 source.n97 9.3005
R988 source.n19 source.n18 9.3005
R989 source.n104 source.n103 9.3005
R990 source.n106 source.n105 9.3005
R991 source.n14 source.n13 9.3005
R992 source.n112 source.n111 9.3005
R993 source.n114 source.n113 9.3005
R994 source.n137 source.n136 9.3005
R995 source.n2 source.n1 9.3005
R996 source.n131 source.n130 9.3005
R997 source.n129 source.n128 9.3005
R998 source.n6 source.n5 9.3005
R999 source.n123 source.n122 9.3005
R1000 source.n121 source.n120 9.3005
R1001 source.n10 source.n9 9.3005
R1002 source.n23 source.n22 9.3005
R1003 source.n90 source.n89 9.3005
R1004 source.n88 source.n87 9.3005
R1005 source.n27 source.n26 9.3005
R1006 source.n82 source.n81 9.3005
R1007 source.n80 source.n79 9.3005
R1008 source.n31 source.n30 9.3005
R1009 source.n74 source.n73 9.3005
R1010 source.n72 source.n71 9.3005
R1011 source.n195 source.n194 9.3005
R1012 source.n190 source.n189 9.3005
R1013 source.n201 source.n200 9.3005
R1014 source.n203 source.n202 9.3005
R1015 source.n186 source.n185 9.3005
R1016 source.n209 source.n208 9.3005
R1017 source.n211 source.n210 9.3005
R1018 source.n183 source.n180 9.3005
R1019 source.n242 source.n241 9.3005
R1020 source.n244 source.n243 9.3005
R1021 source.n165 source.n164 9.3005
R1022 source.n250 source.n249 9.3005
R1023 source.n252 source.n251 9.3005
R1024 source.n160 source.n159 9.3005
R1025 source.n258 source.n257 9.3005
R1026 source.n260 source.n259 9.3005
R1027 source.n283 source.n282 9.3005
R1028 source.n148 source.n147 9.3005
R1029 source.n277 source.n276 9.3005
R1030 source.n275 source.n274 9.3005
R1031 source.n152 source.n151 9.3005
R1032 source.n269 source.n268 9.3005
R1033 source.n267 source.n266 9.3005
R1034 source.n156 source.n155 9.3005
R1035 source.n169 source.n168 9.3005
R1036 source.n236 source.n235 9.3005
R1037 source.n234 source.n233 9.3005
R1038 source.n173 source.n172 9.3005
R1039 source.n228 source.n227 9.3005
R1040 source.n226 source.n225 9.3005
R1041 source.n177 source.n176 9.3005
R1042 source.n220 source.n219 9.3005
R1043 source.n218 source.n217 9.3005
R1044 source.n496 source.n495 8.92171
R1045 source.n529 source.n470 8.92171
R1046 source.n542 source.n462 8.92171
R1047 source.n576 source.n575 8.92171
R1048 source.n350 source.n349 8.92171
R1049 source.n383 source.n324 8.92171
R1050 source.n396 source.n316 8.92171
R1051 source.n430 source.n429 8.92171
R1052 source.n132 source.n131 8.92171
R1053 source.n99 source.n19 8.92171
R1054 source.n86 source.n27 8.92171
R1055 source.n54 source.n53 8.92171
R1056 source.n278 source.n277 8.92171
R1057 source.n245 source.n165 8.92171
R1058 source.n232 source.n173 8.92171
R1059 source.n200 source.n199 8.92171
R1060 source.n492 source.n486 8.14595
R1061 source.n530 source.n468 8.14595
R1062 source.n541 source.n464 8.14595
R1063 source.n579 source.n446 8.14595
R1064 source.n346 source.n340 8.14595
R1065 source.n384 source.n322 8.14595
R1066 source.n395 source.n318 8.14595
R1067 source.n433 source.n300 8.14595
R1068 source.n135 source.n2 8.14595
R1069 source.n98 source.n21 8.14595
R1070 source.n87 source.n25 8.14595
R1071 source.n50 source.n44 8.14595
R1072 source.n281 source.n148 8.14595
R1073 source.n244 source.n167 8.14595
R1074 source.n233 source.n171 8.14595
R1075 source.n196 source.n190 8.14595
R1076 source.n491 source.n488 7.3702
R1077 source.n534 source.n533 7.3702
R1078 source.n538 source.n537 7.3702
R1079 source.n580 source.n444 7.3702
R1080 source.n345 source.n342 7.3702
R1081 source.n388 source.n387 7.3702
R1082 source.n392 source.n391 7.3702
R1083 source.n434 source.n298 7.3702
R1084 source.n136 source.n0 7.3702
R1085 source.n95 source.n94 7.3702
R1086 source.n91 source.n90 7.3702
R1087 source.n49 source.n46 7.3702
R1088 source.n282 source.n146 7.3702
R1089 source.n241 source.n240 7.3702
R1090 source.n237 source.n236 7.3702
R1091 source.n195 source.n192 7.3702
R1092 source.n534 source.n466 6.59444
R1093 source.n537 source.n466 6.59444
R1094 source.n582 source.n444 6.59444
R1095 source.n388 source.n320 6.59444
R1096 source.n391 source.n320 6.59444
R1097 source.n436 source.n298 6.59444
R1098 source.n138 source.n0 6.59444
R1099 source.n94 source.n23 6.59444
R1100 source.n91 source.n23 6.59444
R1101 source.n284 source.n146 6.59444
R1102 source.n240 source.n169 6.59444
R1103 source.n237 source.n169 6.59444
R1104 source.n492 source.n491 5.81868
R1105 source.n533 source.n468 5.81868
R1106 source.n538 source.n464 5.81868
R1107 source.n580 source.n579 5.81868
R1108 source.n346 source.n345 5.81868
R1109 source.n387 source.n322 5.81868
R1110 source.n392 source.n318 5.81868
R1111 source.n434 source.n433 5.81868
R1112 source.n136 source.n135 5.81868
R1113 source.n95 source.n21 5.81868
R1114 source.n90 source.n25 5.81868
R1115 source.n50 source.n49 5.81868
R1116 source.n282 source.n281 5.81868
R1117 source.n241 source.n167 5.81868
R1118 source.n236 source.n171 5.81868
R1119 source.n196 source.n195 5.81868
R1120 source.n584 source.n583 5.66429
R1121 source.n495 source.n486 5.04292
R1122 source.n530 source.n529 5.04292
R1123 source.n542 source.n541 5.04292
R1124 source.n576 source.n446 5.04292
R1125 source.n349 source.n340 5.04292
R1126 source.n384 source.n383 5.04292
R1127 source.n396 source.n395 5.04292
R1128 source.n430 source.n300 5.04292
R1129 source.n132 source.n2 5.04292
R1130 source.n99 source.n98 5.04292
R1131 source.n87 source.n86 5.04292
R1132 source.n53 source.n44 5.04292
R1133 source.n278 source.n148 5.04292
R1134 source.n245 source.n244 5.04292
R1135 source.n233 source.n232 5.04292
R1136 source.n199 source.n190 5.04292
R1137 source.n496 source.n484 4.26717
R1138 source.n526 source.n470 4.26717
R1139 source.n545 source.n462 4.26717
R1140 source.n575 source.n448 4.26717
R1141 source.n350 source.n338 4.26717
R1142 source.n380 source.n324 4.26717
R1143 source.n399 source.n316 4.26717
R1144 source.n429 source.n302 4.26717
R1145 source.n131 source.n4 4.26717
R1146 source.n102 source.n19 4.26717
R1147 source.n83 source.n27 4.26717
R1148 source.n54 source.n42 4.26717
R1149 source.n277 source.n150 4.26717
R1150 source.n248 source.n165 4.26717
R1151 source.n229 source.n173 4.26717
R1152 source.n200 source.n188 4.26717
R1153 source.n500 source.n499 3.49141
R1154 source.n525 source.n472 3.49141
R1155 source.n546 source.n460 3.49141
R1156 source.n572 source.n571 3.49141
R1157 source.n354 source.n353 3.49141
R1158 source.n379 source.n326 3.49141
R1159 source.n400 source.n314 3.49141
R1160 source.n426 source.n425 3.49141
R1161 source.n128 source.n127 3.49141
R1162 source.n103 source.n17 3.49141
R1163 source.n82 source.n29 3.49141
R1164 source.n58 source.n57 3.49141
R1165 source.n274 source.n273 3.49141
R1166 source.n249 source.n163 3.49141
R1167 source.n228 source.n175 3.49141
R1168 source.n204 source.n203 3.49141
R1169 source.n48 source.n47 2.84303
R1170 source.n194 source.n193 2.84303
R1171 source.n490 source.n489 2.84303
R1172 source.n344 source.n343 2.84303
R1173 source.n503 source.n482 2.71565
R1174 source.n522 source.n521 2.71565
R1175 source.n550 source.n549 2.71565
R1176 source.n568 source.n450 2.71565
R1177 source.n357 source.n336 2.71565
R1178 source.n376 source.n375 2.71565
R1179 source.n404 source.n403 2.71565
R1180 source.n422 source.n304 2.71565
R1181 source.n124 source.n6 2.71565
R1182 source.n107 source.n106 2.71565
R1183 source.n79 source.n78 2.71565
R1184 source.n61 source.n40 2.71565
R1185 source.n270 source.n152 2.71565
R1186 source.n253 source.n252 2.71565
R1187 source.n225 source.n224 2.71565
R1188 source.n207 source.n186 2.71565
R1189 source.n504 source.n480 1.93989
R1190 source.n518 source.n474 1.93989
R1191 source.n554 source.n458 1.93989
R1192 source.n567 source.n452 1.93989
R1193 source.n358 source.n334 1.93989
R1194 source.n372 source.n328 1.93989
R1195 source.n408 source.n312 1.93989
R1196 source.n421 source.n306 1.93989
R1197 source.n123 source.n8 1.93989
R1198 source.n110 source.n14 1.93989
R1199 source.n75 source.n31 1.93989
R1200 source.n62 source.n38 1.93989
R1201 source.n269 source.n154 1.93989
R1202 source.n256 source.n160 1.93989
R1203 source.n221 source.n177 1.93989
R1204 source.n208 source.n184 1.93989
R1205 source.n509 source.n507 1.16414
R1206 source.n517 source.n476 1.16414
R1207 source.n555 source.n456 1.16414
R1208 source.n564 source.n563 1.16414
R1209 source.n363 source.n361 1.16414
R1210 source.n371 source.n330 1.16414
R1211 source.n409 source.n310 1.16414
R1212 source.n418 source.n417 1.16414
R1213 source.n120 source.n119 1.16414
R1214 source.n111 source.n12 1.16414
R1215 source.n74 source.n33 1.16414
R1216 source.n66 source.n65 1.16414
R1217 source.n266 source.n265 1.16414
R1218 source.n257 source.n158 1.16414
R1219 source.n220 source.n179 1.16414
R1220 source.n212 source.n211 1.16414
R1221 source.n285 source.n145 0.87119
R1222 source.n439 source.n437 0.87119
R1223 source.n291 source.n289 0.802224
R1224 source.n289 source.n287 0.802224
R1225 source.n287 source.n285 0.802224
R1226 source.n145 source.n143 0.802224
R1227 source.n143 source.n141 0.802224
R1228 source.n141 source.n139 0.802224
R1229 source.n295 source.n293 0.802224
R1230 source.n297 source.n295 0.802224
R1231 source.n437 source.n297 0.802224
R1232 source.n441 source.n439 0.802224
R1233 source.n443 source.n441 0.802224
R1234 source.n583 source.n443 0.802224
R1235 source.n442 source.t0 0.7925
R1236 source.n442 source.t10 0.7925
R1237 source.n440 source.t3 0.7925
R1238 source.n440 source.t5 0.7925
R1239 source.n438 source.t13 0.7925
R1240 source.n438 source.t9 0.7925
R1241 source.n296 source.t16 0.7925
R1242 source.n296 source.t21 0.7925
R1243 source.n294 source.t24 0.7925
R1244 source.n294 source.t27 0.7925
R1245 source.n292 source.t15 0.7925
R1246 source.n292 source.t23 0.7925
R1247 source.n140 source.t22 0.7925
R1248 source.n140 source.t25 0.7925
R1249 source.n142 source.t19 0.7925
R1250 source.n142 source.t20 0.7925
R1251 source.n144 source.t17 0.7925
R1252 source.n144 source.t18 0.7925
R1253 source.n286 source.t11 0.7925
R1254 source.n286 source.t4 0.7925
R1255 source.n288 source.t12 0.7925
R1256 source.n288 source.t8 0.7925
R1257 source.n290 source.t1 0.7925
R1258 source.n290 source.t2 0.7925
R1259 source.n508 source.n478 0.388379
R1260 source.n514 source.n513 0.388379
R1261 source.n559 source.n558 0.388379
R1262 source.n560 source.n454 0.388379
R1263 source.n362 source.n332 0.388379
R1264 source.n368 source.n367 0.388379
R1265 source.n413 source.n412 0.388379
R1266 source.n414 source.n308 0.388379
R1267 source.n116 source.n10 0.388379
R1268 source.n115 source.n114 0.388379
R1269 source.n71 source.n70 0.388379
R1270 source.n37 source.n35 0.388379
R1271 source.n262 source.n156 0.388379
R1272 source.n261 source.n260 0.388379
R1273 source.n217 source.n216 0.388379
R1274 source.n183 source.n181 0.388379
R1275 source source.n584 0.188
R1276 source.n490 source.n485 0.155672
R1277 source.n497 source.n485 0.155672
R1278 source.n498 source.n497 0.155672
R1279 source.n498 source.n481 0.155672
R1280 source.n505 source.n481 0.155672
R1281 source.n506 source.n505 0.155672
R1282 source.n506 source.n477 0.155672
R1283 source.n515 source.n477 0.155672
R1284 source.n516 source.n515 0.155672
R1285 source.n516 source.n473 0.155672
R1286 source.n523 source.n473 0.155672
R1287 source.n524 source.n523 0.155672
R1288 source.n524 source.n469 0.155672
R1289 source.n531 source.n469 0.155672
R1290 source.n532 source.n531 0.155672
R1291 source.n532 source.n465 0.155672
R1292 source.n539 source.n465 0.155672
R1293 source.n540 source.n539 0.155672
R1294 source.n540 source.n461 0.155672
R1295 source.n547 source.n461 0.155672
R1296 source.n548 source.n547 0.155672
R1297 source.n548 source.n457 0.155672
R1298 source.n556 source.n457 0.155672
R1299 source.n557 source.n556 0.155672
R1300 source.n557 source.n453 0.155672
R1301 source.n565 source.n453 0.155672
R1302 source.n566 source.n565 0.155672
R1303 source.n566 source.n449 0.155672
R1304 source.n573 source.n449 0.155672
R1305 source.n574 source.n573 0.155672
R1306 source.n574 source.n445 0.155672
R1307 source.n581 source.n445 0.155672
R1308 source.n344 source.n339 0.155672
R1309 source.n351 source.n339 0.155672
R1310 source.n352 source.n351 0.155672
R1311 source.n352 source.n335 0.155672
R1312 source.n359 source.n335 0.155672
R1313 source.n360 source.n359 0.155672
R1314 source.n360 source.n331 0.155672
R1315 source.n369 source.n331 0.155672
R1316 source.n370 source.n369 0.155672
R1317 source.n370 source.n327 0.155672
R1318 source.n377 source.n327 0.155672
R1319 source.n378 source.n377 0.155672
R1320 source.n378 source.n323 0.155672
R1321 source.n385 source.n323 0.155672
R1322 source.n386 source.n385 0.155672
R1323 source.n386 source.n319 0.155672
R1324 source.n393 source.n319 0.155672
R1325 source.n394 source.n393 0.155672
R1326 source.n394 source.n315 0.155672
R1327 source.n401 source.n315 0.155672
R1328 source.n402 source.n401 0.155672
R1329 source.n402 source.n311 0.155672
R1330 source.n410 source.n311 0.155672
R1331 source.n411 source.n410 0.155672
R1332 source.n411 source.n307 0.155672
R1333 source.n419 source.n307 0.155672
R1334 source.n420 source.n419 0.155672
R1335 source.n420 source.n303 0.155672
R1336 source.n427 source.n303 0.155672
R1337 source.n428 source.n427 0.155672
R1338 source.n428 source.n299 0.155672
R1339 source.n435 source.n299 0.155672
R1340 source.n137 source.n1 0.155672
R1341 source.n130 source.n1 0.155672
R1342 source.n130 source.n129 0.155672
R1343 source.n129 source.n5 0.155672
R1344 source.n122 source.n5 0.155672
R1345 source.n122 source.n121 0.155672
R1346 source.n121 source.n9 0.155672
R1347 source.n113 source.n9 0.155672
R1348 source.n113 source.n112 0.155672
R1349 source.n112 source.n13 0.155672
R1350 source.n105 source.n13 0.155672
R1351 source.n105 source.n104 0.155672
R1352 source.n104 source.n18 0.155672
R1353 source.n97 source.n18 0.155672
R1354 source.n97 source.n96 0.155672
R1355 source.n96 source.n22 0.155672
R1356 source.n89 source.n22 0.155672
R1357 source.n89 source.n88 0.155672
R1358 source.n88 source.n26 0.155672
R1359 source.n81 source.n26 0.155672
R1360 source.n81 source.n80 0.155672
R1361 source.n80 source.n30 0.155672
R1362 source.n73 source.n30 0.155672
R1363 source.n73 source.n72 0.155672
R1364 source.n72 source.n34 0.155672
R1365 source.n64 source.n34 0.155672
R1366 source.n64 source.n63 0.155672
R1367 source.n63 source.n39 0.155672
R1368 source.n56 source.n39 0.155672
R1369 source.n56 source.n55 0.155672
R1370 source.n55 source.n43 0.155672
R1371 source.n48 source.n43 0.155672
R1372 source.n283 source.n147 0.155672
R1373 source.n276 source.n147 0.155672
R1374 source.n276 source.n275 0.155672
R1375 source.n275 source.n151 0.155672
R1376 source.n268 source.n151 0.155672
R1377 source.n268 source.n267 0.155672
R1378 source.n267 source.n155 0.155672
R1379 source.n259 source.n155 0.155672
R1380 source.n259 source.n258 0.155672
R1381 source.n258 source.n159 0.155672
R1382 source.n251 source.n159 0.155672
R1383 source.n251 source.n250 0.155672
R1384 source.n250 source.n164 0.155672
R1385 source.n243 source.n164 0.155672
R1386 source.n243 source.n242 0.155672
R1387 source.n242 source.n168 0.155672
R1388 source.n235 source.n168 0.155672
R1389 source.n235 source.n234 0.155672
R1390 source.n234 source.n172 0.155672
R1391 source.n227 source.n172 0.155672
R1392 source.n227 source.n226 0.155672
R1393 source.n226 source.n176 0.155672
R1394 source.n219 source.n176 0.155672
R1395 source.n219 source.n218 0.155672
R1396 source.n218 source.n180 0.155672
R1397 source.n210 source.n180 0.155672
R1398 source.n210 source.n209 0.155672
R1399 source.n209 source.n185 0.155672
R1400 source.n202 source.n185 0.155672
R1401 source.n202 source.n201 0.155672
R1402 source.n201 source.n189 0.155672
R1403 source.n194 source.n189 0.155672
R1404 minus.n5 minus.t10 1093.48
R1405 minus.n23 minus.t12 1093.48
R1406 minus.n4 minus.t9 1069.64
R1407 minus.n8 minus.t8 1069.64
R1408 minus.n9 minus.t7 1069.64
R1409 minus.n10 minus.t3 1069.64
R1410 minus.n14 minus.t5 1069.64
R1411 minus.n16 minus.t4 1069.64
R1412 minus.n22 minus.t2 1069.64
R1413 minus.n26 minus.t6 1069.64
R1414 minus.n27 minus.t13 1069.64
R1415 minus.n28 minus.t1 1069.64
R1416 minus.n32 minus.t0 1069.64
R1417 minus.n34 minus.t11 1069.64
R1418 minus.n17 minus.n16 161.3
R1419 minus.n15 minus.n0 161.3
R1420 minus.n14 minus.n13 161.3
R1421 minus.n12 minus.n1 161.3
R1422 minus.n11 minus.n10 161.3
R1423 minus.n8 minus.n7 161.3
R1424 minus.n6 minus.n3 161.3
R1425 minus.n35 minus.n34 161.3
R1426 minus.n33 minus.n18 161.3
R1427 minus.n32 minus.n31 161.3
R1428 minus.n30 minus.n19 161.3
R1429 minus.n29 minus.n28 161.3
R1430 minus.n26 minus.n25 161.3
R1431 minus.n24 minus.n21 161.3
R1432 minus.n9 minus.n2 80.6037
R1433 minus.n27 minus.n20 80.6037
R1434 minus.n9 minus.n8 48.2005
R1435 minus.n10 minus.n9 48.2005
R1436 minus.n27 minus.n26 48.2005
R1437 minus.n28 minus.n27 48.2005
R1438 minus.n36 minus.n17 47.3925
R1439 minus.n4 minus.n3 45.2793
R1440 minus.n14 minus.n1 45.2793
R1441 minus.n22 minus.n21 45.2793
R1442 minus.n32 minus.n19 45.2793
R1443 minus.n6 minus.n5 44.9119
R1444 minus.n24 minus.n23 44.9119
R1445 minus.n16 minus.n15 35.055
R1446 minus.n34 minus.n33 35.055
R1447 minus.n5 minus.n4 17.739
R1448 minus.n23 minus.n22 17.739
R1449 minus.n15 minus.n14 13.146
R1450 minus.n33 minus.n32 13.146
R1451 minus.n36 minus.n35 6.57436
R1452 minus.n8 minus.n3 2.92171
R1453 minus.n10 minus.n1 2.92171
R1454 minus.n26 minus.n21 2.92171
R1455 minus.n28 minus.n19 2.92171
R1456 minus.n11 minus.n2 0.285035
R1457 minus.n7 minus.n2 0.285035
R1458 minus.n25 minus.n20 0.285035
R1459 minus.n29 minus.n20 0.285035
R1460 minus.n17 minus.n0 0.189894
R1461 minus.n13 minus.n0 0.189894
R1462 minus.n13 minus.n12 0.189894
R1463 minus.n12 minus.n11 0.189894
R1464 minus.n7 minus.n6 0.189894
R1465 minus.n25 minus.n24 0.189894
R1466 minus.n30 minus.n29 0.189894
R1467 minus.n31 minus.n30 0.189894
R1468 minus.n31 minus.n18 0.189894
R1469 minus.n35 minus.n18 0.189894
R1470 minus minus.n36 0.188
R1471 drain_right.n134 drain_right.n0 289.615
R1472 drain_right.n284 drain_right.n150 289.615
R1473 drain_right.n44 drain_right.n43 185
R1474 drain_right.n49 drain_right.n48 185
R1475 drain_right.n51 drain_right.n50 185
R1476 drain_right.n40 drain_right.n39 185
R1477 drain_right.n57 drain_right.n56 185
R1478 drain_right.n59 drain_right.n58 185
R1479 drain_right.n36 drain_right.n35 185
R1480 drain_right.n66 drain_right.n65 185
R1481 drain_right.n67 drain_right.n34 185
R1482 drain_right.n69 drain_right.n68 185
R1483 drain_right.n32 drain_right.n31 185
R1484 drain_right.n75 drain_right.n74 185
R1485 drain_right.n77 drain_right.n76 185
R1486 drain_right.n28 drain_right.n27 185
R1487 drain_right.n83 drain_right.n82 185
R1488 drain_right.n85 drain_right.n84 185
R1489 drain_right.n24 drain_right.n23 185
R1490 drain_right.n91 drain_right.n90 185
R1491 drain_right.n93 drain_right.n92 185
R1492 drain_right.n20 drain_right.n19 185
R1493 drain_right.n99 drain_right.n98 185
R1494 drain_right.n101 drain_right.n100 185
R1495 drain_right.n16 drain_right.n15 185
R1496 drain_right.n107 drain_right.n106 185
R1497 drain_right.n110 drain_right.n109 185
R1498 drain_right.n108 drain_right.n12 185
R1499 drain_right.n115 drain_right.n11 185
R1500 drain_right.n117 drain_right.n116 185
R1501 drain_right.n119 drain_right.n118 185
R1502 drain_right.n8 drain_right.n7 185
R1503 drain_right.n125 drain_right.n124 185
R1504 drain_right.n127 drain_right.n126 185
R1505 drain_right.n4 drain_right.n3 185
R1506 drain_right.n133 drain_right.n132 185
R1507 drain_right.n135 drain_right.n134 185
R1508 drain_right.n285 drain_right.n284 185
R1509 drain_right.n283 drain_right.n282 185
R1510 drain_right.n154 drain_right.n153 185
R1511 drain_right.n277 drain_right.n276 185
R1512 drain_right.n275 drain_right.n274 185
R1513 drain_right.n158 drain_right.n157 185
R1514 drain_right.n269 drain_right.n268 185
R1515 drain_right.n267 drain_right.n266 185
R1516 drain_right.n265 drain_right.n161 185
R1517 drain_right.n165 drain_right.n162 185
R1518 drain_right.n260 drain_right.n259 185
R1519 drain_right.n258 drain_right.n257 185
R1520 drain_right.n167 drain_right.n166 185
R1521 drain_right.n252 drain_right.n251 185
R1522 drain_right.n250 drain_right.n249 185
R1523 drain_right.n171 drain_right.n170 185
R1524 drain_right.n244 drain_right.n243 185
R1525 drain_right.n242 drain_right.n241 185
R1526 drain_right.n175 drain_right.n174 185
R1527 drain_right.n236 drain_right.n235 185
R1528 drain_right.n234 drain_right.n233 185
R1529 drain_right.n179 drain_right.n178 185
R1530 drain_right.n228 drain_right.n227 185
R1531 drain_right.n226 drain_right.n225 185
R1532 drain_right.n183 drain_right.n182 185
R1533 drain_right.n220 drain_right.n219 185
R1534 drain_right.n218 drain_right.n185 185
R1535 drain_right.n217 drain_right.n216 185
R1536 drain_right.n188 drain_right.n186 185
R1537 drain_right.n211 drain_right.n210 185
R1538 drain_right.n209 drain_right.n208 185
R1539 drain_right.n192 drain_right.n191 185
R1540 drain_right.n203 drain_right.n202 185
R1541 drain_right.n201 drain_right.n200 185
R1542 drain_right.n196 drain_right.n195 185
R1543 drain_right.n45 drain_right.t1 149.524
R1544 drain_right.n197 drain_right.t9 149.524
R1545 drain_right.n49 drain_right.n43 104.615
R1546 drain_right.n50 drain_right.n49 104.615
R1547 drain_right.n50 drain_right.n39 104.615
R1548 drain_right.n57 drain_right.n39 104.615
R1549 drain_right.n58 drain_right.n57 104.615
R1550 drain_right.n58 drain_right.n35 104.615
R1551 drain_right.n66 drain_right.n35 104.615
R1552 drain_right.n67 drain_right.n66 104.615
R1553 drain_right.n68 drain_right.n67 104.615
R1554 drain_right.n68 drain_right.n31 104.615
R1555 drain_right.n75 drain_right.n31 104.615
R1556 drain_right.n76 drain_right.n75 104.615
R1557 drain_right.n76 drain_right.n27 104.615
R1558 drain_right.n83 drain_right.n27 104.615
R1559 drain_right.n84 drain_right.n83 104.615
R1560 drain_right.n84 drain_right.n23 104.615
R1561 drain_right.n91 drain_right.n23 104.615
R1562 drain_right.n92 drain_right.n91 104.615
R1563 drain_right.n92 drain_right.n19 104.615
R1564 drain_right.n99 drain_right.n19 104.615
R1565 drain_right.n100 drain_right.n99 104.615
R1566 drain_right.n100 drain_right.n15 104.615
R1567 drain_right.n107 drain_right.n15 104.615
R1568 drain_right.n109 drain_right.n107 104.615
R1569 drain_right.n109 drain_right.n108 104.615
R1570 drain_right.n108 drain_right.n11 104.615
R1571 drain_right.n117 drain_right.n11 104.615
R1572 drain_right.n118 drain_right.n117 104.615
R1573 drain_right.n118 drain_right.n7 104.615
R1574 drain_right.n125 drain_right.n7 104.615
R1575 drain_right.n126 drain_right.n125 104.615
R1576 drain_right.n126 drain_right.n3 104.615
R1577 drain_right.n133 drain_right.n3 104.615
R1578 drain_right.n134 drain_right.n133 104.615
R1579 drain_right.n284 drain_right.n283 104.615
R1580 drain_right.n283 drain_right.n153 104.615
R1581 drain_right.n276 drain_right.n153 104.615
R1582 drain_right.n276 drain_right.n275 104.615
R1583 drain_right.n275 drain_right.n157 104.615
R1584 drain_right.n268 drain_right.n157 104.615
R1585 drain_right.n268 drain_right.n267 104.615
R1586 drain_right.n267 drain_right.n161 104.615
R1587 drain_right.n165 drain_right.n161 104.615
R1588 drain_right.n259 drain_right.n165 104.615
R1589 drain_right.n259 drain_right.n258 104.615
R1590 drain_right.n258 drain_right.n166 104.615
R1591 drain_right.n251 drain_right.n166 104.615
R1592 drain_right.n251 drain_right.n250 104.615
R1593 drain_right.n250 drain_right.n170 104.615
R1594 drain_right.n243 drain_right.n170 104.615
R1595 drain_right.n243 drain_right.n242 104.615
R1596 drain_right.n242 drain_right.n174 104.615
R1597 drain_right.n235 drain_right.n174 104.615
R1598 drain_right.n235 drain_right.n234 104.615
R1599 drain_right.n234 drain_right.n178 104.615
R1600 drain_right.n227 drain_right.n178 104.615
R1601 drain_right.n227 drain_right.n226 104.615
R1602 drain_right.n226 drain_right.n182 104.615
R1603 drain_right.n219 drain_right.n182 104.615
R1604 drain_right.n219 drain_right.n218 104.615
R1605 drain_right.n218 drain_right.n217 104.615
R1606 drain_right.n217 drain_right.n186 104.615
R1607 drain_right.n210 drain_right.n186 104.615
R1608 drain_right.n210 drain_right.n209 104.615
R1609 drain_right.n209 drain_right.n191 104.615
R1610 drain_right.n202 drain_right.n191 104.615
R1611 drain_right.n202 drain_right.n201 104.615
R1612 drain_right.n201 drain_right.n195 104.615
R1613 drain_right.n143 drain_right.n141 59.5172
R1614 drain_right.n147 drain_right.n145 59.517
R1615 drain_right.n143 drain_right.n142 58.7154
R1616 drain_right.n140 drain_right.n139 58.7154
R1617 drain_right.n147 drain_right.n146 58.7154
R1618 drain_right.n149 drain_right.n148 58.7154
R1619 drain_right.t1 drain_right.n43 52.3082
R1620 drain_right.t9 drain_right.n195 52.3082
R1621 drain_right.n140 drain_right.n138 48.1143
R1622 drain_right.n289 drain_right.n288 47.3126
R1623 drain_right drain_right.n144 41.2722
R1624 drain_right.n69 drain_right.n34 13.1884
R1625 drain_right.n116 drain_right.n115 13.1884
R1626 drain_right.n266 drain_right.n265 13.1884
R1627 drain_right.n220 drain_right.n185 13.1884
R1628 drain_right.n65 drain_right.n64 12.8005
R1629 drain_right.n70 drain_right.n32 12.8005
R1630 drain_right.n114 drain_right.n12 12.8005
R1631 drain_right.n119 drain_right.n10 12.8005
R1632 drain_right.n269 drain_right.n160 12.8005
R1633 drain_right.n264 drain_right.n162 12.8005
R1634 drain_right.n221 drain_right.n183 12.8005
R1635 drain_right.n216 drain_right.n187 12.8005
R1636 drain_right.n63 drain_right.n36 12.0247
R1637 drain_right.n74 drain_right.n73 12.0247
R1638 drain_right.n111 drain_right.n110 12.0247
R1639 drain_right.n120 drain_right.n8 12.0247
R1640 drain_right.n270 drain_right.n158 12.0247
R1641 drain_right.n261 drain_right.n260 12.0247
R1642 drain_right.n225 drain_right.n224 12.0247
R1643 drain_right.n215 drain_right.n188 12.0247
R1644 drain_right.n60 drain_right.n59 11.249
R1645 drain_right.n77 drain_right.n30 11.249
R1646 drain_right.n106 drain_right.n14 11.249
R1647 drain_right.n124 drain_right.n123 11.249
R1648 drain_right.n274 drain_right.n273 11.249
R1649 drain_right.n257 drain_right.n164 11.249
R1650 drain_right.n228 drain_right.n181 11.249
R1651 drain_right.n212 drain_right.n211 11.249
R1652 drain_right.n56 drain_right.n38 10.4732
R1653 drain_right.n78 drain_right.n28 10.4732
R1654 drain_right.n105 drain_right.n16 10.4732
R1655 drain_right.n127 drain_right.n6 10.4732
R1656 drain_right.n277 drain_right.n156 10.4732
R1657 drain_right.n256 drain_right.n167 10.4732
R1658 drain_right.n229 drain_right.n179 10.4732
R1659 drain_right.n208 drain_right.n190 10.4732
R1660 drain_right.n45 drain_right.n44 10.2747
R1661 drain_right.n197 drain_right.n196 10.2747
R1662 drain_right.n55 drain_right.n40 9.69747
R1663 drain_right.n82 drain_right.n81 9.69747
R1664 drain_right.n102 drain_right.n101 9.69747
R1665 drain_right.n128 drain_right.n4 9.69747
R1666 drain_right.n278 drain_right.n154 9.69747
R1667 drain_right.n253 drain_right.n252 9.69747
R1668 drain_right.n233 drain_right.n232 9.69747
R1669 drain_right.n207 drain_right.n192 9.69747
R1670 drain_right.n138 drain_right.n137 9.45567
R1671 drain_right.n288 drain_right.n287 9.45567
R1672 drain_right.n2 drain_right.n1 9.3005
R1673 drain_right.n131 drain_right.n130 9.3005
R1674 drain_right.n129 drain_right.n128 9.3005
R1675 drain_right.n6 drain_right.n5 9.3005
R1676 drain_right.n123 drain_right.n122 9.3005
R1677 drain_right.n121 drain_right.n120 9.3005
R1678 drain_right.n10 drain_right.n9 9.3005
R1679 drain_right.n89 drain_right.n88 9.3005
R1680 drain_right.n87 drain_right.n86 9.3005
R1681 drain_right.n26 drain_right.n25 9.3005
R1682 drain_right.n81 drain_right.n80 9.3005
R1683 drain_right.n79 drain_right.n78 9.3005
R1684 drain_right.n30 drain_right.n29 9.3005
R1685 drain_right.n73 drain_right.n72 9.3005
R1686 drain_right.n71 drain_right.n70 9.3005
R1687 drain_right.n47 drain_right.n46 9.3005
R1688 drain_right.n42 drain_right.n41 9.3005
R1689 drain_right.n53 drain_right.n52 9.3005
R1690 drain_right.n55 drain_right.n54 9.3005
R1691 drain_right.n38 drain_right.n37 9.3005
R1692 drain_right.n61 drain_right.n60 9.3005
R1693 drain_right.n63 drain_right.n62 9.3005
R1694 drain_right.n64 drain_right.n33 9.3005
R1695 drain_right.n22 drain_right.n21 9.3005
R1696 drain_right.n95 drain_right.n94 9.3005
R1697 drain_right.n97 drain_right.n96 9.3005
R1698 drain_right.n18 drain_right.n17 9.3005
R1699 drain_right.n103 drain_right.n102 9.3005
R1700 drain_right.n105 drain_right.n104 9.3005
R1701 drain_right.n14 drain_right.n13 9.3005
R1702 drain_right.n112 drain_right.n111 9.3005
R1703 drain_right.n114 drain_right.n113 9.3005
R1704 drain_right.n137 drain_right.n136 9.3005
R1705 drain_right.n199 drain_right.n198 9.3005
R1706 drain_right.n194 drain_right.n193 9.3005
R1707 drain_right.n205 drain_right.n204 9.3005
R1708 drain_right.n207 drain_right.n206 9.3005
R1709 drain_right.n190 drain_right.n189 9.3005
R1710 drain_right.n213 drain_right.n212 9.3005
R1711 drain_right.n215 drain_right.n214 9.3005
R1712 drain_right.n187 drain_right.n184 9.3005
R1713 drain_right.n246 drain_right.n245 9.3005
R1714 drain_right.n248 drain_right.n247 9.3005
R1715 drain_right.n169 drain_right.n168 9.3005
R1716 drain_right.n254 drain_right.n253 9.3005
R1717 drain_right.n256 drain_right.n255 9.3005
R1718 drain_right.n164 drain_right.n163 9.3005
R1719 drain_right.n262 drain_right.n261 9.3005
R1720 drain_right.n264 drain_right.n263 9.3005
R1721 drain_right.n287 drain_right.n286 9.3005
R1722 drain_right.n152 drain_right.n151 9.3005
R1723 drain_right.n281 drain_right.n280 9.3005
R1724 drain_right.n279 drain_right.n278 9.3005
R1725 drain_right.n156 drain_right.n155 9.3005
R1726 drain_right.n273 drain_right.n272 9.3005
R1727 drain_right.n271 drain_right.n270 9.3005
R1728 drain_right.n160 drain_right.n159 9.3005
R1729 drain_right.n173 drain_right.n172 9.3005
R1730 drain_right.n240 drain_right.n239 9.3005
R1731 drain_right.n238 drain_right.n237 9.3005
R1732 drain_right.n177 drain_right.n176 9.3005
R1733 drain_right.n232 drain_right.n231 9.3005
R1734 drain_right.n230 drain_right.n229 9.3005
R1735 drain_right.n181 drain_right.n180 9.3005
R1736 drain_right.n224 drain_right.n223 9.3005
R1737 drain_right.n222 drain_right.n221 9.3005
R1738 drain_right.n52 drain_right.n51 8.92171
R1739 drain_right.n85 drain_right.n26 8.92171
R1740 drain_right.n98 drain_right.n18 8.92171
R1741 drain_right.n132 drain_right.n131 8.92171
R1742 drain_right.n282 drain_right.n281 8.92171
R1743 drain_right.n249 drain_right.n169 8.92171
R1744 drain_right.n236 drain_right.n177 8.92171
R1745 drain_right.n204 drain_right.n203 8.92171
R1746 drain_right.n48 drain_right.n42 8.14595
R1747 drain_right.n86 drain_right.n24 8.14595
R1748 drain_right.n97 drain_right.n20 8.14595
R1749 drain_right.n135 drain_right.n2 8.14595
R1750 drain_right.n285 drain_right.n152 8.14595
R1751 drain_right.n248 drain_right.n171 8.14595
R1752 drain_right.n237 drain_right.n175 8.14595
R1753 drain_right.n200 drain_right.n194 8.14595
R1754 drain_right.n47 drain_right.n44 7.3702
R1755 drain_right.n90 drain_right.n89 7.3702
R1756 drain_right.n94 drain_right.n93 7.3702
R1757 drain_right.n136 drain_right.n0 7.3702
R1758 drain_right.n286 drain_right.n150 7.3702
R1759 drain_right.n245 drain_right.n244 7.3702
R1760 drain_right.n241 drain_right.n240 7.3702
R1761 drain_right.n199 drain_right.n196 7.3702
R1762 drain_right.n90 drain_right.n22 6.59444
R1763 drain_right.n93 drain_right.n22 6.59444
R1764 drain_right.n138 drain_right.n0 6.59444
R1765 drain_right.n288 drain_right.n150 6.59444
R1766 drain_right.n244 drain_right.n173 6.59444
R1767 drain_right.n241 drain_right.n173 6.59444
R1768 drain_right drain_right.n289 6.05408
R1769 drain_right.n48 drain_right.n47 5.81868
R1770 drain_right.n89 drain_right.n24 5.81868
R1771 drain_right.n94 drain_right.n20 5.81868
R1772 drain_right.n136 drain_right.n135 5.81868
R1773 drain_right.n286 drain_right.n285 5.81868
R1774 drain_right.n245 drain_right.n171 5.81868
R1775 drain_right.n240 drain_right.n175 5.81868
R1776 drain_right.n200 drain_right.n199 5.81868
R1777 drain_right.n51 drain_right.n42 5.04292
R1778 drain_right.n86 drain_right.n85 5.04292
R1779 drain_right.n98 drain_right.n97 5.04292
R1780 drain_right.n132 drain_right.n2 5.04292
R1781 drain_right.n282 drain_right.n152 5.04292
R1782 drain_right.n249 drain_right.n248 5.04292
R1783 drain_right.n237 drain_right.n236 5.04292
R1784 drain_right.n203 drain_right.n194 5.04292
R1785 drain_right.n52 drain_right.n40 4.26717
R1786 drain_right.n82 drain_right.n26 4.26717
R1787 drain_right.n101 drain_right.n18 4.26717
R1788 drain_right.n131 drain_right.n4 4.26717
R1789 drain_right.n281 drain_right.n154 4.26717
R1790 drain_right.n252 drain_right.n169 4.26717
R1791 drain_right.n233 drain_right.n177 4.26717
R1792 drain_right.n204 drain_right.n192 4.26717
R1793 drain_right.n56 drain_right.n55 3.49141
R1794 drain_right.n81 drain_right.n28 3.49141
R1795 drain_right.n102 drain_right.n16 3.49141
R1796 drain_right.n128 drain_right.n127 3.49141
R1797 drain_right.n278 drain_right.n277 3.49141
R1798 drain_right.n253 drain_right.n167 3.49141
R1799 drain_right.n232 drain_right.n179 3.49141
R1800 drain_right.n208 drain_right.n207 3.49141
R1801 drain_right.n198 drain_right.n197 2.84303
R1802 drain_right.n46 drain_right.n45 2.84303
R1803 drain_right.n59 drain_right.n38 2.71565
R1804 drain_right.n78 drain_right.n77 2.71565
R1805 drain_right.n106 drain_right.n105 2.71565
R1806 drain_right.n124 drain_right.n6 2.71565
R1807 drain_right.n274 drain_right.n156 2.71565
R1808 drain_right.n257 drain_right.n256 2.71565
R1809 drain_right.n229 drain_right.n228 2.71565
R1810 drain_right.n211 drain_right.n190 2.71565
R1811 drain_right.n60 drain_right.n36 1.93989
R1812 drain_right.n74 drain_right.n30 1.93989
R1813 drain_right.n110 drain_right.n14 1.93989
R1814 drain_right.n123 drain_right.n8 1.93989
R1815 drain_right.n273 drain_right.n158 1.93989
R1816 drain_right.n260 drain_right.n164 1.93989
R1817 drain_right.n225 drain_right.n181 1.93989
R1818 drain_right.n212 drain_right.n188 1.93989
R1819 drain_right.n65 drain_right.n63 1.16414
R1820 drain_right.n73 drain_right.n32 1.16414
R1821 drain_right.n111 drain_right.n12 1.16414
R1822 drain_right.n120 drain_right.n119 1.16414
R1823 drain_right.n270 drain_right.n269 1.16414
R1824 drain_right.n261 drain_right.n162 1.16414
R1825 drain_right.n224 drain_right.n183 1.16414
R1826 drain_right.n216 drain_right.n215 1.16414
R1827 drain_right.n289 drain_right.n149 0.802224
R1828 drain_right.n149 drain_right.n147 0.802224
R1829 drain_right.n141 drain_right.t13 0.7925
R1830 drain_right.n141 drain_right.t2 0.7925
R1831 drain_right.n142 drain_right.t0 0.7925
R1832 drain_right.n142 drain_right.t12 0.7925
R1833 drain_right.n139 drain_right.t11 0.7925
R1834 drain_right.n139 drain_right.t7 0.7925
R1835 drain_right.n145 drain_right.t4 0.7925
R1836 drain_right.n145 drain_right.t3 0.7925
R1837 drain_right.n146 drain_right.t6 0.7925
R1838 drain_right.n146 drain_right.t5 0.7925
R1839 drain_right.n148 drain_right.t8 0.7925
R1840 drain_right.n148 drain_right.t10 0.7925
R1841 drain_right.n144 drain_right.n140 0.546447
R1842 drain_right.n64 drain_right.n34 0.388379
R1843 drain_right.n70 drain_right.n69 0.388379
R1844 drain_right.n115 drain_right.n114 0.388379
R1845 drain_right.n116 drain_right.n10 0.388379
R1846 drain_right.n266 drain_right.n160 0.388379
R1847 drain_right.n265 drain_right.n264 0.388379
R1848 drain_right.n221 drain_right.n220 0.388379
R1849 drain_right.n187 drain_right.n185 0.388379
R1850 drain_right.n46 drain_right.n41 0.155672
R1851 drain_right.n53 drain_right.n41 0.155672
R1852 drain_right.n54 drain_right.n53 0.155672
R1853 drain_right.n54 drain_right.n37 0.155672
R1854 drain_right.n61 drain_right.n37 0.155672
R1855 drain_right.n62 drain_right.n61 0.155672
R1856 drain_right.n62 drain_right.n33 0.155672
R1857 drain_right.n71 drain_right.n33 0.155672
R1858 drain_right.n72 drain_right.n71 0.155672
R1859 drain_right.n72 drain_right.n29 0.155672
R1860 drain_right.n79 drain_right.n29 0.155672
R1861 drain_right.n80 drain_right.n79 0.155672
R1862 drain_right.n80 drain_right.n25 0.155672
R1863 drain_right.n87 drain_right.n25 0.155672
R1864 drain_right.n88 drain_right.n87 0.155672
R1865 drain_right.n88 drain_right.n21 0.155672
R1866 drain_right.n95 drain_right.n21 0.155672
R1867 drain_right.n96 drain_right.n95 0.155672
R1868 drain_right.n96 drain_right.n17 0.155672
R1869 drain_right.n103 drain_right.n17 0.155672
R1870 drain_right.n104 drain_right.n103 0.155672
R1871 drain_right.n104 drain_right.n13 0.155672
R1872 drain_right.n112 drain_right.n13 0.155672
R1873 drain_right.n113 drain_right.n112 0.155672
R1874 drain_right.n113 drain_right.n9 0.155672
R1875 drain_right.n121 drain_right.n9 0.155672
R1876 drain_right.n122 drain_right.n121 0.155672
R1877 drain_right.n122 drain_right.n5 0.155672
R1878 drain_right.n129 drain_right.n5 0.155672
R1879 drain_right.n130 drain_right.n129 0.155672
R1880 drain_right.n130 drain_right.n1 0.155672
R1881 drain_right.n137 drain_right.n1 0.155672
R1882 drain_right.n287 drain_right.n151 0.155672
R1883 drain_right.n280 drain_right.n151 0.155672
R1884 drain_right.n280 drain_right.n279 0.155672
R1885 drain_right.n279 drain_right.n155 0.155672
R1886 drain_right.n272 drain_right.n155 0.155672
R1887 drain_right.n272 drain_right.n271 0.155672
R1888 drain_right.n271 drain_right.n159 0.155672
R1889 drain_right.n263 drain_right.n159 0.155672
R1890 drain_right.n263 drain_right.n262 0.155672
R1891 drain_right.n262 drain_right.n163 0.155672
R1892 drain_right.n255 drain_right.n163 0.155672
R1893 drain_right.n255 drain_right.n254 0.155672
R1894 drain_right.n254 drain_right.n168 0.155672
R1895 drain_right.n247 drain_right.n168 0.155672
R1896 drain_right.n247 drain_right.n246 0.155672
R1897 drain_right.n246 drain_right.n172 0.155672
R1898 drain_right.n239 drain_right.n172 0.155672
R1899 drain_right.n239 drain_right.n238 0.155672
R1900 drain_right.n238 drain_right.n176 0.155672
R1901 drain_right.n231 drain_right.n176 0.155672
R1902 drain_right.n231 drain_right.n230 0.155672
R1903 drain_right.n230 drain_right.n180 0.155672
R1904 drain_right.n223 drain_right.n180 0.155672
R1905 drain_right.n223 drain_right.n222 0.155672
R1906 drain_right.n222 drain_right.n184 0.155672
R1907 drain_right.n214 drain_right.n184 0.155672
R1908 drain_right.n214 drain_right.n213 0.155672
R1909 drain_right.n213 drain_right.n189 0.155672
R1910 drain_right.n206 drain_right.n189 0.155672
R1911 drain_right.n206 drain_right.n205 0.155672
R1912 drain_right.n205 drain_right.n193 0.155672
R1913 drain_right.n198 drain_right.n193 0.155672
R1914 drain_right.n144 drain_right.n143 0.145585
C0 minus drain_left 0.172803f
C1 drain_right drain_left 1.15268f
C2 plus drain_left 16.9329f
C3 source drain_left 38.4673f
C4 drain_right minus 16.721401f
C5 plus minus 8.30565f
C6 minus source 16.114f
C7 drain_right plus 0.37654f
C8 drain_right source 38.4513f
C9 plus source 16.129099f
C10 drain_right a_n2204_n5888# 11.04566f
C11 drain_left a_n2204_n5888# 11.374969f
C12 source a_n2204_n5888# 11.246991f
C13 minus a_n2204_n5888# 9.59493f
C14 plus a_n2204_n5888# 12.06242f
C15 drain_right.n0 a_n2204_n5888# 0.035452f
C16 drain_right.n1 a_n2204_n5888# 0.025716f
C17 drain_right.n2 a_n2204_n5888# 0.013819f
C18 drain_right.n3 a_n2204_n5888# 0.032662f
C19 drain_right.n4 a_n2204_n5888# 0.014631f
C20 drain_right.n5 a_n2204_n5888# 0.025716f
C21 drain_right.n6 a_n2204_n5888# 0.013819f
C22 drain_right.n7 a_n2204_n5888# 0.032662f
C23 drain_right.n8 a_n2204_n5888# 0.014631f
C24 drain_right.n9 a_n2204_n5888# 0.025716f
C25 drain_right.n10 a_n2204_n5888# 0.013819f
C26 drain_right.n11 a_n2204_n5888# 0.032662f
C27 drain_right.n12 a_n2204_n5888# 0.014631f
C28 drain_right.n13 a_n2204_n5888# 0.025716f
C29 drain_right.n14 a_n2204_n5888# 0.013819f
C30 drain_right.n15 a_n2204_n5888# 0.032662f
C31 drain_right.n16 a_n2204_n5888# 0.014631f
C32 drain_right.n17 a_n2204_n5888# 0.025716f
C33 drain_right.n18 a_n2204_n5888# 0.013819f
C34 drain_right.n19 a_n2204_n5888# 0.032662f
C35 drain_right.n20 a_n2204_n5888# 0.014631f
C36 drain_right.n21 a_n2204_n5888# 0.025716f
C37 drain_right.n22 a_n2204_n5888# 0.013819f
C38 drain_right.n23 a_n2204_n5888# 0.032662f
C39 drain_right.n24 a_n2204_n5888# 0.014631f
C40 drain_right.n25 a_n2204_n5888# 0.025716f
C41 drain_right.n26 a_n2204_n5888# 0.013819f
C42 drain_right.n27 a_n2204_n5888# 0.032662f
C43 drain_right.n28 a_n2204_n5888# 0.014631f
C44 drain_right.n29 a_n2204_n5888# 0.025716f
C45 drain_right.n30 a_n2204_n5888# 0.013819f
C46 drain_right.n31 a_n2204_n5888# 0.032662f
C47 drain_right.n32 a_n2204_n5888# 0.014631f
C48 drain_right.n33 a_n2204_n5888# 0.025716f
C49 drain_right.n34 a_n2204_n5888# 0.014225f
C50 drain_right.n35 a_n2204_n5888# 0.032662f
C51 drain_right.n36 a_n2204_n5888# 0.014631f
C52 drain_right.n37 a_n2204_n5888# 0.025716f
C53 drain_right.n38 a_n2204_n5888# 0.013819f
C54 drain_right.n39 a_n2204_n5888# 0.032662f
C55 drain_right.n40 a_n2204_n5888# 0.014631f
C56 drain_right.n41 a_n2204_n5888# 0.025716f
C57 drain_right.n42 a_n2204_n5888# 0.013819f
C58 drain_right.n43 a_n2204_n5888# 0.024497f
C59 drain_right.n44 a_n2204_n5888# 0.02309f
C60 drain_right.t1 a_n2204_n5888# 0.056965f
C61 drain_right.n45 a_n2204_n5888# 0.313756f
C62 drain_right.n46 a_n2204_n5888# 2.78428f
C63 drain_right.n47 a_n2204_n5888# 0.013819f
C64 drain_right.n48 a_n2204_n5888# 0.014631f
C65 drain_right.n49 a_n2204_n5888# 0.032662f
C66 drain_right.n50 a_n2204_n5888# 0.032662f
C67 drain_right.n51 a_n2204_n5888# 0.014631f
C68 drain_right.n52 a_n2204_n5888# 0.013819f
C69 drain_right.n53 a_n2204_n5888# 0.025716f
C70 drain_right.n54 a_n2204_n5888# 0.025716f
C71 drain_right.n55 a_n2204_n5888# 0.013819f
C72 drain_right.n56 a_n2204_n5888# 0.014631f
C73 drain_right.n57 a_n2204_n5888# 0.032662f
C74 drain_right.n58 a_n2204_n5888# 0.032662f
C75 drain_right.n59 a_n2204_n5888# 0.014631f
C76 drain_right.n60 a_n2204_n5888# 0.013819f
C77 drain_right.n61 a_n2204_n5888# 0.025716f
C78 drain_right.n62 a_n2204_n5888# 0.025716f
C79 drain_right.n63 a_n2204_n5888# 0.013819f
C80 drain_right.n64 a_n2204_n5888# 0.013819f
C81 drain_right.n65 a_n2204_n5888# 0.014631f
C82 drain_right.n66 a_n2204_n5888# 0.032662f
C83 drain_right.n67 a_n2204_n5888# 0.032662f
C84 drain_right.n68 a_n2204_n5888# 0.032662f
C85 drain_right.n69 a_n2204_n5888# 0.014225f
C86 drain_right.n70 a_n2204_n5888# 0.013819f
C87 drain_right.n71 a_n2204_n5888# 0.025716f
C88 drain_right.n72 a_n2204_n5888# 0.025716f
C89 drain_right.n73 a_n2204_n5888# 0.013819f
C90 drain_right.n74 a_n2204_n5888# 0.014631f
C91 drain_right.n75 a_n2204_n5888# 0.032662f
C92 drain_right.n76 a_n2204_n5888# 0.032662f
C93 drain_right.n77 a_n2204_n5888# 0.014631f
C94 drain_right.n78 a_n2204_n5888# 0.013819f
C95 drain_right.n79 a_n2204_n5888# 0.025716f
C96 drain_right.n80 a_n2204_n5888# 0.025716f
C97 drain_right.n81 a_n2204_n5888# 0.013819f
C98 drain_right.n82 a_n2204_n5888# 0.014631f
C99 drain_right.n83 a_n2204_n5888# 0.032662f
C100 drain_right.n84 a_n2204_n5888# 0.032662f
C101 drain_right.n85 a_n2204_n5888# 0.014631f
C102 drain_right.n86 a_n2204_n5888# 0.013819f
C103 drain_right.n87 a_n2204_n5888# 0.025716f
C104 drain_right.n88 a_n2204_n5888# 0.025716f
C105 drain_right.n89 a_n2204_n5888# 0.013819f
C106 drain_right.n90 a_n2204_n5888# 0.014631f
C107 drain_right.n91 a_n2204_n5888# 0.032662f
C108 drain_right.n92 a_n2204_n5888# 0.032662f
C109 drain_right.n93 a_n2204_n5888# 0.014631f
C110 drain_right.n94 a_n2204_n5888# 0.013819f
C111 drain_right.n95 a_n2204_n5888# 0.025716f
C112 drain_right.n96 a_n2204_n5888# 0.025716f
C113 drain_right.n97 a_n2204_n5888# 0.013819f
C114 drain_right.n98 a_n2204_n5888# 0.014631f
C115 drain_right.n99 a_n2204_n5888# 0.032662f
C116 drain_right.n100 a_n2204_n5888# 0.032662f
C117 drain_right.n101 a_n2204_n5888# 0.014631f
C118 drain_right.n102 a_n2204_n5888# 0.013819f
C119 drain_right.n103 a_n2204_n5888# 0.025716f
C120 drain_right.n104 a_n2204_n5888# 0.025716f
C121 drain_right.n105 a_n2204_n5888# 0.013819f
C122 drain_right.n106 a_n2204_n5888# 0.014631f
C123 drain_right.n107 a_n2204_n5888# 0.032662f
C124 drain_right.n108 a_n2204_n5888# 0.032662f
C125 drain_right.n109 a_n2204_n5888# 0.032662f
C126 drain_right.n110 a_n2204_n5888# 0.014631f
C127 drain_right.n111 a_n2204_n5888# 0.013819f
C128 drain_right.n112 a_n2204_n5888# 0.025716f
C129 drain_right.n113 a_n2204_n5888# 0.025716f
C130 drain_right.n114 a_n2204_n5888# 0.013819f
C131 drain_right.n115 a_n2204_n5888# 0.014225f
C132 drain_right.n116 a_n2204_n5888# 0.014225f
C133 drain_right.n117 a_n2204_n5888# 0.032662f
C134 drain_right.n118 a_n2204_n5888# 0.032662f
C135 drain_right.n119 a_n2204_n5888# 0.014631f
C136 drain_right.n120 a_n2204_n5888# 0.013819f
C137 drain_right.n121 a_n2204_n5888# 0.025716f
C138 drain_right.n122 a_n2204_n5888# 0.025716f
C139 drain_right.n123 a_n2204_n5888# 0.013819f
C140 drain_right.n124 a_n2204_n5888# 0.014631f
C141 drain_right.n125 a_n2204_n5888# 0.032662f
C142 drain_right.n126 a_n2204_n5888# 0.032662f
C143 drain_right.n127 a_n2204_n5888# 0.014631f
C144 drain_right.n128 a_n2204_n5888# 0.013819f
C145 drain_right.n129 a_n2204_n5888# 0.025716f
C146 drain_right.n130 a_n2204_n5888# 0.025716f
C147 drain_right.n131 a_n2204_n5888# 0.013819f
C148 drain_right.n132 a_n2204_n5888# 0.014631f
C149 drain_right.n133 a_n2204_n5888# 0.032662f
C150 drain_right.n134 a_n2204_n5888# 0.069481f
C151 drain_right.n135 a_n2204_n5888# 0.014631f
C152 drain_right.n136 a_n2204_n5888# 0.013819f
C153 drain_right.n137 a_n2204_n5888# 0.056631f
C154 drain_right.n138 a_n2204_n5888# 0.058348f
C155 drain_right.t11 a_n2204_n5888# 0.508038f
C156 drain_right.t7 a_n2204_n5888# 0.508038f
C157 drain_right.n139 a_n2204_n5888# 4.68212f
C158 drain_right.n140 a_n2204_n5888# 0.442576f
C159 drain_right.t13 a_n2204_n5888# 0.508038f
C160 drain_right.t2 a_n2204_n5888# 0.508038f
C161 drain_right.n141 a_n2204_n5888# 4.68698f
C162 drain_right.t0 a_n2204_n5888# 0.508038f
C163 drain_right.t12 a_n2204_n5888# 0.508038f
C164 drain_right.n142 a_n2204_n5888# 4.68212f
C165 drain_right.n143 a_n2204_n5888# 0.65568f
C166 drain_right.n144 a_n2204_n5888# 2.16085f
C167 drain_right.t4 a_n2204_n5888# 0.508038f
C168 drain_right.t3 a_n2204_n5888# 0.508038f
C169 drain_right.n145 a_n2204_n5888# 4.68697f
C170 drain_right.t6 a_n2204_n5888# 0.508038f
C171 drain_right.t5 a_n2204_n5888# 0.508038f
C172 drain_right.n146 a_n2204_n5888# 4.68212f
C173 drain_right.n147 a_n2204_n5888# 0.70599f
C174 drain_right.t8 a_n2204_n5888# 0.508038f
C175 drain_right.t10 a_n2204_n5888# 0.508038f
C176 drain_right.n148 a_n2204_n5888# 4.68212f
C177 drain_right.n149 a_n2204_n5888# 0.350239f
C178 drain_right.n150 a_n2204_n5888# 0.035452f
C179 drain_right.n151 a_n2204_n5888# 0.025716f
C180 drain_right.n152 a_n2204_n5888# 0.013819f
C181 drain_right.n153 a_n2204_n5888# 0.032662f
C182 drain_right.n154 a_n2204_n5888# 0.014631f
C183 drain_right.n155 a_n2204_n5888# 0.025716f
C184 drain_right.n156 a_n2204_n5888# 0.013819f
C185 drain_right.n157 a_n2204_n5888# 0.032662f
C186 drain_right.n158 a_n2204_n5888# 0.014631f
C187 drain_right.n159 a_n2204_n5888# 0.025716f
C188 drain_right.n160 a_n2204_n5888# 0.013819f
C189 drain_right.n161 a_n2204_n5888# 0.032662f
C190 drain_right.n162 a_n2204_n5888# 0.014631f
C191 drain_right.n163 a_n2204_n5888# 0.025716f
C192 drain_right.n164 a_n2204_n5888# 0.013819f
C193 drain_right.n165 a_n2204_n5888# 0.032662f
C194 drain_right.n166 a_n2204_n5888# 0.032662f
C195 drain_right.n167 a_n2204_n5888# 0.014631f
C196 drain_right.n168 a_n2204_n5888# 0.025716f
C197 drain_right.n169 a_n2204_n5888# 0.013819f
C198 drain_right.n170 a_n2204_n5888# 0.032662f
C199 drain_right.n171 a_n2204_n5888# 0.014631f
C200 drain_right.n172 a_n2204_n5888# 0.025716f
C201 drain_right.n173 a_n2204_n5888# 0.013819f
C202 drain_right.n174 a_n2204_n5888# 0.032662f
C203 drain_right.n175 a_n2204_n5888# 0.014631f
C204 drain_right.n176 a_n2204_n5888# 0.025716f
C205 drain_right.n177 a_n2204_n5888# 0.013819f
C206 drain_right.n178 a_n2204_n5888# 0.032662f
C207 drain_right.n179 a_n2204_n5888# 0.014631f
C208 drain_right.n180 a_n2204_n5888# 0.025716f
C209 drain_right.n181 a_n2204_n5888# 0.013819f
C210 drain_right.n182 a_n2204_n5888# 0.032662f
C211 drain_right.n183 a_n2204_n5888# 0.014631f
C212 drain_right.n184 a_n2204_n5888# 0.025716f
C213 drain_right.n185 a_n2204_n5888# 0.014225f
C214 drain_right.n186 a_n2204_n5888# 0.032662f
C215 drain_right.n187 a_n2204_n5888# 0.013819f
C216 drain_right.n188 a_n2204_n5888# 0.014631f
C217 drain_right.n189 a_n2204_n5888# 0.025716f
C218 drain_right.n190 a_n2204_n5888# 0.013819f
C219 drain_right.n191 a_n2204_n5888# 0.032662f
C220 drain_right.n192 a_n2204_n5888# 0.014631f
C221 drain_right.n193 a_n2204_n5888# 0.025716f
C222 drain_right.n194 a_n2204_n5888# 0.013819f
C223 drain_right.n195 a_n2204_n5888# 0.024497f
C224 drain_right.n196 a_n2204_n5888# 0.02309f
C225 drain_right.t9 a_n2204_n5888# 0.056965f
C226 drain_right.n197 a_n2204_n5888# 0.313756f
C227 drain_right.n198 a_n2204_n5888# 2.78428f
C228 drain_right.n199 a_n2204_n5888# 0.013819f
C229 drain_right.n200 a_n2204_n5888# 0.014631f
C230 drain_right.n201 a_n2204_n5888# 0.032662f
C231 drain_right.n202 a_n2204_n5888# 0.032662f
C232 drain_right.n203 a_n2204_n5888# 0.014631f
C233 drain_right.n204 a_n2204_n5888# 0.013819f
C234 drain_right.n205 a_n2204_n5888# 0.025716f
C235 drain_right.n206 a_n2204_n5888# 0.025716f
C236 drain_right.n207 a_n2204_n5888# 0.013819f
C237 drain_right.n208 a_n2204_n5888# 0.014631f
C238 drain_right.n209 a_n2204_n5888# 0.032662f
C239 drain_right.n210 a_n2204_n5888# 0.032662f
C240 drain_right.n211 a_n2204_n5888# 0.014631f
C241 drain_right.n212 a_n2204_n5888# 0.013819f
C242 drain_right.n213 a_n2204_n5888# 0.025716f
C243 drain_right.n214 a_n2204_n5888# 0.025716f
C244 drain_right.n215 a_n2204_n5888# 0.013819f
C245 drain_right.n216 a_n2204_n5888# 0.014631f
C246 drain_right.n217 a_n2204_n5888# 0.032662f
C247 drain_right.n218 a_n2204_n5888# 0.032662f
C248 drain_right.n219 a_n2204_n5888# 0.032662f
C249 drain_right.n220 a_n2204_n5888# 0.014225f
C250 drain_right.n221 a_n2204_n5888# 0.013819f
C251 drain_right.n222 a_n2204_n5888# 0.025716f
C252 drain_right.n223 a_n2204_n5888# 0.025716f
C253 drain_right.n224 a_n2204_n5888# 0.013819f
C254 drain_right.n225 a_n2204_n5888# 0.014631f
C255 drain_right.n226 a_n2204_n5888# 0.032662f
C256 drain_right.n227 a_n2204_n5888# 0.032662f
C257 drain_right.n228 a_n2204_n5888# 0.014631f
C258 drain_right.n229 a_n2204_n5888# 0.013819f
C259 drain_right.n230 a_n2204_n5888# 0.025716f
C260 drain_right.n231 a_n2204_n5888# 0.025716f
C261 drain_right.n232 a_n2204_n5888# 0.013819f
C262 drain_right.n233 a_n2204_n5888# 0.014631f
C263 drain_right.n234 a_n2204_n5888# 0.032662f
C264 drain_right.n235 a_n2204_n5888# 0.032662f
C265 drain_right.n236 a_n2204_n5888# 0.014631f
C266 drain_right.n237 a_n2204_n5888# 0.013819f
C267 drain_right.n238 a_n2204_n5888# 0.025716f
C268 drain_right.n239 a_n2204_n5888# 0.025716f
C269 drain_right.n240 a_n2204_n5888# 0.013819f
C270 drain_right.n241 a_n2204_n5888# 0.014631f
C271 drain_right.n242 a_n2204_n5888# 0.032662f
C272 drain_right.n243 a_n2204_n5888# 0.032662f
C273 drain_right.n244 a_n2204_n5888# 0.014631f
C274 drain_right.n245 a_n2204_n5888# 0.013819f
C275 drain_right.n246 a_n2204_n5888# 0.025716f
C276 drain_right.n247 a_n2204_n5888# 0.025716f
C277 drain_right.n248 a_n2204_n5888# 0.013819f
C278 drain_right.n249 a_n2204_n5888# 0.014631f
C279 drain_right.n250 a_n2204_n5888# 0.032662f
C280 drain_right.n251 a_n2204_n5888# 0.032662f
C281 drain_right.n252 a_n2204_n5888# 0.014631f
C282 drain_right.n253 a_n2204_n5888# 0.013819f
C283 drain_right.n254 a_n2204_n5888# 0.025716f
C284 drain_right.n255 a_n2204_n5888# 0.025716f
C285 drain_right.n256 a_n2204_n5888# 0.013819f
C286 drain_right.n257 a_n2204_n5888# 0.014631f
C287 drain_right.n258 a_n2204_n5888# 0.032662f
C288 drain_right.n259 a_n2204_n5888# 0.032662f
C289 drain_right.n260 a_n2204_n5888# 0.014631f
C290 drain_right.n261 a_n2204_n5888# 0.013819f
C291 drain_right.n262 a_n2204_n5888# 0.025716f
C292 drain_right.n263 a_n2204_n5888# 0.025716f
C293 drain_right.n264 a_n2204_n5888# 0.013819f
C294 drain_right.n265 a_n2204_n5888# 0.014225f
C295 drain_right.n266 a_n2204_n5888# 0.014225f
C296 drain_right.n267 a_n2204_n5888# 0.032662f
C297 drain_right.n268 a_n2204_n5888# 0.032662f
C298 drain_right.n269 a_n2204_n5888# 0.014631f
C299 drain_right.n270 a_n2204_n5888# 0.013819f
C300 drain_right.n271 a_n2204_n5888# 0.025716f
C301 drain_right.n272 a_n2204_n5888# 0.025716f
C302 drain_right.n273 a_n2204_n5888# 0.013819f
C303 drain_right.n274 a_n2204_n5888# 0.014631f
C304 drain_right.n275 a_n2204_n5888# 0.032662f
C305 drain_right.n276 a_n2204_n5888# 0.032662f
C306 drain_right.n277 a_n2204_n5888# 0.014631f
C307 drain_right.n278 a_n2204_n5888# 0.013819f
C308 drain_right.n279 a_n2204_n5888# 0.025716f
C309 drain_right.n280 a_n2204_n5888# 0.025716f
C310 drain_right.n281 a_n2204_n5888# 0.013819f
C311 drain_right.n282 a_n2204_n5888# 0.014631f
C312 drain_right.n283 a_n2204_n5888# 0.032662f
C313 drain_right.n284 a_n2204_n5888# 0.069481f
C314 drain_right.n285 a_n2204_n5888# 0.014631f
C315 drain_right.n286 a_n2204_n5888# 0.013819f
C316 drain_right.n287 a_n2204_n5888# 0.056631f
C317 drain_right.n288 a_n2204_n5888# 0.056443f
C318 drain_right.n289 a_n2204_n5888# 0.345275f
C319 minus.n0 a_n2204_n5888# 0.042927f
C320 minus.n1 a_n2204_n5888# 0.009741f
C321 minus.t5 a_n2204_n5888# 1.81969f
C322 minus.n2 a_n2204_n5888# 0.057147f
C323 minus.n3 a_n2204_n5888# 0.009741f
C324 minus.t8 a_n2204_n5888# 1.81969f
C325 minus.t10 a_n2204_n5888# 1.8342f
C326 minus.t9 a_n2204_n5888# 1.81969f
C327 minus.n4 a_n2204_n5888# 0.67352f
C328 minus.n5 a_n2204_n5888# 0.65473f
C329 minus.n6 a_n2204_n5888# 0.17562f
C330 minus.n7 a_n2204_n5888# 0.057281f
C331 minus.n8 a_n2204_n5888# 0.666879f
C332 minus.t7 a_n2204_n5888# 1.81969f
C333 minus.n9 a_n2204_n5888# 0.676091f
C334 minus.t3 a_n2204_n5888# 1.81969f
C335 minus.n10 a_n2204_n5888# 0.666879f
C336 minus.n11 a_n2204_n5888# 0.057281f
C337 minus.n12 a_n2204_n5888# 0.042927f
C338 minus.n13 a_n2204_n5888# 0.042927f
C339 minus.n14 a_n2204_n5888# 0.668203f
C340 minus.n15 a_n2204_n5888# 0.009741f
C341 minus.t4 a_n2204_n5888# 1.81969f
C342 minus.n16 a_n2204_n5888# 0.663968f
C343 minus.n17 a_n2204_n5888# 2.26437f
C344 minus.n18 a_n2204_n5888# 0.042927f
C345 minus.n19 a_n2204_n5888# 0.009741f
C346 minus.n20 a_n2204_n5888# 0.057147f
C347 minus.n21 a_n2204_n5888# 0.009741f
C348 minus.t12 a_n2204_n5888# 1.8342f
C349 minus.t2 a_n2204_n5888# 1.81969f
C350 minus.n22 a_n2204_n5888# 0.67352f
C351 minus.n23 a_n2204_n5888# 0.65473f
C352 minus.n24 a_n2204_n5888# 0.17562f
C353 minus.n25 a_n2204_n5888# 0.057281f
C354 minus.t6 a_n2204_n5888# 1.81969f
C355 minus.n26 a_n2204_n5888# 0.666879f
C356 minus.t13 a_n2204_n5888# 1.81969f
C357 minus.n27 a_n2204_n5888# 0.676091f
C358 minus.t1 a_n2204_n5888# 1.81969f
C359 minus.n28 a_n2204_n5888# 0.666879f
C360 minus.n29 a_n2204_n5888# 0.057281f
C361 minus.n30 a_n2204_n5888# 0.042927f
C362 minus.n31 a_n2204_n5888# 0.042927f
C363 minus.t0 a_n2204_n5888# 1.81969f
C364 minus.n32 a_n2204_n5888# 0.668203f
C365 minus.n33 a_n2204_n5888# 0.009741f
C366 minus.t11 a_n2204_n5888# 1.81969f
C367 minus.n34 a_n2204_n5888# 0.663968f
C368 minus.n35 a_n2204_n5888# 0.288141f
C369 minus.n36 a_n2204_n5888# 2.6634f
C370 source.n0 a_n2204_n5888# 0.036027f
C371 source.n1 a_n2204_n5888# 0.026133f
C372 source.n2 a_n2204_n5888# 0.014043f
C373 source.n3 a_n2204_n5888# 0.033192f
C374 source.n4 a_n2204_n5888# 0.014869f
C375 source.n5 a_n2204_n5888# 0.026133f
C376 source.n6 a_n2204_n5888# 0.014043f
C377 source.n7 a_n2204_n5888# 0.033192f
C378 source.n8 a_n2204_n5888# 0.014869f
C379 source.n9 a_n2204_n5888# 0.026133f
C380 source.n10 a_n2204_n5888# 0.014043f
C381 source.n11 a_n2204_n5888# 0.033192f
C382 source.n12 a_n2204_n5888# 0.014869f
C383 source.n13 a_n2204_n5888# 0.026133f
C384 source.n14 a_n2204_n5888# 0.014043f
C385 source.n15 a_n2204_n5888# 0.033192f
C386 source.n16 a_n2204_n5888# 0.033192f
C387 source.n17 a_n2204_n5888# 0.014869f
C388 source.n18 a_n2204_n5888# 0.026133f
C389 source.n19 a_n2204_n5888# 0.014043f
C390 source.n20 a_n2204_n5888# 0.033192f
C391 source.n21 a_n2204_n5888# 0.014869f
C392 source.n22 a_n2204_n5888# 0.026133f
C393 source.n23 a_n2204_n5888# 0.014043f
C394 source.n24 a_n2204_n5888# 0.033192f
C395 source.n25 a_n2204_n5888# 0.014869f
C396 source.n26 a_n2204_n5888# 0.026133f
C397 source.n27 a_n2204_n5888# 0.014043f
C398 source.n28 a_n2204_n5888# 0.033192f
C399 source.n29 a_n2204_n5888# 0.014869f
C400 source.n30 a_n2204_n5888# 0.026133f
C401 source.n31 a_n2204_n5888# 0.014043f
C402 source.n32 a_n2204_n5888# 0.033192f
C403 source.n33 a_n2204_n5888# 0.014869f
C404 source.n34 a_n2204_n5888# 0.026133f
C405 source.n35 a_n2204_n5888# 0.014456f
C406 source.n36 a_n2204_n5888# 0.033192f
C407 source.n37 a_n2204_n5888# 0.014043f
C408 source.n38 a_n2204_n5888# 0.014869f
C409 source.n39 a_n2204_n5888# 0.026133f
C410 source.n40 a_n2204_n5888# 0.014043f
C411 source.n41 a_n2204_n5888# 0.033192f
C412 source.n42 a_n2204_n5888# 0.014869f
C413 source.n43 a_n2204_n5888# 0.026133f
C414 source.n44 a_n2204_n5888# 0.014043f
C415 source.n45 a_n2204_n5888# 0.024894f
C416 source.n46 a_n2204_n5888# 0.023464f
C417 source.t26 a_n2204_n5888# 0.057889f
C418 source.n47 a_n2204_n5888# 0.318846f
C419 source.n48 a_n2204_n5888# 2.82945f
C420 source.n49 a_n2204_n5888# 0.014043f
C421 source.n50 a_n2204_n5888# 0.014869f
C422 source.n51 a_n2204_n5888# 0.033192f
C423 source.n52 a_n2204_n5888# 0.033192f
C424 source.n53 a_n2204_n5888# 0.014869f
C425 source.n54 a_n2204_n5888# 0.014043f
C426 source.n55 a_n2204_n5888# 0.026133f
C427 source.n56 a_n2204_n5888# 0.026133f
C428 source.n57 a_n2204_n5888# 0.014043f
C429 source.n58 a_n2204_n5888# 0.014869f
C430 source.n59 a_n2204_n5888# 0.033192f
C431 source.n60 a_n2204_n5888# 0.033192f
C432 source.n61 a_n2204_n5888# 0.014869f
C433 source.n62 a_n2204_n5888# 0.014043f
C434 source.n63 a_n2204_n5888# 0.026133f
C435 source.n64 a_n2204_n5888# 0.026133f
C436 source.n65 a_n2204_n5888# 0.014043f
C437 source.n66 a_n2204_n5888# 0.014869f
C438 source.n67 a_n2204_n5888# 0.033192f
C439 source.n68 a_n2204_n5888# 0.033192f
C440 source.n69 a_n2204_n5888# 0.033192f
C441 source.n70 a_n2204_n5888# 0.014456f
C442 source.n71 a_n2204_n5888# 0.014043f
C443 source.n72 a_n2204_n5888# 0.026133f
C444 source.n73 a_n2204_n5888# 0.026133f
C445 source.n74 a_n2204_n5888# 0.014043f
C446 source.n75 a_n2204_n5888# 0.014869f
C447 source.n76 a_n2204_n5888# 0.033192f
C448 source.n77 a_n2204_n5888# 0.033192f
C449 source.n78 a_n2204_n5888# 0.014869f
C450 source.n79 a_n2204_n5888# 0.014043f
C451 source.n80 a_n2204_n5888# 0.026133f
C452 source.n81 a_n2204_n5888# 0.026133f
C453 source.n82 a_n2204_n5888# 0.014043f
C454 source.n83 a_n2204_n5888# 0.014869f
C455 source.n84 a_n2204_n5888# 0.033192f
C456 source.n85 a_n2204_n5888# 0.033192f
C457 source.n86 a_n2204_n5888# 0.014869f
C458 source.n87 a_n2204_n5888# 0.014043f
C459 source.n88 a_n2204_n5888# 0.026133f
C460 source.n89 a_n2204_n5888# 0.026133f
C461 source.n90 a_n2204_n5888# 0.014043f
C462 source.n91 a_n2204_n5888# 0.014869f
C463 source.n92 a_n2204_n5888# 0.033192f
C464 source.n93 a_n2204_n5888# 0.033192f
C465 source.n94 a_n2204_n5888# 0.014869f
C466 source.n95 a_n2204_n5888# 0.014043f
C467 source.n96 a_n2204_n5888# 0.026133f
C468 source.n97 a_n2204_n5888# 0.026133f
C469 source.n98 a_n2204_n5888# 0.014043f
C470 source.n99 a_n2204_n5888# 0.014869f
C471 source.n100 a_n2204_n5888# 0.033192f
C472 source.n101 a_n2204_n5888# 0.033192f
C473 source.n102 a_n2204_n5888# 0.014869f
C474 source.n103 a_n2204_n5888# 0.014043f
C475 source.n104 a_n2204_n5888# 0.026133f
C476 source.n105 a_n2204_n5888# 0.026133f
C477 source.n106 a_n2204_n5888# 0.014043f
C478 source.n107 a_n2204_n5888# 0.014869f
C479 source.n108 a_n2204_n5888# 0.033192f
C480 source.n109 a_n2204_n5888# 0.033192f
C481 source.n110 a_n2204_n5888# 0.014869f
C482 source.n111 a_n2204_n5888# 0.014043f
C483 source.n112 a_n2204_n5888# 0.026133f
C484 source.n113 a_n2204_n5888# 0.026133f
C485 source.n114 a_n2204_n5888# 0.014043f
C486 source.n115 a_n2204_n5888# 0.014456f
C487 source.n116 a_n2204_n5888# 0.014456f
C488 source.n117 a_n2204_n5888# 0.033192f
C489 source.n118 a_n2204_n5888# 0.033192f
C490 source.n119 a_n2204_n5888# 0.014869f
C491 source.n120 a_n2204_n5888# 0.014043f
C492 source.n121 a_n2204_n5888# 0.026133f
C493 source.n122 a_n2204_n5888# 0.026133f
C494 source.n123 a_n2204_n5888# 0.014043f
C495 source.n124 a_n2204_n5888# 0.014869f
C496 source.n125 a_n2204_n5888# 0.033192f
C497 source.n126 a_n2204_n5888# 0.033192f
C498 source.n127 a_n2204_n5888# 0.014869f
C499 source.n128 a_n2204_n5888# 0.014043f
C500 source.n129 a_n2204_n5888# 0.026133f
C501 source.n130 a_n2204_n5888# 0.026133f
C502 source.n131 a_n2204_n5888# 0.014043f
C503 source.n132 a_n2204_n5888# 0.014869f
C504 source.n133 a_n2204_n5888# 0.033192f
C505 source.n134 a_n2204_n5888# 0.070608f
C506 source.n135 a_n2204_n5888# 0.014869f
C507 source.n136 a_n2204_n5888# 0.014043f
C508 source.n137 a_n2204_n5888# 0.057549f
C509 source.n138 a_n2204_n5888# 0.03929f
C510 source.n139 a_n2204_n5888# 2.08758f
C511 source.t22 a_n2204_n5888# 0.51628f
C512 source.t25 a_n2204_n5888# 0.51628f
C513 source.n140 a_n2204_n5888# 4.67241f
C514 source.n141 a_n2204_n5888# 0.406074f
C515 source.t19 a_n2204_n5888# 0.51628f
C516 source.t20 a_n2204_n5888# 0.51628f
C517 source.n142 a_n2204_n5888# 4.67241f
C518 source.n143 a_n2204_n5888# 0.406074f
C519 source.t17 a_n2204_n5888# 0.51628f
C520 source.t18 a_n2204_n5888# 0.51628f
C521 source.n144 a_n2204_n5888# 4.67241f
C522 source.n145 a_n2204_n5888# 0.411881f
C523 source.n146 a_n2204_n5888# 0.036027f
C524 source.n147 a_n2204_n5888# 0.026133f
C525 source.n148 a_n2204_n5888# 0.014043f
C526 source.n149 a_n2204_n5888# 0.033192f
C527 source.n150 a_n2204_n5888# 0.014869f
C528 source.n151 a_n2204_n5888# 0.026133f
C529 source.n152 a_n2204_n5888# 0.014043f
C530 source.n153 a_n2204_n5888# 0.033192f
C531 source.n154 a_n2204_n5888# 0.014869f
C532 source.n155 a_n2204_n5888# 0.026133f
C533 source.n156 a_n2204_n5888# 0.014043f
C534 source.n157 a_n2204_n5888# 0.033192f
C535 source.n158 a_n2204_n5888# 0.014869f
C536 source.n159 a_n2204_n5888# 0.026133f
C537 source.n160 a_n2204_n5888# 0.014043f
C538 source.n161 a_n2204_n5888# 0.033192f
C539 source.n162 a_n2204_n5888# 0.033192f
C540 source.n163 a_n2204_n5888# 0.014869f
C541 source.n164 a_n2204_n5888# 0.026133f
C542 source.n165 a_n2204_n5888# 0.014043f
C543 source.n166 a_n2204_n5888# 0.033192f
C544 source.n167 a_n2204_n5888# 0.014869f
C545 source.n168 a_n2204_n5888# 0.026133f
C546 source.n169 a_n2204_n5888# 0.014043f
C547 source.n170 a_n2204_n5888# 0.033192f
C548 source.n171 a_n2204_n5888# 0.014869f
C549 source.n172 a_n2204_n5888# 0.026133f
C550 source.n173 a_n2204_n5888# 0.014043f
C551 source.n174 a_n2204_n5888# 0.033192f
C552 source.n175 a_n2204_n5888# 0.014869f
C553 source.n176 a_n2204_n5888# 0.026133f
C554 source.n177 a_n2204_n5888# 0.014043f
C555 source.n178 a_n2204_n5888# 0.033192f
C556 source.n179 a_n2204_n5888# 0.014869f
C557 source.n180 a_n2204_n5888# 0.026133f
C558 source.n181 a_n2204_n5888# 0.014456f
C559 source.n182 a_n2204_n5888# 0.033192f
C560 source.n183 a_n2204_n5888# 0.014043f
C561 source.n184 a_n2204_n5888# 0.014869f
C562 source.n185 a_n2204_n5888# 0.026133f
C563 source.n186 a_n2204_n5888# 0.014043f
C564 source.n187 a_n2204_n5888# 0.033192f
C565 source.n188 a_n2204_n5888# 0.014869f
C566 source.n189 a_n2204_n5888# 0.026133f
C567 source.n190 a_n2204_n5888# 0.014043f
C568 source.n191 a_n2204_n5888# 0.024894f
C569 source.n192 a_n2204_n5888# 0.023464f
C570 source.t7 a_n2204_n5888# 0.057889f
C571 source.n193 a_n2204_n5888# 0.318846f
C572 source.n194 a_n2204_n5888# 2.82945f
C573 source.n195 a_n2204_n5888# 0.014043f
C574 source.n196 a_n2204_n5888# 0.014869f
C575 source.n197 a_n2204_n5888# 0.033192f
C576 source.n198 a_n2204_n5888# 0.033192f
C577 source.n199 a_n2204_n5888# 0.014869f
C578 source.n200 a_n2204_n5888# 0.014043f
C579 source.n201 a_n2204_n5888# 0.026133f
C580 source.n202 a_n2204_n5888# 0.026133f
C581 source.n203 a_n2204_n5888# 0.014043f
C582 source.n204 a_n2204_n5888# 0.014869f
C583 source.n205 a_n2204_n5888# 0.033192f
C584 source.n206 a_n2204_n5888# 0.033192f
C585 source.n207 a_n2204_n5888# 0.014869f
C586 source.n208 a_n2204_n5888# 0.014043f
C587 source.n209 a_n2204_n5888# 0.026133f
C588 source.n210 a_n2204_n5888# 0.026133f
C589 source.n211 a_n2204_n5888# 0.014043f
C590 source.n212 a_n2204_n5888# 0.014869f
C591 source.n213 a_n2204_n5888# 0.033192f
C592 source.n214 a_n2204_n5888# 0.033192f
C593 source.n215 a_n2204_n5888# 0.033192f
C594 source.n216 a_n2204_n5888# 0.014456f
C595 source.n217 a_n2204_n5888# 0.014043f
C596 source.n218 a_n2204_n5888# 0.026133f
C597 source.n219 a_n2204_n5888# 0.026133f
C598 source.n220 a_n2204_n5888# 0.014043f
C599 source.n221 a_n2204_n5888# 0.014869f
C600 source.n222 a_n2204_n5888# 0.033192f
C601 source.n223 a_n2204_n5888# 0.033192f
C602 source.n224 a_n2204_n5888# 0.014869f
C603 source.n225 a_n2204_n5888# 0.014043f
C604 source.n226 a_n2204_n5888# 0.026133f
C605 source.n227 a_n2204_n5888# 0.026133f
C606 source.n228 a_n2204_n5888# 0.014043f
C607 source.n229 a_n2204_n5888# 0.014869f
C608 source.n230 a_n2204_n5888# 0.033192f
C609 source.n231 a_n2204_n5888# 0.033192f
C610 source.n232 a_n2204_n5888# 0.014869f
C611 source.n233 a_n2204_n5888# 0.014043f
C612 source.n234 a_n2204_n5888# 0.026133f
C613 source.n235 a_n2204_n5888# 0.026133f
C614 source.n236 a_n2204_n5888# 0.014043f
C615 source.n237 a_n2204_n5888# 0.014869f
C616 source.n238 a_n2204_n5888# 0.033192f
C617 source.n239 a_n2204_n5888# 0.033192f
C618 source.n240 a_n2204_n5888# 0.014869f
C619 source.n241 a_n2204_n5888# 0.014043f
C620 source.n242 a_n2204_n5888# 0.026133f
C621 source.n243 a_n2204_n5888# 0.026133f
C622 source.n244 a_n2204_n5888# 0.014043f
C623 source.n245 a_n2204_n5888# 0.014869f
C624 source.n246 a_n2204_n5888# 0.033192f
C625 source.n247 a_n2204_n5888# 0.033192f
C626 source.n248 a_n2204_n5888# 0.014869f
C627 source.n249 a_n2204_n5888# 0.014043f
C628 source.n250 a_n2204_n5888# 0.026133f
C629 source.n251 a_n2204_n5888# 0.026133f
C630 source.n252 a_n2204_n5888# 0.014043f
C631 source.n253 a_n2204_n5888# 0.014869f
C632 source.n254 a_n2204_n5888# 0.033192f
C633 source.n255 a_n2204_n5888# 0.033192f
C634 source.n256 a_n2204_n5888# 0.014869f
C635 source.n257 a_n2204_n5888# 0.014043f
C636 source.n258 a_n2204_n5888# 0.026133f
C637 source.n259 a_n2204_n5888# 0.026133f
C638 source.n260 a_n2204_n5888# 0.014043f
C639 source.n261 a_n2204_n5888# 0.014456f
C640 source.n262 a_n2204_n5888# 0.014456f
C641 source.n263 a_n2204_n5888# 0.033192f
C642 source.n264 a_n2204_n5888# 0.033192f
C643 source.n265 a_n2204_n5888# 0.014869f
C644 source.n266 a_n2204_n5888# 0.014043f
C645 source.n267 a_n2204_n5888# 0.026133f
C646 source.n268 a_n2204_n5888# 0.026133f
C647 source.n269 a_n2204_n5888# 0.014043f
C648 source.n270 a_n2204_n5888# 0.014869f
C649 source.n271 a_n2204_n5888# 0.033192f
C650 source.n272 a_n2204_n5888# 0.033192f
C651 source.n273 a_n2204_n5888# 0.014869f
C652 source.n274 a_n2204_n5888# 0.014043f
C653 source.n275 a_n2204_n5888# 0.026133f
C654 source.n276 a_n2204_n5888# 0.026133f
C655 source.n277 a_n2204_n5888# 0.014043f
C656 source.n278 a_n2204_n5888# 0.014869f
C657 source.n279 a_n2204_n5888# 0.033192f
C658 source.n280 a_n2204_n5888# 0.070608f
C659 source.n281 a_n2204_n5888# 0.014869f
C660 source.n282 a_n2204_n5888# 0.014043f
C661 source.n283 a_n2204_n5888# 0.057549f
C662 source.n284 a_n2204_n5888# 0.03929f
C663 source.n285 a_n2204_n5888# 0.161538f
C664 source.t11 a_n2204_n5888# 0.51628f
C665 source.t4 a_n2204_n5888# 0.51628f
C666 source.n286 a_n2204_n5888# 4.67241f
C667 source.n287 a_n2204_n5888# 0.406074f
C668 source.t12 a_n2204_n5888# 0.51628f
C669 source.t8 a_n2204_n5888# 0.51628f
C670 source.n288 a_n2204_n5888# 4.67241f
C671 source.n289 a_n2204_n5888# 0.406074f
C672 source.t1 a_n2204_n5888# 0.51628f
C673 source.t2 a_n2204_n5888# 0.51628f
C674 source.n290 a_n2204_n5888# 4.67241f
C675 source.n291 a_n2204_n5888# 2.89872f
C676 source.t15 a_n2204_n5888# 0.51628f
C677 source.t23 a_n2204_n5888# 0.51628f
C678 source.n292 a_n2204_n5888# 4.67241f
C679 source.n293 a_n2204_n5888# 2.89873f
C680 source.t24 a_n2204_n5888# 0.51628f
C681 source.t27 a_n2204_n5888# 0.51628f
C682 source.n294 a_n2204_n5888# 4.67241f
C683 source.n295 a_n2204_n5888# 0.406076f
C684 source.t16 a_n2204_n5888# 0.51628f
C685 source.t21 a_n2204_n5888# 0.51628f
C686 source.n296 a_n2204_n5888# 4.67241f
C687 source.n297 a_n2204_n5888# 0.406076f
C688 source.n298 a_n2204_n5888# 0.036027f
C689 source.n299 a_n2204_n5888# 0.026133f
C690 source.n300 a_n2204_n5888# 0.014043f
C691 source.n301 a_n2204_n5888# 0.033192f
C692 source.n302 a_n2204_n5888# 0.014869f
C693 source.n303 a_n2204_n5888# 0.026133f
C694 source.n304 a_n2204_n5888# 0.014043f
C695 source.n305 a_n2204_n5888# 0.033192f
C696 source.n306 a_n2204_n5888# 0.014869f
C697 source.n307 a_n2204_n5888# 0.026133f
C698 source.n308 a_n2204_n5888# 0.014043f
C699 source.n309 a_n2204_n5888# 0.033192f
C700 source.n310 a_n2204_n5888# 0.014869f
C701 source.n311 a_n2204_n5888# 0.026133f
C702 source.n312 a_n2204_n5888# 0.014043f
C703 source.n313 a_n2204_n5888# 0.033192f
C704 source.n314 a_n2204_n5888# 0.014869f
C705 source.n315 a_n2204_n5888# 0.026133f
C706 source.n316 a_n2204_n5888# 0.014043f
C707 source.n317 a_n2204_n5888# 0.033192f
C708 source.n318 a_n2204_n5888# 0.014869f
C709 source.n319 a_n2204_n5888# 0.026133f
C710 source.n320 a_n2204_n5888# 0.014043f
C711 source.n321 a_n2204_n5888# 0.033192f
C712 source.n322 a_n2204_n5888# 0.014869f
C713 source.n323 a_n2204_n5888# 0.026133f
C714 source.n324 a_n2204_n5888# 0.014043f
C715 source.n325 a_n2204_n5888# 0.033192f
C716 source.n326 a_n2204_n5888# 0.014869f
C717 source.n327 a_n2204_n5888# 0.026133f
C718 source.n328 a_n2204_n5888# 0.014043f
C719 source.n329 a_n2204_n5888# 0.033192f
C720 source.n330 a_n2204_n5888# 0.014869f
C721 source.n331 a_n2204_n5888# 0.026133f
C722 source.n332 a_n2204_n5888# 0.014456f
C723 source.n333 a_n2204_n5888# 0.033192f
C724 source.n334 a_n2204_n5888# 0.014869f
C725 source.n335 a_n2204_n5888# 0.026133f
C726 source.n336 a_n2204_n5888# 0.014043f
C727 source.n337 a_n2204_n5888# 0.033192f
C728 source.n338 a_n2204_n5888# 0.014869f
C729 source.n339 a_n2204_n5888# 0.026133f
C730 source.n340 a_n2204_n5888# 0.014043f
C731 source.n341 a_n2204_n5888# 0.024894f
C732 source.n342 a_n2204_n5888# 0.023464f
C733 source.t14 a_n2204_n5888# 0.057889f
C734 source.n343 a_n2204_n5888# 0.318846f
C735 source.n344 a_n2204_n5888# 2.82945f
C736 source.n345 a_n2204_n5888# 0.014043f
C737 source.n346 a_n2204_n5888# 0.014869f
C738 source.n347 a_n2204_n5888# 0.033192f
C739 source.n348 a_n2204_n5888# 0.033192f
C740 source.n349 a_n2204_n5888# 0.014869f
C741 source.n350 a_n2204_n5888# 0.014043f
C742 source.n351 a_n2204_n5888# 0.026133f
C743 source.n352 a_n2204_n5888# 0.026133f
C744 source.n353 a_n2204_n5888# 0.014043f
C745 source.n354 a_n2204_n5888# 0.014869f
C746 source.n355 a_n2204_n5888# 0.033192f
C747 source.n356 a_n2204_n5888# 0.033192f
C748 source.n357 a_n2204_n5888# 0.014869f
C749 source.n358 a_n2204_n5888# 0.014043f
C750 source.n359 a_n2204_n5888# 0.026133f
C751 source.n360 a_n2204_n5888# 0.026133f
C752 source.n361 a_n2204_n5888# 0.014043f
C753 source.n362 a_n2204_n5888# 0.014043f
C754 source.n363 a_n2204_n5888# 0.014869f
C755 source.n364 a_n2204_n5888# 0.033192f
C756 source.n365 a_n2204_n5888# 0.033192f
C757 source.n366 a_n2204_n5888# 0.033192f
C758 source.n367 a_n2204_n5888# 0.014456f
C759 source.n368 a_n2204_n5888# 0.014043f
C760 source.n369 a_n2204_n5888# 0.026133f
C761 source.n370 a_n2204_n5888# 0.026133f
C762 source.n371 a_n2204_n5888# 0.014043f
C763 source.n372 a_n2204_n5888# 0.014869f
C764 source.n373 a_n2204_n5888# 0.033192f
C765 source.n374 a_n2204_n5888# 0.033192f
C766 source.n375 a_n2204_n5888# 0.014869f
C767 source.n376 a_n2204_n5888# 0.014043f
C768 source.n377 a_n2204_n5888# 0.026133f
C769 source.n378 a_n2204_n5888# 0.026133f
C770 source.n379 a_n2204_n5888# 0.014043f
C771 source.n380 a_n2204_n5888# 0.014869f
C772 source.n381 a_n2204_n5888# 0.033192f
C773 source.n382 a_n2204_n5888# 0.033192f
C774 source.n383 a_n2204_n5888# 0.014869f
C775 source.n384 a_n2204_n5888# 0.014043f
C776 source.n385 a_n2204_n5888# 0.026133f
C777 source.n386 a_n2204_n5888# 0.026133f
C778 source.n387 a_n2204_n5888# 0.014043f
C779 source.n388 a_n2204_n5888# 0.014869f
C780 source.n389 a_n2204_n5888# 0.033192f
C781 source.n390 a_n2204_n5888# 0.033192f
C782 source.n391 a_n2204_n5888# 0.014869f
C783 source.n392 a_n2204_n5888# 0.014043f
C784 source.n393 a_n2204_n5888# 0.026133f
C785 source.n394 a_n2204_n5888# 0.026133f
C786 source.n395 a_n2204_n5888# 0.014043f
C787 source.n396 a_n2204_n5888# 0.014869f
C788 source.n397 a_n2204_n5888# 0.033192f
C789 source.n398 a_n2204_n5888# 0.033192f
C790 source.n399 a_n2204_n5888# 0.014869f
C791 source.n400 a_n2204_n5888# 0.014043f
C792 source.n401 a_n2204_n5888# 0.026133f
C793 source.n402 a_n2204_n5888# 0.026133f
C794 source.n403 a_n2204_n5888# 0.014043f
C795 source.n404 a_n2204_n5888# 0.014869f
C796 source.n405 a_n2204_n5888# 0.033192f
C797 source.n406 a_n2204_n5888# 0.033192f
C798 source.n407 a_n2204_n5888# 0.033192f
C799 source.n408 a_n2204_n5888# 0.014869f
C800 source.n409 a_n2204_n5888# 0.014043f
C801 source.n410 a_n2204_n5888# 0.026133f
C802 source.n411 a_n2204_n5888# 0.026133f
C803 source.n412 a_n2204_n5888# 0.014043f
C804 source.n413 a_n2204_n5888# 0.014456f
C805 source.n414 a_n2204_n5888# 0.014456f
C806 source.n415 a_n2204_n5888# 0.033192f
C807 source.n416 a_n2204_n5888# 0.033192f
C808 source.n417 a_n2204_n5888# 0.014869f
C809 source.n418 a_n2204_n5888# 0.014043f
C810 source.n419 a_n2204_n5888# 0.026133f
C811 source.n420 a_n2204_n5888# 0.026133f
C812 source.n421 a_n2204_n5888# 0.014043f
C813 source.n422 a_n2204_n5888# 0.014869f
C814 source.n423 a_n2204_n5888# 0.033192f
C815 source.n424 a_n2204_n5888# 0.033192f
C816 source.n425 a_n2204_n5888# 0.014869f
C817 source.n426 a_n2204_n5888# 0.014043f
C818 source.n427 a_n2204_n5888# 0.026133f
C819 source.n428 a_n2204_n5888# 0.026133f
C820 source.n429 a_n2204_n5888# 0.014043f
C821 source.n430 a_n2204_n5888# 0.014869f
C822 source.n431 a_n2204_n5888# 0.033192f
C823 source.n432 a_n2204_n5888# 0.070608f
C824 source.n433 a_n2204_n5888# 0.014869f
C825 source.n434 a_n2204_n5888# 0.014043f
C826 source.n435 a_n2204_n5888# 0.057549f
C827 source.n436 a_n2204_n5888# 0.03929f
C828 source.n437 a_n2204_n5888# 0.161538f
C829 source.t13 a_n2204_n5888# 0.51628f
C830 source.t9 a_n2204_n5888# 0.51628f
C831 source.n438 a_n2204_n5888# 4.67241f
C832 source.n439 a_n2204_n5888# 0.411883f
C833 source.t3 a_n2204_n5888# 0.51628f
C834 source.t5 a_n2204_n5888# 0.51628f
C835 source.n440 a_n2204_n5888# 4.67241f
C836 source.n441 a_n2204_n5888# 0.406076f
C837 source.t0 a_n2204_n5888# 0.51628f
C838 source.t10 a_n2204_n5888# 0.51628f
C839 source.n442 a_n2204_n5888# 4.67241f
C840 source.n443 a_n2204_n5888# 0.406076f
C841 source.n444 a_n2204_n5888# 0.036027f
C842 source.n445 a_n2204_n5888# 0.026133f
C843 source.n446 a_n2204_n5888# 0.014043f
C844 source.n447 a_n2204_n5888# 0.033192f
C845 source.n448 a_n2204_n5888# 0.014869f
C846 source.n449 a_n2204_n5888# 0.026133f
C847 source.n450 a_n2204_n5888# 0.014043f
C848 source.n451 a_n2204_n5888# 0.033192f
C849 source.n452 a_n2204_n5888# 0.014869f
C850 source.n453 a_n2204_n5888# 0.026133f
C851 source.n454 a_n2204_n5888# 0.014043f
C852 source.n455 a_n2204_n5888# 0.033192f
C853 source.n456 a_n2204_n5888# 0.014869f
C854 source.n457 a_n2204_n5888# 0.026133f
C855 source.n458 a_n2204_n5888# 0.014043f
C856 source.n459 a_n2204_n5888# 0.033192f
C857 source.n460 a_n2204_n5888# 0.014869f
C858 source.n461 a_n2204_n5888# 0.026133f
C859 source.n462 a_n2204_n5888# 0.014043f
C860 source.n463 a_n2204_n5888# 0.033192f
C861 source.n464 a_n2204_n5888# 0.014869f
C862 source.n465 a_n2204_n5888# 0.026133f
C863 source.n466 a_n2204_n5888# 0.014043f
C864 source.n467 a_n2204_n5888# 0.033192f
C865 source.n468 a_n2204_n5888# 0.014869f
C866 source.n469 a_n2204_n5888# 0.026133f
C867 source.n470 a_n2204_n5888# 0.014043f
C868 source.n471 a_n2204_n5888# 0.033192f
C869 source.n472 a_n2204_n5888# 0.014869f
C870 source.n473 a_n2204_n5888# 0.026133f
C871 source.n474 a_n2204_n5888# 0.014043f
C872 source.n475 a_n2204_n5888# 0.033192f
C873 source.n476 a_n2204_n5888# 0.014869f
C874 source.n477 a_n2204_n5888# 0.026133f
C875 source.n478 a_n2204_n5888# 0.014456f
C876 source.n479 a_n2204_n5888# 0.033192f
C877 source.n480 a_n2204_n5888# 0.014869f
C878 source.n481 a_n2204_n5888# 0.026133f
C879 source.n482 a_n2204_n5888# 0.014043f
C880 source.n483 a_n2204_n5888# 0.033192f
C881 source.n484 a_n2204_n5888# 0.014869f
C882 source.n485 a_n2204_n5888# 0.026133f
C883 source.n486 a_n2204_n5888# 0.014043f
C884 source.n487 a_n2204_n5888# 0.024894f
C885 source.n488 a_n2204_n5888# 0.023464f
C886 source.t6 a_n2204_n5888# 0.057889f
C887 source.n489 a_n2204_n5888# 0.318846f
C888 source.n490 a_n2204_n5888# 2.82945f
C889 source.n491 a_n2204_n5888# 0.014043f
C890 source.n492 a_n2204_n5888# 0.014869f
C891 source.n493 a_n2204_n5888# 0.033192f
C892 source.n494 a_n2204_n5888# 0.033192f
C893 source.n495 a_n2204_n5888# 0.014869f
C894 source.n496 a_n2204_n5888# 0.014043f
C895 source.n497 a_n2204_n5888# 0.026133f
C896 source.n498 a_n2204_n5888# 0.026133f
C897 source.n499 a_n2204_n5888# 0.014043f
C898 source.n500 a_n2204_n5888# 0.014869f
C899 source.n501 a_n2204_n5888# 0.033192f
C900 source.n502 a_n2204_n5888# 0.033192f
C901 source.n503 a_n2204_n5888# 0.014869f
C902 source.n504 a_n2204_n5888# 0.014043f
C903 source.n505 a_n2204_n5888# 0.026133f
C904 source.n506 a_n2204_n5888# 0.026133f
C905 source.n507 a_n2204_n5888# 0.014043f
C906 source.n508 a_n2204_n5888# 0.014043f
C907 source.n509 a_n2204_n5888# 0.014869f
C908 source.n510 a_n2204_n5888# 0.033192f
C909 source.n511 a_n2204_n5888# 0.033192f
C910 source.n512 a_n2204_n5888# 0.033192f
C911 source.n513 a_n2204_n5888# 0.014456f
C912 source.n514 a_n2204_n5888# 0.014043f
C913 source.n515 a_n2204_n5888# 0.026133f
C914 source.n516 a_n2204_n5888# 0.026133f
C915 source.n517 a_n2204_n5888# 0.014043f
C916 source.n518 a_n2204_n5888# 0.014869f
C917 source.n519 a_n2204_n5888# 0.033192f
C918 source.n520 a_n2204_n5888# 0.033192f
C919 source.n521 a_n2204_n5888# 0.014869f
C920 source.n522 a_n2204_n5888# 0.014043f
C921 source.n523 a_n2204_n5888# 0.026133f
C922 source.n524 a_n2204_n5888# 0.026133f
C923 source.n525 a_n2204_n5888# 0.014043f
C924 source.n526 a_n2204_n5888# 0.014869f
C925 source.n527 a_n2204_n5888# 0.033192f
C926 source.n528 a_n2204_n5888# 0.033192f
C927 source.n529 a_n2204_n5888# 0.014869f
C928 source.n530 a_n2204_n5888# 0.014043f
C929 source.n531 a_n2204_n5888# 0.026133f
C930 source.n532 a_n2204_n5888# 0.026133f
C931 source.n533 a_n2204_n5888# 0.014043f
C932 source.n534 a_n2204_n5888# 0.014869f
C933 source.n535 a_n2204_n5888# 0.033192f
C934 source.n536 a_n2204_n5888# 0.033192f
C935 source.n537 a_n2204_n5888# 0.014869f
C936 source.n538 a_n2204_n5888# 0.014043f
C937 source.n539 a_n2204_n5888# 0.026133f
C938 source.n540 a_n2204_n5888# 0.026133f
C939 source.n541 a_n2204_n5888# 0.014043f
C940 source.n542 a_n2204_n5888# 0.014869f
C941 source.n543 a_n2204_n5888# 0.033192f
C942 source.n544 a_n2204_n5888# 0.033192f
C943 source.n545 a_n2204_n5888# 0.014869f
C944 source.n546 a_n2204_n5888# 0.014043f
C945 source.n547 a_n2204_n5888# 0.026133f
C946 source.n548 a_n2204_n5888# 0.026133f
C947 source.n549 a_n2204_n5888# 0.014043f
C948 source.n550 a_n2204_n5888# 0.014869f
C949 source.n551 a_n2204_n5888# 0.033192f
C950 source.n552 a_n2204_n5888# 0.033192f
C951 source.n553 a_n2204_n5888# 0.033192f
C952 source.n554 a_n2204_n5888# 0.014869f
C953 source.n555 a_n2204_n5888# 0.014043f
C954 source.n556 a_n2204_n5888# 0.026133f
C955 source.n557 a_n2204_n5888# 0.026133f
C956 source.n558 a_n2204_n5888# 0.014043f
C957 source.n559 a_n2204_n5888# 0.014456f
C958 source.n560 a_n2204_n5888# 0.014456f
C959 source.n561 a_n2204_n5888# 0.033192f
C960 source.n562 a_n2204_n5888# 0.033192f
C961 source.n563 a_n2204_n5888# 0.014869f
C962 source.n564 a_n2204_n5888# 0.014043f
C963 source.n565 a_n2204_n5888# 0.026133f
C964 source.n566 a_n2204_n5888# 0.026133f
C965 source.n567 a_n2204_n5888# 0.014043f
C966 source.n568 a_n2204_n5888# 0.014869f
C967 source.n569 a_n2204_n5888# 0.033192f
C968 source.n570 a_n2204_n5888# 0.033192f
C969 source.n571 a_n2204_n5888# 0.014869f
C970 source.n572 a_n2204_n5888# 0.014043f
C971 source.n573 a_n2204_n5888# 0.026133f
C972 source.n574 a_n2204_n5888# 0.026133f
C973 source.n575 a_n2204_n5888# 0.014043f
C974 source.n576 a_n2204_n5888# 0.014869f
C975 source.n577 a_n2204_n5888# 0.033192f
C976 source.n578 a_n2204_n5888# 0.070608f
C977 source.n579 a_n2204_n5888# 0.014869f
C978 source.n580 a_n2204_n5888# 0.014043f
C979 source.n581 a_n2204_n5888# 0.057549f
C980 source.n582 a_n2204_n5888# 0.03929f
C981 source.n583 a_n2204_n5888# 0.292562f
C982 source.n584 a_n2204_n5888# 2.80019f
C983 drain_left.n0 a_n2204_n5888# 0.035516f
C984 drain_left.n1 a_n2204_n5888# 0.025762f
C985 drain_left.n2 a_n2204_n5888# 0.013844f
C986 drain_left.n3 a_n2204_n5888# 0.032721f
C987 drain_left.n4 a_n2204_n5888# 0.014658f
C988 drain_left.n5 a_n2204_n5888# 0.025762f
C989 drain_left.n6 a_n2204_n5888# 0.013844f
C990 drain_left.n7 a_n2204_n5888# 0.032721f
C991 drain_left.n8 a_n2204_n5888# 0.014658f
C992 drain_left.n9 a_n2204_n5888# 0.025762f
C993 drain_left.n10 a_n2204_n5888# 0.013844f
C994 drain_left.n11 a_n2204_n5888# 0.032721f
C995 drain_left.n12 a_n2204_n5888# 0.014658f
C996 drain_left.n13 a_n2204_n5888# 0.025762f
C997 drain_left.n14 a_n2204_n5888# 0.013844f
C998 drain_left.n15 a_n2204_n5888# 0.032721f
C999 drain_left.n16 a_n2204_n5888# 0.014658f
C1000 drain_left.n17 a_n2204_n5888# 0.025762f
C1001 drain_left.n18 a_n2204_n5888# 0.013844f
C1002 drain_left.n19 a_n2204_n5888# 0.032721f
C1003 drain_left.n20 a_n2204_n5888# 0.014658f
C1004 drain_left.n21 a_n2204_n5888# 0.025762f
C1005 drain_left.n22 a_n2204_n5888# 0.013844f
C1006 drain_left.n23 a_n2204_n5888# 0.032721f
C1007 drain_left.n24 a_n2204_n5888# 0.014658f
C1008 drain_left.n25 a_n2204_n5888# 0.025762f
C1009 drain_left.n26 a_n2204_n5888# 0.013844f
C1010 drain_left.n27 a_n2204_n5888# 0.032721f
C1011 drain_left.n28 a_n2204_n5888# 0.014658f
C1012 drain_left.n29 a_n2204_n5888# 0.025762f
C1013 drain_left.n30 a_n2204_n5888# 0.013844f
C1014 drain_left.n31 a_n2204_n5888# 0.032721f
C1015 drain_left.n32 a_n2204_n5888# 0.014658f
C1016 drain_left.n33 a_n2204_n5888# 0.025762f
C1017 drain_left.n34 a_n2204_n5888# 0.014251f
C1018 drain_left.n35 a_n2204_n5888# 0.032721f
C1019 drain_left.n36 a_n2204_n5888# 0.014658f
C1020 drain_left.n37 a_n2204_n5888# 0.025762f
C1021 drain_left.n38 a_n2204_n5888# 0.013844f
C1022 drain_left.n39 a_n2204_n5888# 0.032721f
C1023 drain_left.n40 a_n2204_n5888# 0.014658f
C1024 drain_left.n41 a_n2204_n5888# 0.025762f
C1025 drain_left.n42 a_n2204_n5888# 0.013844f
C1026 drain_left.n43 a_n2204_n5888# 0.024541f
C1027 drain_left.n44 a_n2204_n5888# 0.023131f
C1028 drain_left.t11 a_n2204_n5888# 0.057067f
C1029 drain_left.n45 a_n2204_n5888# 0.31432f
C1030 drain_left.n46 a_n2204_n5888# 2.78928f
C1031 drain_left.n47 a_n2204_n5888# 0.013844f
C1032 drain_left.n48 a_n2204_n5888# 0.014658f
C1033 drain_left.n49 a_n2204_n5888# 0.032721f
C1034 drain_left.n50 a_n2204_n5888# 0.032721f
C1035 drain_left.n51 a_n2204_n5888# 0.014658f
C1036 drain_left.n52 a_n2204_n5888# 0.013844f
C1037 drain_left.n53 a_n2204_n5888# 0.025762f
C1038 drain_left.n54 a_n2204_n5888# 0.025762f
C1039 drain_left.n55 a_n2204_n5888# 0.013844f
C1040 drain_left.n56 a_n2204_n5888# 0.014658f
C1041 drain_left.n57 a_n2204_n5888# 0.032721f
C1042 drain_left.n58 a_n2204_n5888# 0.032721f
C1043 drain_left.n59 a_n2204_n5888# 0.014658f
C1044 drain_left.n60 a_n2204_n5888# 0.013844f
C1045 drain_left.n61 a_n2204_n5888# 0.025762f
C1046 drain_left.n62 a_n2204_n5888# 0.025762f
C1047 drain_left.n63 a_n2204_n5888# 0.013844f
C1048 drain_left.n64 a_n2204_n5888# 0.013844f
C1049 drain_left.n65 a_n2204_n5888# 0.014658f
C1050 drain_left.n66 a_n2204_n5888# 0.032721f
C1051 drain_left.n67 a_n2204_n5888# 0.032721f
C1052 drain_left.n68 a_n2204_n5888# 0.032721f
C1053 drain_left.n69 a_n2204_n5888# 0.014251f
C1054 drain_left.n70 a_n2204_n5888# 0.013844f
C1055 drain_left.n71 a_n2204_n5888# 0.025762f
C1056 drain_left.n72 a_n2204_n5888# 0.025762f
C1057 drain_left.n73 a_n2204_n5888# 0.013844f
C1058 drain_left.n74 a_n2204_n5888# 0.014658f
C1059 drain_left.n75 a_n2204_n5888# 0.032721f
C1060 drain_left.n76 a_n2204_n5888# 0.032721f
C1061 drain_left.n77 a_n2204_n5888# 0.014658f
C1062 drain_left.n78 a_n2204_n5888# 0.013844f
C1063 drain_left.n79 a_n2204_n5888# 0.025762f
C1064 drain_left.n80 a_n2204_n5888# 0.025762f
C1065 drain_left.n81 a_n2204_n5888# 0.013844f
C1066 drain_left.n82 a_n2204_n5888# 0.014658f
C1067 drain_left.n83 a_n2204_n5888# 0.032721f
C1068 drain_left.n84 a_n2204_n5888# 0.032721f
C1069 drain_left.n85 a_n2204_n5888# 0.014658f
C1070 drain_left.n86 a_n2204_n5888# 0.013844f
C1071 drain_left.n87 a_n2204_n5888# 0.025762f
C1072 drain_left.n88 a_n2204_n5888# 0.025762f
C1073 drain_left.n89 a_n2204_n5888# 0.013844f
C1074 drain_left.n90 a_n2204_n5888# 0.014658f
C1075 drain_left.n91 a_n2204_n5888# 0.032721f
C1076 drain_left.n92 a_n2204_n5888# 0.032721f
C1077 drain_left.n93 a_n2204_n5888# 0.014658f
C1078 drain_left.n94 a_n2204_n5888# 0.013844f
C1079 drain_left.n95 a_n2204_n5888# 0.025762f
C1080 drain_left.n96 a_n2204_n5888# 0.025762f
C1081 drain_left.n97 a_n2204_n5888# 0.013844f
C1082 drain_left.n98 a_n2204_n5888# 0.014658f
C1083 drain_left.n99 a_n2204_n5888# 0.032721f
C1084 drain_left.n100 a_n2204_n5888# 0.032721f
C1085 drain_left.n101 a_n2204_n5888# 0.014658f
C1086 drain_left.n102 a_n2204_n5888# 0.013844f
C1087 drain_left.n103 a_n2204_n5888# 0.025762f
C1088 drain_left.n104 a_n2204_n5888# 0.025762f
C1089 drain_left.n105 a_n2204_n5888# 0.013844f
C1090 drain_left.n106 a_n2204_n5888# 0.014658f
C1091 drain_left.n107 a_n2204_n5888# 0.032721f
C1092 drain_left.n108 a_n2204_n5888# 0.032721f
C1093 drain_left.n109 a_n2204_n5888# 0.032721f
C1094 drain_left.n110 a_n2204_n5888# 0.014658f
C1095 drain_left.n111 a_n2204_n5888# 0.013844f
C1096 drain_left.n112 a_n2204_n5888# 0.025762f
C1097 drain_left.n113 a_n2204_n5888# 0.025762f
C1098 drain_left.n114 a_n2204_n5888# 0.013844f
C1099 drain_left.n115 a_n2204_n5888# 0.014251f
C1100 drain_left.n116 a_n2204_n5888# 0.014251f
C1101 drain_left.n117 a_n2204_n5888# 0.032721f
C1102 drain_left.n118 a_n2204_n5888# 0.032721f
C1103 drain_left.n119 a_n2204_n5888# 0.014658f
C1104 drain_left.n120 a_n2204_n5888# 0.013844f
C1105 drain_left.n121 a_n2204_n5888# 0.025762f
C1106 drain_left.n122 a_n2204_n5888# 0.025762f
C1107 drain_left.n123 a_n2204_n5888# 0.013844f
C1108 drain_left.n124 a_n2204_n5888# 0.014658f
C1109 drain_left.n125 a_n2204_n5888# 0.032721f
C1110 drain_left.n126 a_n2204_n5888# 0.032721f
C1111 drain_left.n127 a_n2204_n5888# 0.014658f
C1112 drain_left.n128 a_n2204_n5888# 0.013844f
C1113 drain_left.n129 a_n2204_n5888# 0.025762f
C1114 drain_left.n130 a_n2204_n5888# 0.025762f
C1115 drain_left.n131 a_n2204_n5888# 0.013844f
C1116 drain_left.n132 a_n2204_n5888# 0.014658f
C1117 drain_left.n133 a_n2204_n5888# 0.032721f
C1118 drain_left.n134 a_n2204_n5888# 0.069606f
C1119 drain_left.n135 a_n2204_n5888# 0.014658f
C1120 drain_left.n136 a_n2204_n5888# 0.013844f
C1121 drain_left.n137 a_n2204_n5888# 0.056733f
C1122 drain_left.n138 a_n2204_n5888# 0.058453f
C1123 drain_left.t3 a_n2204_n5888# 0.508952f
C1124 drain_left.t0 a_n2204_n5888# 0.508952f
C1125 drain_left.n139 a_n2204_n5888# 4.69054f
C1126 drain_left.n140 a_n2204_n5888# 0.443371f
C1127 drain_left.t7 a_n2204_n5888# 0.508952f
C1128 drain_left.t10 a_n2204_n5888# 0.508952f
C1129 drain_left.n141 a_n2204_n5888# 4.6954f
C1130 drain_left.t5 a_n2204_n5888# 0.508952f
C1131 drain_left.t12 a_n2204_n5888# 0.508952f
C1132 drain_left.n142 a_n2204_n5888# 4.69054f
C1133 drain_left.n143 a_n2204_n5888# 0.656858f
C1134 drain_left.n144 a_n2204_n5888# 2.21791f
C1135 drain_left.n145 a_n2204_n5888# 0.035516f
C1136 drain_left.n146 a_n2204_n5888# 0.025762f
C1137 drain_left.n147 a_n2204_n5888# 0.013844f
C1138 drain_left.n148 a_n2204_n5888# 0.032721f
C1139 drain_left.n149 a_n2204_n5888# 0.014658f
C1140 drain_left.n150 a_n2204_n5888# 0.025762f
C1141 drain_left.n151 a_n2204_n5888# 0.013844f
C1142 drain_left.n152 a_n2204_n5888# 0.032721f
C1143 drain_left.n153 a_n2204_n5888# 0.014658f
C1144 drain_left.n154 a_n2204_n5888# 0.025762f
C1145 drain_left.n155 a_n2204_n5888# 0.013844f
C1146 drain_left.n156 a_n2204_n5888# 0.032721f
C1147 drain_left.n157 a_n2204_n5888# 0.014658f
C1148 drain_left.n158 a_n2204_n5888# 0.025762f
C1149 drain_left.n159 a_n2204_n5888# 0.013844f
C1150 drain_left.n160 a_n2204_n5888# 0.032721f
C1151 drain_left.n161 a_n2204_n5888# 0.032721f
C1152 drain_left.n162 a_n2204_n5888# 0.014658f
C1153 drain_left.n163 a_n2204_n5888# 0.025762f
C1154 drain_left.n164 a_n2204_n5888# 0.013844f
C1155 drain_left.n165 a_n2204_n5888# 0.032721f
C1156 drain_left.n166 a_n2204_n5888# 0.014658f
C1157 drain_left.n167 a_n2204_n5888# 0.025762f
C1158 drain_left.n168 a_n2204_n5888# 0.013844f
C1159 drain_left.n169 a_n2204_n5888# 0.032721f
C1160 drain_left.n170 a_n2204_n5888# 0.014658f
C1161 drain_left.n171 a_n2204_n5888# 0.025762f
C1162 drain_left.n172 a_n2204_n5888# 0.013844f
C1163 drain_left.n173 a_n2204_n5888# 0.032721f
C1164 drain_left.n174 a_n2204_n5888# 0.014658f
C1165 drain_left.n175 a_n2204_n5888# 0.025762f
C1166 drain_left.n176 a_n2204_n5888# 0.013844f
C1167 drain_left.n177 a_n2204_n5888# 0.032721f
C1168 drain_left.n178 a_n2204_n5888# 0.014658f
C1169 drain_left.n179 a_n2204_n5888# 0.025762f
C1170 drain_left.n180 a_n2204_n5888# 0.014251f
C1171 drain_left.n181 a_n2204_n5888# 0.032721f
C1172 drain_left.n182 a_n2204_n5888# 0.013844f
C1173 drain_left.n183 a_n2204_n5888# 0.014658f
C1174 drain_left.n184 a_n2204_n5888# 0.025762f
C1175 drain_left.n185 a_n2204_n5888# 0.013844f
C1176 drain_left.n186 a_n2204_n5888# 0.032721f
C1177 drain_left.n187 a_n2204_n5888# 0.014658f
C1178 drain_left.n188 a_n2204_n5888# 0.025762f
C1179 drain_left.n189 a_n2204_n5888# 0.013844f
C1180 drain_left.n190 a_n2204_n5888# 0.024541f
C1181 drain_left.n191 a_n2204_n5888# 0.023131f
C1182 drain_left.t13 a_n2204_n5888# 0.057067f
C1183 drain_left.n192 a_n2204_n5888# 0.31432f
C1184 drain_left.n193 a_n2204_n5888# 2.78928f
C1185 drain_left.n194 a_n2204_n5888# 0.013844f
C1186 drain_left.n195 a_n2204_n5888# 0.014658f
C1187 drain_left.n196 a_n2204_n5888# 0.032721f
C1188 drain_left.n197 a_n2204_n5888# 0.032721f
C1189 drain_left.n198 a_n2204_n5888# 0.014658f
C1190 drain_left.n199 a_n2204_n5888# 0.013844f
C1191 drain_left.n200 a_n2204_n5888# 0.025762f
C1192 drain_left.n201 a_n2204_n5888# 0.025762f
C1193 drain_left.n202 a_n2204_n5888# 0.013844f
C1194 drain_left.n203 a_n2204_n5888# 0.014658f
C1195 drain_left.n204 a_n2204_n5888# 0.032721f
C1196 drain_left.n205 a_n2204_n5888# 0.032721f
C1197 drain_left.n206 a_n2204_n5888# 0.014658f
C1198 drain_left.n207 a_n2204_n5888# 0.013844f
C1199 drain_left.n208 a_n2204_n5888# 0.025762f
C1200 drain_left.n209 a_n2204_n5888# 0.025762f
C1201 drain_left.n210 a_n2204_n5888# 0.013844f
C1202 drain_left.n211 a_n2204_n5888# 0.014658f
C1203 drain_left.n212 a_n2204_n5888# 0.032721f
C1204 drain_left.n213 a_n2204_n5888# 0.032721f
C1205 drain_left.n214 a_n2204_n5888# 0.032721f
C1206 drain_left.n215 a_n2204_n5888# 0.014251f
C1207 drain_left.n216 a_n2204_n5888# 0.013844f
C1208 drain_left.n217 a_n2204_n5888# 0.025762f
C1209 drain_left.n218 a_n2204_n5888# 0.025762f
C1210 drain_left.n219 a_n2204_n5888# 0.013844f
C1211 drain_left.n220 a_n2204_n5888# 0.014658f
C1212 drain_left.n221 a_n2204_n5888# 0.032721f
C1213 drain_left.n222 a_n2204_n5888# 0.032721f
C1214 drain_left.n223 a_n2204_n5888# 0.014658f
C1215 drain_left.n224 a_n2204_n5888# 0.013844f
C1216 drain_left.n225 a_n2204_n5888# 0.025762f
C1217 drain_left.n226 a_n2204_n5888# 0.025762f
C1218 drain_left.n227 a_n2204_n5888# 0.013844f
C1219 drain_left.n228 a_n2204_n5888# 0.014658f
C1220 drain_left.n229 a_n2204_n5888# 0.032721f
C1221 drain_left.n230 a_n2204_n5888# 0.032721f
C1222 drain_left.n231 a_n2204_n5888# 0.014658f
C1223 drain_left.n232 a_n2204_n5888# 0.013844f
C1224 drain_left.n233 a_n2204_n5888# 0.025762f
C1225 drain_left.n234 a_n2204_n5888# 0.025762f
C1226 drain_left.n235 a_n2204_n5888# 0.013844f
C1227 drain_left.n236 a_n2204_n5888# 0.014658f
C1228 drain_left.n237 a_n2204_n5888# 0.032721f
C1229 drain_left.n238 a_n2204_n5888# 0.032721f
C1230 drain_left.n239 a_n2204_n5888# 0.014658f
C1231 drain_left.n240 a_n2204_n5888# 0.013844f
C1232 drain_left.n241 a_n2204_n5888# 0.025762f
C1233 drain_left.n242 a_n2204_n5888# 0.025762f
C1234 drain_left.n243 a_n2204_n5888# 0.013844f
C1235 drain_left.n244 a_n2204_n5888# 0.014658f
C1236 drain_left.n245 a_n2204_n5888# 0.032721f
C1237 drain_left.n246 a_n2204_n5888# 0.032721f
C1238 drain_left.n247 a_n2204_n5888# 0.014658f
C1239 drain_left.n248 a_n2204_n5888# 0.013844f
C1240 drain_left.n249 a_n2204_n5888# 0.025762f
C1241 drain_left.n250 a_n2204_n5888# 0.025762f
C1242 drain_left.n251 a_n2204_n5888# 0.013844f
C1243 drain_left.n252 a_n2204_n5888# 0.014658f
C1244 drain_left.n253 a_n2204_n5888# 0.032721f
C1245 drain_left.n254 a_n2204_n5888# 0.032721f
C1246 drain_left.n255 a_n2204_n5888# 0.014658f
C1247 drain_left.n256 a_n2204_n5888# 0.013844f
C1248 drain_left.n257 a_n2204_n5888# 0.025762f
C1249 drain_left.n258 a_n2204_n5888# 0.025762f
C1250 drain_left.n259 a_n2204_n5888# 0.013844f
C1251 drain_left.n260 a_n2204_n5888# 0.014251f
C1252 drain_left.n261 a_n2204_n5888# 0.014251f
C1253 drain_left.n262 a_n2204_n5888# 0.032721f
C1254 drain_left.n263 a_n2204_n5888# 0.032721f
C1255 drain_left.n264 a_n2204_n5888# 0.014658f
C1256 drain_left.n265 a_n2204_n5888# 0.013844f
C1257 drain_left.n266 a_n2204_n5888# 0.025762f
C1258 drain_left.n267 a_n2204_n5888# 0.025762f
C1259 drain_left.n268 a_n2204_n5888# 0.013844f
C1260 drain_left.n269 a_n2204_n5888# 0.014658f
C1261 drain_left.n270 a_n2204_n5888# 0.032721f
C1262 drain_left.n271 a_n2204_n5888# 0.032721f
C1263 drain_left.n272 a_n2204_n5888# 0.014658f
C1264 drain_left.n273 a_n2204_n5888# 0.013844f
C1265 drain_left.n274 a_n2204_n5888# 0.025762f
C1266 drain_left.n275 a_n2204_n5888# 0.025762f
C1267 drain_left.n276 a_n2204_n5888# 0.013844f
C1268 drain_left.n277 a_n2204_n5888# 0.014658f
C1269 drain_left.n278 a_n2204_n5888# 0.032721f
C1270 drain_left.n279 a_n2204_n5888# 0.069606f
C1271 drain_left.n280 a_n2204_n5888# 0.014658f
C1272 drain_left.n281 a_n2204_n5888# 0.013844f
C1273 drain_left.n282 a_n2204_n5888# 0.056733f
C1274 drain_left.n283 a_n2204_n5888# 0.058453f
C1275 drain_left.t8 a_n2204_n5888# 0.508952f
C1276 drain_left.t9 a_n2204_n5888# 0.508952f
C1277 drain_left.n284 a_n2204_n5888# 4.69054f
C1278 drain_left.n285 a_n2204_n5888# 0.463508f
C1279 drain_left.t6 a_n2204_n5888# 0.508952f
C1280 drain_left.t2 a_n2204_n5888# 0.508952f
C1281 drain_left.n286 a_n2204_n5888# 4.69054f
C1282 drain_left.n287 a_n2204_n5888# 0.350869f
C1283 drain_left.t1 a_n2204_n5888# 0.508952f
C1284 drain_left.t4 a_n2204_n5888# 0.508952f
C1285 drain_left.n288 a_n2204_n5888# 4.69053f
C1286 drain_left.n289 a_n2204_n5888# 0.575525f
C1287 plus.n0 a_n2204_n5888# 0.043227f
C1288 plus.t1 a_n2204_n5888# 1.83242f
C1289 plus.t2 a_n2204_n5888# 1.83242f
C1290 plus.n1 a_n2204_n5888# 0.043227f
C1291 plus.t5 a_n2204_n5888# 1.83242f
C1292 plus.n2 a_n2204_n5888# 0.671543f
C1293 plus.n3 a_n2204_n5888# 0.057682f
C1294 plus.t7 a_n2204_n5888# 1.83242f
C1295 plus.t8 a_n2204_n5888# 1.83242f
C1296 plus.t9 a_n2204_n5888# 1.83242f
C1297 plus.n4 a_n2204_n5888# 0.67823f
C1298 plus.t10 a_n2204_n5888# 1.84703f
C1299 plus.n5 a_n2204_n5888# 0.659308f
C1300 plus.n6 a_n2204_n5888# 0.176848f
C1301 plus.n7 a_n2204_n5888# 0.009809f
C1302 plus.n8 a_n2204_n5888# 0.671543f
C1303 plus.n9 a_n2204_n5888# 0.680819f
C1304 plus.n10 a_n2204_n5888# 0.057547f
C1305 plus.n11 a_n2204_n5888# 0.057682f
C1306 plus.n12 a_n2204_n5888# 0.043227f
C1307 plus.n13 a_n2204_n5888# 0.009809f
C1308 plus.n14 a_n2204_n5888# 0.672876f
C1309 plus.n15 a_n2204_n5888# 0.009809f
C1310 plus.n16 a_n2204_n5888# 0.668611f
C1311 plus.n17 a_n2204_n5888# 0.778859f
C1312 plus.n18 a_n2204_n5888# 0.043227f
C1313 plus.t12 a_n2204_n5888# 1.83242f
C1314 plus.n19 a_n2204_n5888# 0.043227f
C1315 plus.t4 a_n2204_n5888# 1.83242f
C1316 plus.t3 a_n2204_n5888# 1.83242f
C1317 plus.n20 a_n2204_n5888# 0.671543f
C1318 plus.n21 a_n2204_n5888# 0.057682f
C1319 plus.t0 a_n2204_n5888# 1.83242f
C1320 plus.t11 a_n2204_n5888# 1.83242f
C1321 plus.t6 a_n2204_n5888# 1.83242f
C1322 plus.n22 a_n2204_n5888# 0.67823f
C1323 plus.t13 a_n2204_n5888# 1.84703f
C1324 plus.n23 a_n2204_n5888# 0.659308f
C1325 plus.n24 a_n2204_n5888# 0.176848f
C1326 plus.n25 a_n2204_n5888# 0.009809f
C1327 plus.n26 a_n2204_n5888# 0.671543f
C1328 plus.n27 a_n2204_n5888# 0.680819f
C1329 plus.n28 a_n2204_n5888# 0.057547f
C1330 plus.n29 a_n2204_n5888# 0.057682f
C1331 plus.n30 a_n2204_n5888# 0.043227f
C1332 plus.n31 a_n2204_n5888# 0.009809f
C1333 plus.n32 a_n2204_n5888# 0.672876f
C1334 plus.n33 a_n2204_n5888# 0.009809f
C1335 plus.n34 a_n2204_n5888# 0.668611f
C1336 plus.n35 a_n2204_n5888# 1.75679f
.ends

