* NGSPICE file created from diffpair672.ext - technology: sky130A

.subckt diffpair672 minus drain_right drain_left source plus
X0 drain_right.t5 minus.t0 source.t8 a_n1220_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X1 a_n1220_n5888# a_n1220_n5888# a_n1220_n5888# a_n1220_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=78 ps=406.24 w=25 l=0.3
X2 drain_right.t4 minus.t1 source.t7 a_n1220_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X3 drain_right.t3 minus.t2 source.t6 a_n1220_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X4 drain_left.t5 plus.t0 source.t3 a_n1220_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
X5 a_n1220_n5888# a_n1220_n5888# a_n1220_n5888# a_n1220_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X6 source.t0 plus.t1 drain_left.t4 a_n1220_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X7 source.t11 plus.t2 drain_left.t3 a_n1220_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X8 drain_right.t2 minus.t3 source.t10 a_n1220_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X9 drain_left.t2 plus.t3 source.t4 a_n1220_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X10 a_n1220_n5888# a_n1220_n5888# a_n1220_n5888# a_n1220_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X11 source.t5 minus.t4 drain_right.t1 a_n1220_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X12 source.t9 minus.t5 drain_right.t0 a_n1220_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=4.125 ps=25.33 w=25 l=0.3
X13 a_n1220_n5888# a_n1220_n5888# a_n1220_n5888# a_n1220_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=0 ps=0 w=25 l=0.3
X14 drain_left.t1 plus.t4 source.t1 a_n1220_n5888# sky130_fd_pr__nfet_01v8 ad=4.125 pd=25.33 as=9.75 ps=50.78 w=25 l=0.3
X15 drain_left.t0 plus.t5 source.t2 a_n1220_n5888# sky130_fd_pr__nfet_01v8 ad=9.75 pd=50.78 as=4.125 ps=25.33 w=25 l=0.3
R0 minus.n2 minus.t0 2168.27
R1 minus.n0 minus.t3 2168.27
R2 minus.n6 minus.t1 2168.27
R3 minus.n4 minus.t2 2168.27
R4 minus.n1 minus.t5 2112.77
R5 minus.n5 minus.t4 2112.77
R6 minus.n3 minus.n0 161.489
R7 minus.n7 minus.n4 161.489
R8 minus.n3 minus.n2 161.3
R9 minus.n7 minus.n6 161.3
R10 minus.n8 minus.n3 43.6236
R11 minus.n2 minus.n1 36.5157
R12 minus.n1 minus.n0 36.5157
R13 minus.n5 minus.n4 36.5157
R14 minus.n6 minus.n5 36.5157
R15 minus.n8 minus.n7 6.5327
R16 minus minus.n8 0.188
R17 source.n562 source.n428 289.615
R18 source.n420 source.n286 289.615
R19 source.n134 source.n0 289.615
R20 source.n276 source.n142 289.615
R21 source.n472 source.n471 185
R22 source.n477 source.n476 185
R23 source.n479 source.n478 185
R24 source.n468 source.n467 185
R25 source.n485 source.n484 185
R26 source.n487 source.n486 185
R27 source.n464 source.n463 185
R28 source.n494 source.n493 185
R29 source.n495 source.n462 185
R30 source.n497 source.n496 185
R31 source.n460 source.n459 185
R32 source.n503 source.n502 185
R33 source.n505 source.n504 185
R34 source.n456 source.n455 185
R35 source.n511 source.n510 185
R36 source.n513 source.n512 185
R37 source.n452 source.n451 185
R38 source.n519 source.n518 185
R39 source.n521 source.n520 185
R40 source.n448 source.n447 185
R41 source.n527 source.n526 185
R42 source.n529 source.n528 185
R43 source.n444 source.n443 185
R44 source.n535 source.n534 185
R45 source.n538 source.n537 185
R46 source.n536 source.n440 185
R47 source.n543 source.n439 185
R48 source.n545 source.n544 185
R49 source.n547 source.n546 185
R50 source.n436 source.n435 185
R51 source.n553 source.n552 185
R52 source.n555 source.n554 185
R53 source.n432 source.n431 185
R54 source.n561 source.n560 185
R55 source.n563 source.n562 185
R56 source.n330 source.n329 185
R57 source.n335 source.n334 185
R58 source.n337 source.n336 185
R59 source.n326 source.n325 185
R60 source.n343 source.n342 185
R61 source.n345 source.n344 185
R62 source.n322 source.n321 185
R63 source.n352 source.n351 185
R64 source.n353 source.n320 185
R65 source.n355 source.n354 185
R66 source.n318 source.n317 185
R67 source.n361 source.n360 185
R68 source.n363 source.n362 185
R69 source.n314 source.n313 185
R70 source.n369 source.n368 185
R71 source.n371 source.n370 185
R72 source.n310 source.n309 185
R73 source.n377 source.n376 185
R74 source.n379 source.n378 185
R75 source.n306 source.n305 185
R76 source.n385 source.n384 185
R77 source.n387 source.n386 185
R78 source.n302 source.n301 185
R79 source.n393 source.n392 185
R80 source.n396 source.n395 185
R81 source.n394 source.n298 185
R82 source.n401 source.n297 185
R83 source.n403 source.n402 185
R84 source.n405 source.n404 185
R85 source.n294 source.n293 185
R86 source.n411 source.n410 185
R87 source.n413 source.n412 185
R88 source.n290 source.n289 185
R89 source.n419 source.n418 185
R90 source.n421 source.n420 185
R91 source.n135 source.n134 185
R92 source.n133 source.n132 185
R93 source.n4 source.n3 185
R94 source.n127 source.n126 185
R95 source.n125 source.n124 185
R96 source.n8 source.n7 185
R97 source.n119 source.n118 185
R98 source.n117 source.n116 185
R99 source.n115 source.n11 185
R100 source.n15 source.n12 185
R101 source.n110 source.n109 185
R102 source.n108 source.n107 185
R103 source.n17 source.n16 185
R104 source.n102 source.n101 185
R105 source.n100 source.n99 185
R106 source.n21 source.n20 185
R107 source.n94 source.n93 185
R108 source.n92 source.n91 185
R109 source.n25 source.n24 185
R110 source.n86 source.n85 185
R111 source.n84 source.n83 185
R112 source.n29 source.n28 185
R113 source.n78 source.n77 185
R114 source.n76 source.n75 185
R115 source.n33 source.n32 185
R116 source.n70 source.n69 185
R117 source.n68 source.n35 185
R118 source.n67 source.n66 185
R119 source.n38 source.n36 185
R120 source.n61 source.n60 185
R121 source.n59 source.n58 185
R122 source.n42 source.n41 185
R123 source.n53 source.n52 185
R124 source.n51 source.n50 185
R125 source.n46 source.n45 185
R126 source.n277 source.n276 185
R127 source.n275 source.n274 185
R128 source.n146 source.n145 185
R129 source.n269 source.n268 185
R130 source.n267 source.n266 185
R131 source.n150 source.n149 185
R132 source.n261 source.n260 185
R133 source.n259 source.n258 185
R134 source.n257 source.n153 185
R135 source.n157 source.n154 185
R136 source.n252 source.n251 185
R137 source.n250 source.n249 185
R138 source.n159 source.n158 185
R139 source.n244 source.n243 185
R140 source.n242 source.n241 185
R141 source.n163 source.n162 185
R142 source.n236 source.n235 185
R143 source.n234 source.n233 185
R144 source.n167 source.n166 185
R145 source.n228 source.n227 185
R146 source.n226 source.n225 185
R147 source.n171 source.n170 185
R148 source.n220 source.n219 185
R149 source.n218 source.n217 185
R150 source.n175 source.n174 185
R151 source.n212 source.n211 185
R152 source.n210 source.n177 185
R153 source.n209 source.n208 185
R154 source.n180 source.n178 185
R155 source.n203 source.n202 185
R156 source.n201 source.n200 185
R157 source.n184 source.n183 185
R158 source.n195 source.n194 185
R159 source.n193 source.n192 185
R160 source.n188 source.n187 185
R161 source.n473 source.t7 149.524
R162 source.n331 source.t1 149.524
R163 source.n47 source.t4 149.524
R164 source.n189 source.t10 149.524
R165 source.n477 source.n471 104.615
R166 source.n478 source.n477 104.615
R167 source.n478 source.n467 104.615
R168 source.n485 source.n467 104.615
R169 source.n486 source.n485 104.615
R170 source.n486 source.n463 104.615
R171 source.n494 source.n463 104.615
R172 source.n495 source.n494 104.615
R173 source.n496 source.n495 104.615
R174 source.n496 source.n459 104.615
R175 source.n503 source.n459 104.615
R176 source.n504 source.n503 104.615
R177 source.n504 source.n455 104.615
R178 source.n511 source.n455 104.615
R179 source.n512 source.n511 104.615
R180 source.n512 source.n451 104.615
R181 source.n519 source.n451 104.615
R182 source.n520 source.n519 104.615
R183 source.n520 source.n447 104.615
R184 source.n527 source.n447 104.615
R185 source.n528 source.n527 104.615
R186 source.n528 source.n443 104.615
R187 source.n535 source.n443 104.615
R188 source.n537 source.n535 104.615
R189 source.n537 source.n536 104.615
R190 source.n536 source.n439 104.615
R191 source.n545 source.n439 104.615
R192 source.n546 source.n545 104.615
R193 source.n546 source.n435 104.615
R194 source.n553 source.n435 104.615
R195 source.n554 source.n553 104.615
R196 source.n554 source.n431 104.615
R197 source.n561 source.n431 104.615
R198 source.n562 source.n561 104.615
R199 source.n335 source.n329 104.615
R200 source.n336 source.n335 104.615
R201 source.n336 source.n325 104.615
R202 source.n343 source.n325 104.615
R203 source.n344 source.n343 104.615
R204 source.n344 source.n321 104.615
R205 source.n352 source.n321 104.615
R206 source.n353 source.n352 104.615
R207 source.n354 source.n353 104.615
R208 source.n354 source.n317 104.615
R209 source.n361 source.n317 104.615
R210 source.n362 source.n361 104.615
R211 source.n362 source.n313 104.615
R212 source.n369 source.n313 104.615
R213 source.n370 source.n369 104.615
R214 source.n370 source.n309 104.615
R215 source.n377 source.n309 104.615
R216 source.n378 source.n377 104.615
R217 source.n378 source.n305 104.615
R218 source.n385 source.n305 104.615
R219 source.n386 source.n385 104.615
R220 source.n386 source.n301 104.615
R221 source.n393 source.n301 104.615
R222 source.n395 source.n393 104.615
R223 source.n395 source.n394 104.615
R224 source.n394 source.n297 104.615
R225 source.n403 source.n297 104.615
R226 source.n404 source.n403 104.615
R227 source.n404 source.n293 104.615
R228 source.n411 source.n293 104.615
R229 source.n412 source.n411 104.615
R230 source.n412 source.n289 104.615
R231 source.n419 source.n289 104.615
R232 source.n420 source.n419 104.615
R233 source.n134 source.n133 104.615
R234 source.n133 source.n3 104.615
R235 source.n126 source.n3 104.615
R236 source.n126 source.n125 104.615
R237 source.n125 source.n7 104.615
R238 source.n118 source.n7 104.615
R239 source.n118 source.n117 104.615
R240 source.n117 source.n11 104.615
R241 source.n15 source.n11 104.615
R242 source.n109 source.n15 104.615
R243 source.n109 source.n108 104.615
R244 source.n108 source.n16 104.615
R245 source.n101 source.n16 104.615
R246 source.n101 source.n100 104.615
R247 source.n100 source.n20 104.615
R248 source.n93 source.n20 104.615
R249 source.n93 source.n92 104.615
R250 source.n92 source.n24 104.615
R251 source.n85 source.n24 104.615
R252 source.n85 source.n84 104.615
R253 source.n84 source.n28 104.615
R254 source.n77 source.n28 104.615
R255 source.n77 source.n76 104.615
R256 source.n76 source.n32 104.615
R257 source.n69 source.n32 104.615
R258 source.n69 source.n68 104.615
R259 source.n68 source.n67 104.615
R260 source.n67 source.n36 104.615
R261 source.n60 source.n36 104.615
R262 source.n60 source.n59 104.615
R263 source.n59 source.n41 104.615
R264 source.n52 source.n41 104.615
R265 source.n52 source.n51 104.615
R266 source.n51 source.n45 104.615
R267 source.n276 source.n275 104.615
R268 source.n275 source.n145 104.615
R269 source.n268 source.n145 104.615
R270 source.n268 source.n267 104.615
R271 source.n267 source.n149 104.615
R272 source.n260 source.n149 104.615
R273 source.n260 source.n259 104.615
R274 source.n259 source.n153 104.615
R275 source.n157 source.n153 104.615
R276 source.n251 source.n157 104.615
R277 source.n251 source.n250 104.615
R278 source.n250 source.n158 104.615
R279 source.n243 source.n158 104.615
R280 source.n243 source.n242 104.615
R281 source.n242 source.n162 104.615
R282 source.n235 source.n162 104.615
R283 source.n235 source.n234 104.615
R284 source.n234 source.n166 104.615
R285 source.n227 source.n166 104.615
R286 source.n227 source.n226 104.615
R287 source.n226 source.n170 104.615
R288 source.n219 source.n170 104.615
R289 source.n219 source.n218 104.615
R290 source.n218 source.n174 104.615
R291 source.n211 source.n174 104.615
R292 source.n211 source.n210 104.615
R293 source.n210 source.n209 104.615
R294 source.n209 source.n178 104.615
R295 source.n202 source.n178 104.615
R296 source.n202 source.n201 104.615
R297 source.n201 source.n183 104.615
R298 source.n194 source.n183 104.615
R299 source.n194 source.n193 104.615
R300 source.n193 source.n187 104.615
R301 source.t7 source.n471 52.3082
R302 source.t1 source.n329 52.3082
R303 source.t4 source.n45 52.3082
R304 source.t10 source.n187 52.3082
R305 source.n427 source.n426 42.0366
R306 source.n285 source.n284 42.0366
R307 source.n141 source.n140 42.0366
R308 source.n283 source.n282 42.0366
R309 source.n285 source.n283 32.2224
R310 source.n567 source.n566 30.6338
R311 source.n425 source.n424 30.6338
R312 source.n139 source.n138 30.6338
R313 source.n281 source.n280 30.6338
R314 source.n568 source.n139 26.1448
R315 source.n497 source.n462 13.1884
R316 source.n544 source.n543 13.1884
R317 source.n355 source.n320 13.1884
R318 source.n402 source.n401 13.1884
R319 source.n116 source.n115 13.1884
R320 source.n70 source.n35 13.1884
R321 source.n258 source.n257 13.1884
R322 source.n212 source.n177 13.1884
R323 source.n493 source.n492 12.8005
R324 source.n498 source.n460 12.8005
R325 source.n542 source.n440 12.8005
R326 source.n547 source.n438 12.8005
R327 source.n351 source.n350 12.8005
R328 source.n356 source.n318 12.8005
R329 source.n400 source.n298 12.8005
R330 source.n405 source.n296 12.8005
R331 source.n119 source.n10 12.8005
R332 source.n114 source.n12 12.8005
R333 source.n71 source.n33 12.8005
R334 source.n66 source.n37 12.8005
R335 source.n261 source.n152 12.8005
R336 source.n256 source.n154 12.8005
R337 source.n213 source.n175 12.8005
R338 source.n208 source.n179 12.8005
R339 source.n491 source.n464 12.0247
R340 source.n502 source.n501 12.0247
R341 source.n539 source.n538 12.0247
R342 source.n548 source.n436 12.0247
R343 source.n349 source.n322 12.0247
R344 source.n360 source.n359 12.0247
R345 source.n397 source.n396 12.0247
R346 source.n406 source.n294 12.0247
R347 source.n120 source.n8 12.0247
R348 source.n111 source.n110 12.0247
R349 source.n75 source.n74 12.0247
R350 source.n65 source.n38 12.0247
R351 source.n262 source.n150 12.0247
R352 source.n253 source.n252 12.0247
R353 source.n217 source.n216 12.0247
R354 source.n207 source.n180 12.0247
R355 source.n488 source.n487 11.249
R356 source.n505 source.n458 11.249
R357 source.n534 source.n442 11.249
R358 source.n552 source.n551 11.249
R359 source.n346 source.n345 11.249
R360 source.n363 source.n316 11.249
R361 source.n392 source.n300 11.249
R362 source.n410 source.n409 11.249
R363 source.n124 source.n123 11.249
R364 source.n107 source.n14 11.249
R365 source.n78 source.n31 11.249
R366 source.n62 source.n61 11.249
R367 source.n266 source.n265 11.249
R368 source.n249 source.n156 11.249
R369 source.n220 source.n173 11.249
R370 source.n204 source.n203 11.249
R371 source.n484 source.n466 10.4732
R372 source.n506 source.n456 10.4732
R373 source.n533 source.n444 10.4732
R374 source.n555 source.n434 10.4732
R375 source.n342 source.n324 10.4732
R376 source.n364 source.n314 10.4732
R377 source.n391 source.n302 10.4732
R378 source.n413 source.n292 10.4732
R379 source.n127 source.n6 10.4732
R380 source.n106 source.n17 10.4732
R381 source.n79 source.n29 10.4732
R382 source.n58 source.n40 10.4732
R383 source.n269 source.n148 10.4732
R384 source.n248 source.n159 10.4732
R385 source.n221 source.n171 10.4732
R386 source.n200 source.n182 10.4732
R387 source.n473 source.n472 10.2747
R388 source.n331 source.n330 10.2747
R389 source.n47 source.n46 10.2747
R390 source.n189 source.n188 10.2747
R391 source.n483 source.n468 9.69747
R392 source.n510 source.n509 9.69747
R393 source.n530 source.n529 9.69747
R394 source.n556 source.n432 9.69747
R395 source.n341 source.n326 9.69747
R396 source.n368 source.n367 9.69747
R397 source.n388 source.n387 9.69747
R398 source.n414 source.n290 9.69747
R399 source.n128 source.n4 9.69747
R400 source.n103 source.n102 9.69747
R401 source.n83 source.n82 9.69747
R402 source.n57 source.n42 9.69747
R403 source.n270 source.n146 9.69747
R404 source.n245 source.n244 9.69747
R405 source.n225 source.n224 9.69747
R406 source.n199 source.n184 9.69747
R407 source.n566 source.n565 9.45567
R408 source.n424 source.n423 9.45567
R409 source.n138 source.n137 9.45567
R410 source.n280 source.n279 9.45567
R411 source.n430 source.n429 9.3005
R412 source.n559 source.n558 9.3005
R413 source.n557 source.n556 9.3005
R414 source.n434 source.n433 9.3005
R415 source.n551 source.n550 9.3005
R416 source.n549 source.n548 9.3005
R417 source.n438 source.n437 9.3005
R418 source.n517 source.n516 9.3005
R419 source.n515 source.n514 9.3005
R420 source.n454 source.n453 9.3005
R421 source.n509 source.n508 9.3005
R422 source.n507 source.n506 9.3005
R423 source.n458 source.n457 9.3005
R424 source.n501 source.n500 9.3005
R425 source.n499 source.n498 9.3005
R426 source.n475 source.n474 9.3005
R427 source.n470 source.n469 9.3005
R428 source.n481 source.n480 9.3005
R429 source.n483 source.n482 9.3005
R430 source.n466 source.n465 9.3005
R431 source.n489 source.n488 9.3005
R432 source.n491 source.n490 9.3005
R433 source.n492 source.n461 9.3005
R434 source.n450 source.n449 9.3005
R435 source.n523 source.n522 9.3005
R436 source.n525 source.n524 9.3005
R437 source.n446 source.n445 9.3005
R438 source.n531 source.n530 9.3005
R439 source.n533 source.n532 9.3005
R440 source.n442 source.n441 9.3005
R441 source.n540 source.n539 9.3005
R442 source.n542 source.n541 9.3005
R443 source.n565 source.n564 9.3005
R444 source.n288 source.n287 9.3005
R445 source.n417 source.n416 9.3005
R446 source.n415 source.n414 9.3005
R447 source.n292 source.n291 9.3005
R448 source.n409 source.n408 9.3005
R449 source.n407 source.n406 9.3005
R450 source.n296 source.n295 9.3005
R451 source.n375 source.n374 9.3005
R452 source.n373 source.n372 9.3005
R453 source.n312 source.n311 9.3005
R454 source.n367 source.n366 9.3005
R455 source.n365 source.n364 9.3005
R456 source.n316 source.n315 9.3005
R457 source.n359 source.n358 9.3005
R458 source.n357 source.n356 9.3005
R459 source.n333 source.n332 9.3005
R460 source.n328 source.n327 9.3005
R461 source.n339 source.n338 9.3005
R462 source.n341 source.n340 9.3005
R463 source.n324 source.n323 9.3005
R464 source.n347 source.n346 9.3005
R465 source.n349 source.n348 9.3005
R466 source.n350 source.n319 9.3005
R467 source.n308 source.n307 9.3005
R468 source.n381 source.n380 9.3005
R469 source.n383 source.n382 9.3005
R470 source.n304 source.n303 9.3005
R471 source.n389 source.n388 9.3005
R472 source.n391 source.n390 9.3005
R473 source.n300 source.n299 9.3005
R474 source.n398 source.n397 9.3005
R475 source.n400 source.n399 9.3005
R476 source.n423 source.n422 9.3005
R477 source.n49 source.n48 9.3005
R478 source.n44 source.n43 9.3005
R479 source.n55 source.n54 9.3005
R480 source.n57 source.n56 9.3005
R481 source.n40 source.n39 9.3005
R482 source.n63 source.n62 9.3005
R483 source.n65 source.n64 9.3005
R484 source.n37 source.n34 9.3005
R485 source.n96 source.n95 9.3005
R486 source.n98 source.n97 9.3005
R487 source.n19 source.n18 9.3005
R488 source.n104 source.n103 9.3005
R489 source.n106 source.n105 9.3005
R490 source.n14 source.n13 9.3005
R491 source.n112 source.n111 9.3005
R492 source.n114 source.n113 9.3005
R493 source.n137 source.n136 9.3005
R494 source.n2 source.n1 9.3005
R495 source.n131 source.n130 9.3005
R496 source.n129 source.n128 9.3005
R497 source.n6 source.n5 9.3005
R498 source.n123 source.n122 9.3005
R499 source.n121 source.n120 9.3005
R500 source.n10 source.n9 9.3005
R501 source.n23 source.n22 9.3005
R502 source.n90 source.n89 9.3005
R503 source.n88 source.n87 9.3005
R504 source.n27 source.n26 9.3005
R505 source.n82 source.n81 9.3005
R506 source.n80 source.n79 9.3005
R507 source.n31 source.n30 9.3005
R508 source.n74 source.n73 9.3005
R509 source.n72 source.n71 9.3005
R510 source.n191 source.n190 9.3005
R511 source.n186 source.n185 9.3005
R512 source.n197 source.n196 9.3005
R513 source.n199 source.n198 9.3005
R514 source.n182 source.n181 9.3005
R515 source.n205 source.n204 9.3005
R516 source.n207 source.n206 9.3005
R517 source.n179 source.n176 9.3005
R518 source.n238 source.n237 9.3005
R519 source.n240 source.n239 9.3005
R520 source.n161 source.n160 9.3005
R521 source.n246 source.n245 9.3005
R522 source.n248 source.n247 9.3005
R523 source.n156 source.n155 9.3005
R524 source.n254 source.n253 9.3005
R525 source.n256 source.n255 9.3005
R526 source.n279 source.n278 9.3005
R527 source.n144 source.n143 9.3005
R528 source.n273 source.n272 9.3005
R529 source.n271 source.n270 9.3005
R530 source.n148 source.n147 9.3005
R531 source.n265 source.n264 9.3005
R532 source.n263 source.n262 9.3005
R533 source.n152 source.n151 9.3005
R534 source.n165 source.n164 9.3005
R535 source.n232 source.n231 9.3005
R536 source.n230 source.n229 9.3005
R537 source.n169 source.n168 9.3005
R538 source.n224 source.n223 9.3005
R539 source.n222 source.n221 9.3005
R540 source.n173 source.n172 9.3005
R541 source.n216 source.n215 9.3005
R542 source.n214 source.n213 9.3005
R543 source.n480 source.n479 8.92171
R544 source.n513 source.n454 8.92171
R545 source.n526 source.n446 8.92171
R546 source.n560 source.n559 8.92171
R547 source.n338 source.n337 8.92171
R548 source.n371 source.n312 8.92171
R549 source.n384 source.n304 8.92171
R550 source.n418 source.n417 8.92171
R551 source.n132 source.n131 8.92171
R552 source.n99 source.n19 8.92171
R553 source.n86 source.n27 8.92171
R554 source.n54 source.n53 8.92171
R555 source.n274 source.n273 8.92171
R556 source.n241 source.n161 8.92171
R557 source.n228 source.n169 8.92171
R558 source.n196 source.n195 8.92171
R559 source.n476 source.n470 8.14595
R560 source.n514 source.n452 8.14595
R561 source.n525 source.n448 8.14595
R562 source.n563 source.n430 8.14595
R563 source.n334 source.n328 8.14595
R564 source.n372 source.n310 8.14595
R565 source.n383 source.n306 8.14595
R566 source.n421 source.n288 8.14595
R567 source.n135 source.n2 8.14595
R568 source.n98 source.n21 8.14595
R569 source.n87 source.n25 8.14595
R570 source.n50 source.n44 8.14595
R571 source.n277 source.n144 8.14595
R572 source.n240 source.n163 8.14595
R573 source.n229 source.n167 8.14595
R574 source.n192 source.n186 8.14595
R575 source.n475 source.n472 7.3702
R576 source.n518 source.n517 7.3702
R577 source.n522 source.n521 7.3702
R578 source.n564 source.n428 7.3702
R579 source.n333 source.n330 7.3702
R580 source.n376 source.n375 7.3702
R581 source.n380 source.n379 7.3702
R582 source.n422 source.n286 7.3702
R583 source.n136 source.n0 7.3702
R584 source.n95 source.n94 7.3702
R585 source.n91 source.n90 7.3702
R586 source.n49 source.n46 7.3702
R587 source.n278 source.n142 7.3702
R588 source.n237 source.n236 7.3702
R589 source.n233 source.n232 7.3702
R590 source.n191 source.n188 7.3702
R591 source.n518 source.n450 6.59444
R592 source.n521 source.n450 6.59444
R593 source.n566 source.n428 6.59444
R594 source.n376 source.n308 6.59444
R595 source.n379 source.n308 6.59444
R596 source.n424 source.n286 6.59444
R597 source.n138 source.n0 6.59444
R598 source.n94 source.n23 6.59444
R599 source.n91 source.n23 6.59444
R600 source.n280 source.n142 6.59444
R601 source.n236 source.n165 6.59444
R602 source.n233 source.n165 6.59444
R603 source.n476 source.n475 5.81868
R604 source.n517 source.n452 5.81868
R605 source.n522 source.n448 5.81868
R606 source.n564 source.n563 5.81868
R607 source.n334 source.n333 5.81868
R608 source.n375 source.n310 5.81868
R609 source.n380 source.n306 5.81868
R610 source.n422 source.n421 5.81868
R611 source.n136 source.n135 5.81868
R612 source.n95 source.n21 5.81868
R613 source.n90 source.n25 5.81868
R614 source.n50 source.n49 5.81868
R615 source.n278 source.n277 5.81868
R616 source.n237 source.n163 5.81868
R617 source.n232 source.n167 5.81868
R618 source.n192 source.n191 5.81868
R619 source.n568 source.n567 5.53498
R620 source.n479 source.n470 5.04292
R621 source.n514 source.n513 5.04292
R622 source.n526 source.n525 5.04292
R623 source.n560 source.n430 5.04292
R624 source.n337 source.n328 5.04292
R625 source.n372 source.n371 5.04292
R626 source.n384 source.n383 5.04292
R627 source.n418 source.n288 5.04292
R628 source.n132 source.n2 5.04292
R629 source.n99 source.n98 5.04292
R630 source.n87 source.n86 5.04292
R631 source.n53 source.n44 5.04292
R632 source.n274 source.n144 5.04292
R633 source.n241 source.n240 5.04292
R634 source.n229 source.n228 5.04292
R635 source.n195 source.n186 5.04292
R636 source.n480 source.n468 4.26717
R637 source.n510 source.n454 4.26717
R638 source.n529 source.n446 4.26717
R639 source.n559 source.n432 4.26717
R640 source.n338 source.n326 4.26717
R641 source.n368 source.n312 4.26717
R642 source.n387 source.n304 4.26717
R643 source.n417 source.n290 4.26717
R644 source.n131 source.n4 4.26717
R645 source.n102 source.n19 4.26717
R646 source.n83 source.n27 4.26717
R647 source.n54 source.n42 4.26717
R648 source.n273 source.n146 4.26717
R649 source.n244 source.n161 4.26717
R650 source.n225 source.n169 4.26717
R651 source.n196 source.n184 4.26717
R652 source.n484 source.n483 3.49141
R653 source.n509 source.n456 3.49141
R654 source.n530 source.n444 3.49141
R655 source.n556 source.n555 3.49141
R656 source.n342 source.n341 3.49141
R657 source.n367 source.n314 3.49141
R658 source.n388 source.n302 3.49141
R659 source.n414 source.n413 3.49141
R660 source.n128 source.n127 3.49141
R661 source.n103 source.n17 3.49141
R662 source.n82 source.n29 3.49141
R663 source.n58 source.n57 3.49141
R664 source.n270 source.n269 3.49141
R665 source.n245 source.n159 3.49141
R666 source.n224 source.n171 3.49141
R667 source.n200 source.n199 3.49141
R668 source.n48 source.n47 2.84303
R669 source.n190 source.n189 2.84303
R670 source.n474 source.n473 2.84303
R671 source.n332 source.n331 2.84303
R672 source.n487 source.n466 2.71565
R673 source.n506 source.n505 2.71565
R674 source.n534 source.n533 2.71565
R675 source.n552 source.n434 2.71565
R676 source.n345 source.n324 2.71565
R677 source.n364 source.n363 2.71565
R678 source.n392 source.n391 2.71565
R679 source.n410 source.n292 2.71565
R680 source.n124 source.n6 2.71565
R681 source.n107 source.n106 2.71565
R682 source.n79 source.n78 2.71565
R683 source.n61 source.n40 2.71565
R684 source.n266 source.n148 2.71565
R685 source.n249 source.n248 2.71565
R686 source.n221 source.n220 2.71565
R687 source.n203 source.n182 2.71565
R688 source.n488 source.n464 1.93989
R689 source.n502 source.n458 1.93989
R690 source.n538 source.n442 1.93989
R691 source.n551 source.n436 1.93989
R692 source.n346 source.n322 1.93989
R693 source.n360 source.n316 1.93989
R694 source.n396 source.n300 1.93989
R695 source.n409 source.n294 1.93989
R696 source.n123 source.n8 1.93989
R697 source.n110 source.n14 1.93989
R698 source.n75 source.n31 1.93989
R699 source.n62 source.n38 1.93989
R700 source.n265 source.n150 1.93989
R701 source.n252 source.n156 1.93989
R702 source.n217 source.n173 1.93989
R703 source.n204 source.n180 1.93989
R704 source.n493 source.n491 1.16414
R705 source.n501 source.n460 1.16414
R706 source.n539 source.n440 1.16414
R707 source.n548 source.n547 1.16414
R708 source.n351 source.n349 1.16414
R709 source.n359 source.n318 1.16414
R710 source.n397 source.n298 1.16414
R711 source.n406 source.n405 1.16414
R712 source.n120 source.n119 1.16414
R713 source.n111 source.n12 1.16414
R714 source.n74 source.n33 1.16414
R715 source.n66 source.n65 1.16414
R716 source.n262 source.n261 1.16414
R717 source.n253 source.n154 1.16414
R718 source.n216 source.n175 1.16414
R719 source.n208 source.n207 1.16414
R720 source.n426 source.t6 0.7925
R721 source.n426 source.t5 0.7925
R722 source.n284 source.t2 0.7925
R723 source.n284 source.t11 0.7925
R724 source.n140 source.t3 0.7925
R725 source.n140 source.t0 0.7925
R726 source.n282 source.t8 0.7925
R727 source.n282 source.t9 0.7925
R728 source.n281 source.n141 0.741879
R729 source.n427 source.n425 0.741879
R730 source.n283 source.n281 0.543603
R731 source.n141 source.n139 0.543603
R732 source.n425 source.n285 0.543603
R733 source.n567 source.n427 0.543603
R734 source.n492 source.n462 0.388379
R735 source.n498 source.n497 0.388379
R736 source.n543 source.n542 0.388379
R737 source.n544 source.n438 0.388379
R738 source.n350 source.n320 0.388379
R739 source.n356 source.n355 0.388379
R740 source.n401 source.n400 0.388379
R741 source.n402 source.n296 0.388379
R742 source.n116 source.n10 0.388379
R743 source.n115 source.n114 0.388379
R744 source.n71 source.n70 0.388379
R745 source.n37 source.n35 0.388379
R746 source.n258 source.n152 0.388379
R747 source.n257 source.n256 0.388379
R748 source.n213 source.n212 0.388379
R749 source.n179 source.n177 0.388379
R750 source source.n568 0.188
R751 source.n474 source.n469 0.155672
R752 source.n481 source.n469 0.155672
R753 source.n482 source.n481 0.155672
R754 source.n482 source.n465 0.155672
R755 source.n489 source.n465 0.155672
R756 source.n490 source.n489 0.155672
R757 source.n490 source.n461 0.155672
R758 source.n499 source.n461 0.155672
R759 source.n500 source.n499 0.155672
R760 source.n500 source.n457 0.155672
R761 source.n507 source.n457 0.155672
R762 source.n508 source.n507 0.155672
R763 source.n508 source.n453 0.155672
R764 source.n515 source.n453 0.155672
R765 source.n516 source.n515 0.155672
R766 source.n516 source.n449 0.155672
R767 source.n523 source.n449 0.155672
R768 source.n524 source.n523 0.155672
R769 source.n524 source.n445 0.155672
R770 source.n531 source.n445 0.155672
R771 source.n532 source.n531 0.155672
R772 source.n532 source.n441 0.155672
R773 source.n540 source.n441 0.155672
R774 source.n541 source.n540 0.155672
R775 source.n541 source.n437 0.155672
R776 source.n549 source.n437 0.155672
R777 source.n550 source.n549 0.155672
R778 source.n550 source.n433 0.155672
R779 source.n557 source.n433 0.155672
R780 source.n558 source.n557 0.155672
R781 source.n558 source.n429 0.155672
R782 source.n565 source.n429 0.155672
R783 source.n332 source.n327 0.155672
R784 source.n339 source.n327 0.155672
R785 source.n340 source.n339 0.155672
R786 source.n340 source.n323 0.155672
R787 source.n347 source.n323 0.155672
R788 source.n348 source.n347 0.155672
R789 source.n348 source.n319 0.155672
R790 source.n357 source.n319 0.155672
R791 source.n358 source.n357 0.155672
R792 source.n358 source.n315 0.155672
R793 source.n365 source.n315 0.155672
R794 source.n366 source.n365 0.155672
R795 source.n366 source.n311 0.155672
R796 source.n373 source.n311 0.155672
R797 source.n374 source.n373 0.155672
R798 source.n374 source.n307 0.155672
R799 source.n381 source.n307 0.155672
R800 source.n382 source.n381 0.155672
R801 source.n382 source.n303 0.155672
R802 source.n389 source.n303 0.155672
R803 source.n390 source.n389 0.155672
R804 source.n390 source.n299 0.155672
R805 source.n398 source.n299 0.155672
R806 source.n399 source.n398 0.155672
R807 source.n399 source.n295 0.155672
R808 source.n407 source.n295 0.155672
R809 source.n408 source.n407 0.155672
R810 source.n408 source.n291 0.155672
R811 source.n415 source.n291 0.155672
R812 source.n416 source.n415 0.155672
R813 source.n416 source.n287 0.155672
R814 source.n423 source.n287 0.155672
R815 source.n137 source.n1 0.155672
R816 source.n130 source.n1 0.155672
R817 source.n130 source.n129 0.155672
R818 source.n129 source.n5 0.155672
R819 source.n122 source.n5 0.155672
R820 source.n122 source.n121 0.155672
R821 source.n121 source.n9 0.155672
R822 source.n113 source.n9 0.155672
R823 source.n113 source.n112 0.155672
R824 source.n112 source.n13 0.155672
R825 source.n105 source.n13 0.155672
R826 source.n105 source.n104 0.155672
R827 source.n104 source.n18 0.155672
R828 source.n97 source.n18 0.155672
R829 source.n97 source.n96 0.155672
R830 source.n96 source.n22 0.155672
R831 source.n89 source.n22 0.155672
R832 source.n89 source.n88 0.155672
R833 source.n88 source.n26 0.155672
R834 source.n81 source.n26 0.155672
R835 source.n81 source.n80 0.155672
R836 source.n80 source.n30 0.155672
R837 source.n73 source.n30 0.155672
R838 source.n73 source.n72 0.155672
R839 source.n72 source.n34 0.155672
R840 source.n64 source.n34 0.155672
R841 source.n64 source.n63 0.155672
R842 source.n63 source.n39 0.155672
R843 source.n56 source.n39 0.155672
R844 source.n56 source.n55 0.155672
R845 source.n55 source.n43 0.155672
R846 source.n48 source.n43 0.155672
R847 source.n279 source.n143 0.155672
R848 source.n272 source.n143 0.155672
R849 source.n272 source.n271 0.155672
R850 source.n271 source.n147 0.155672
R851 source.n264 source.n147 0.155672
R852 source.n264 source.n263 0.155672
R853 source.n263 source.n151 0.155672
R854 source.n255 source.n151 0.155672
R855 source.n255 source.n254 0.155672
R856 source.n254 source.n155 0.155672
R857 source.n247 source.n155 0.155672
R858 source.n247 source.n246 0.155672
R859 source.n246 source.n160 0.155672
R860 source.n239 source.n160 0.155672
R861 source.n239 source.n238 0.155672
R862 source.n238 source.n164 0.155672
R863 source.n231 source.n164 0.155672
R864 source.n231 source.n230 0.155672
R865 source.n230 source.n168 0.155672
R866 source.n223 source.n168 0.155672
R867 source.n223 source.n222 0.155672
R868 source.n222 source.n172 0.155672
R869 source.n215 source.n172 0.155672
R870 source.n215 source.n214 0.155672
R871 source.n214 source.n176 0.155672
R872 source.n206 source.n176 0.155672
R873 source.n206 source.n205 0.155672
R874 source.n205 source.n181 0.155672
R875 source.n198 source.n181 0.155672
R876 source.n198 source.n197 0.155672
R877 source.n197 source.n185 0.155672
R878 source.n190 source.n185 0.155672
R879 drain_right.n134 drain_right.n0 289.615
R880 drain_right.n276 drain_right.n142 289.615
R881 drain_right.n44 drain_right.n43 185
R882 drain_right.n49 drain_right.n48 185
R883 drain_right.n51 drain_right.n50 185
R884 drain_right.n40 drain_right.n39 185
R885 drain_right.n57 drain_right.n56 185
R886 drain_right.n59 drain_right.n58 185
R887 drain_right.n36 drain_right.n35 185
R888 drain_right.n66 drain_right.n65 185
R889 drain_right.n67 drain_right.n34 185
R890 drain_right.n69 drain_right.n68 185
R891 drain_right.n32 drain_right.n31 185
R892 drain_right.n75 drain_right.n74 185
R893 drain_right.n77 drain_right.n76 185
R894 drain_right.n28 drain_right.n27 185
R895 drain_right.n83 drain_right.n82 185
R896 drain_right.n85 drain_right.n84 185
R897 drain_right.n24 drain_right.n23 185
R898 drain_right.n91 drain_right.n90 185
R899 drain_right.n93 drain_right.n92 185
R900 drain_right.n20 drain_right.n19 185
R901 drain_right.n99 drain_right.n98 185
R902 drain_right.n101 drain_right.n100 185
R903 drain_right.n16 drain_right.n15 185
R904 drain_right.n107 drain_right.n106 185
R905 drain_right.n110 drain_right.n109 185
R906 drain_right.n108 drain_right.n12 185
R907 drain_right.n115 drain_right.n11 185
R908 drain_right.n117 drain_right.n116 185
R909 drain_right.n119 drain_right.n118 185
R910 drain_right.n8 drain_right.n7 185
R911 drain_right.n125 drain_right.n124 185
R912 drain_right.n127 drain_right.n126 185
R913 drain_right.n4 drain_right.n3 185
R914 drain_right.n133 drain_right.n132 185
R915 drain_right.n135 drain_right.n134 185
R916 drain_right.n277 drain_right.n276 185
R917 drain_right.n275 drain_right.n274 185
R918 drain_right.n146 drain_right.n145 185
R919 drain_right.n269 drain_right.n268 185
R920 drain_right.n267 drain_right.n266 185
R921 drain_right.n150 drain_right.n149 185
R922 drain_right.n261 drain_right.n260 185
R923 drain_right.n259 drain_right.n258 185
R924 drain_right.n257 drain_right.n153 185
R925 drain_right.n157 drain_right.n154 185
R926 drain_right.n252 drain_right.n251 185
R927 drain_right.n250 drain_right.n249 185
R928 drain_right.n159 drain_right.n158 185
R929 drain_right.n244 drain_right.n243 185
R930 drain_right.n242 drain_right.n241 185
R931 drain_right.n163 drain_right.n162 185
R932 drain_right.n236 drain_right.n235 185
R933 drain_right.n234 drain_right.n233 185
R934 drain_right.n167 drain_right.n166 185
R935 drain_right.n228 drain_right.n227 185
R936 drain_right.n226 drain_right.n225 185
R937 drain_right.n171 drain_right.n170 185
R938 drain_right.n220 drain_right.n219 185
R939 drain_right.n218 drain_right.n217 185
R940 drain_right.n175 drain_right.n174 185
R941 drain_right.n212 drain_right.n211 185
R942 drain_right.n210 drain_right.n177 185
R943 drain_right.n209 drain_right.n208 185
R944 drain_right.n180 drain_right.n178 185
R945 drain_right.n203 drain_right.n202 185
R946 drain_right.n201 drain_right.n200 185
R947 drain_right.n184 drain_right.n183 185
R948 drain_right.n195 drain_right.n194 185
R949 drain_right.n193 drain_right.n192 185
R950 drain_right.n188 drain_right.n187 185
R951 drain_right.n45 drain_right.t3 149.524
R952 drain_right.n189 drain_right.t5 149.524
R953 drain_right.n49 drain_right.n43 104.615
R954 drain_right.n50 drain_right.n49 104.615
R955 drain_right.n50 drain_right.n39 104.615
R956 drain_right.n57 drain_right.n39 104.615
R957 drain_right.n58 drain_right.n57 104.615
R958 drain_right.n58 drain_right.n35 104.615
R959 drain_right.n66 drain_right.n35 104.615
R960 drain_right.n67 drain_right.n66 104.615
R961 drain_right.n68 drain_right.n67 104.615
R962 drain_right.n68 drain_right.n31 104.615
R963 drain_right.n75 drain_right.n31 104.615
R964 drain_right.n76 drain_right.n75 104.615
R965 drain_right.n76 drain_right.n27 104.615
R966 drain_right.n83 drain_right.n27 104.615
R967 drain_right.n84 drain_right.n83 104.615
R968 drain_right.n84 drain_right.n23 104.615
R969 drain_right.n91 drain_right.n23 104.615
R970 drain_right.n92 drain_right.n91 104.615
R971 drain_right.n92 drain_right.n19 104.615
R972 drain_right.n99 drain_right.n19 104.615
R973 drain_right.n100 drain_right.n99 104.615
R974 drain_right.n100 drain_right.n15 104.615
R975 drain_right.n107 drain_right.n15 104.615
R976 drain_right.n109 drain_right.n107 104.615
R977 drain_right.n109 drain_right.n108 104.615
R978 drain_right.n108 drain_right.n11 104.615
R979 drain_right.n117 drain_right.n11 104.615
R980 drain_right.n118 drain_right.n117 104.615
R981 drain_right.n118 drain_right.n7 104.615
R982 drain_right.n125 drain_right.n7 104.615
R983 drain_right.n126 drain_right.n125 104.615
R984 drain_right.n126 drain_right.n3 104.615
R985 drain_right.n133 drain_right.n3 104.615
R986 drain_right.n134 drain_right.n133 104.615
R987 drain_right.n276 drain_right.n275 104.615
R988 drain_right.n275 drain_right.n145 104.615
R989 drain_right.n268 drain_right.n145 104.615
R990 drain_right.n268 drain_right.n267 104.615
R991 drain_right.n267 drain_right.n149 104.615
R992 drain_right.n260 drain_right.n149 104.615
R993 drain_right.n260 drain_right.n259 104.615
R994 drain_right.n259 drain_right.n153 104.615
R995 drain_right.n157 drain_right.n153 104.615
R996 drain_right.n251 drain_right.n157 104.615
R997 drain_right.n251 drain_right.n250 104.615
R998 drain_right.n250 drain_right.n158 104.615
R999 drain_right.n243 drain_right.n158 104.615
R1000 drain_right.n243 drain_right.n242 104.615
R1001 drain_right.n242 drain_right.n162 104.615
R1002 drain_right.n235 drain_right.n162 104.615
R1003 drain_right.n235 drain_right.n234 104.615
R1004 drain_right.n234 drain_right.n166 104.615
R1005 drain_right.n227 drain_right.n166 104.615
R1006 drain_right.n227 drain_right.n226 104.615
R1007 drain_right.n226 drain_right.n170 104.615
R1008 drain_right.n219 drain_right.n170 104.615
R1009 drain_right.n219 drain_right.n218 104.615
R1010 drain_right.n218 drain_right.n174 104.615
R1011 drain_right.n211 drain_right.n174 104.615
R1012 drain_right.n211 drain_right.n210 104.615
R1013 drain_right.n210 drain_right.n209 104.615
R1014 drain_right.n209 drain_right.n178 104.615
R1015 drain_right.n202 drain_right.n178 104.615
R1016 drain_right.n202 drain_right.n201 104.615
R1017 drain_right.n201 drain_right.n183 104.615
R1018 drain_right.n194 drain_right.n183 104.615
R1019 drain_right.n194 drain_right.n193 104.615
R1020 drain_right.n193 drain_right.n187 104.615
R1021 drain_right.n281 drain_right.n141 59.2584
R1022 drain_right.n140 drain_right.n139 58.7959
R1023 drain_right.t3 drain_right.n43 52.3082
R1024 drain_right.t5 drain_right.n187 52.3082
R1025 drain_right.n140 drain_right.n138 47.6646
R1026 drain_right.n281 drain_right.n280 47.3126
R1027 drain_right drain_right.n140 38.1559
R1028 drain_right.n69 drain_right.n34 13.1884
R1029 drain_right.n116 drain_right.n115 13.1884
R1030 drain_right.n258 drain_right.n257 13.1884
R1031 drain_right.n212 drain_right.n177 13.1884
R1032 drain_right.n65 drain_right.n64 12.8005
R1033 drain_right.n70 drain_right.n32 12.8005
R1034 drain_right.n114 drain_right.n12 12.8005
R1035 drain_right.n119 drain_right.n10 12.8005
R1036 drain_right.n261 drain_right.n152 12.8005
R1037 drain_right.n256 drain_right.n154 12.8005
R1038 drain_right.n213 drain_right.n175 12.8005
R1039 drain_right.n208 drain_right.n179 12.8005
R1040 drain_right.n63 drain_right.n36 12.0247
R1041 drain_right.n74 drain_right.n73 12.0247
R1042 drain_right.n111 drain_right.n110 12.0247
R1043 drain_right.n120 drain_right.n8 12.0247
R1044 drain_right.n262 drain_right.n150 12.0247
R1045 drain_right.n253 drain_right.n252 12.0247
R1046 drain_right.n217 drain_right.n216 12.0247
R1047 drain_right.n207 drain_right.n180 12.0247
R1048 drain_right.n60 drain_right.n59 11.249
R1049 drain_right.n77 drain_right.n30 11.249
R1050 drain_right.n106 drain_right.n14 11.249
R1051 drain_right.n124 drain_right.n123 11.249
R1052 drain_right.n266 drain_right.n265 11.249
R1053 drain_right.n249 drain_right.n156 11.249
R1054 drain_right.n220 drain_right.n173 11.249
R1055 drain_right.n204 drain_right.n203 11.249
R1056 drain_right.n56 drain_right.n38 10.4732
R1057 drain_right.n78 drain_right.n28 10.4732
R1058 drain_right.n105 drain_right.n16 10.4732
R1059 drain_right.n127 drain_right.n6 10.4732
R1060 drain_right.n269 drain_right.n148 10.4732
R1061 drain_right.n248 drain_right.n159 10.4732
R1062 drain_right.n221 drain_right.n171 10.4732
R1063 drain_right.n200 drain_right.n182 10.4732
R1064 drain_right.n45 drain_right.n44 10.2747
R1065 drain_right.n189 drain_right.n188 10.2747
R1066 drain_right.n55 drain_right.n40 9.69747
R1067 drain_right.n82 drain_right.n81 9.69747
R1068 drain_right.n102 drain_right.n101 9.69747
R1069 drain_right.n128 drain_right.n4 9.69747
R1070 drain_right.n270 drain_right.n146 9.69747
R1071 drain_right.n245 drain_right.n244 9.69747
R1072 drain_right.n225 drain_right.n224 9.69747
R1073 drain_right.n199 drain_right.n184 9.69747
R1074 drain_right.n138 drain_right.n137 9.45567
R1075 drain_right.n280 drain_right.n279 9.45567
R1076 drain_right.n2 drain_right.n1 9.3005
R1077 drain_right.n131 drain_right.n130 9.3005
R1078 drain_right.n129 drain_right.n128 9.3005
R1079 drain_right.n6 drain_right.n5 9.3005
R1080 drain_right.n123 drain_right.n122 9.3005
R1081 drain_right.n121 drain_right.n120 9.3005
R1082 drain_right.n10 drain_right.n9 9.3005
R1083 drain_right.n89 drain_right.n88 9.3005
R1084 drain_right.n87 drain_right.n86 9.3005
R1085 drain_right.n26 drain_right.n25 9.3005
R1086 drain_right.n81 drain_right.n80 9.3005
R1087 drain_right.n79 drain_right.n78 9.3005
R1088 drain_right.n30 drain_right.n29 9.3005
R1089 drain_right.n73 drain_right.n72 9.3005
R1090 drain_right.n71 drain_right.n70 9.3005
R1091 drain_right.n47 drain_right.n46 9.3005
R1092 drain_right.n42 drain_right.n41 9.3005
R1093 drain_right.n53 drain_right.n52 9.3005
R1094 drain_right.n55 drain_right.n54 9.3005
R1095 drain_right.n38 drain_right.n37 9.3005
R1096 drain_right.n61 drain_right.n60 9.3005
R1097 drain_right.n63 drain_right.n62 9.3005
R1098 drain_right.n64 drain_right.n33 9.3005
R1099 drain_right.n22 drain_right.n21 9.3005
R1100 drain_right.n95 drain_right.n94 9.3005
R1101 drain_right.n97 drain_right.n96 9.3005
R1102 drain_right.n18 drain_right.n17 9.3005
R1103 drain_right.n103 drain_right.n102 9.3005
R1104 drain_right.n105 drain_right.n104 9.3005
R1105 drain_right.n14 drain_right.n13 9.3005
R1106 drain_right.n112 drain_right.n111 9.3005
R1107 drain_right.n114 drain_right.n113 9.3005
R1108 drain_right.n137 drain_right.n136 9.3005
R1109 drain_right.n191 drain_right.n190 9.3005
R1110 drain_right.n186 drain_right.n185 9.3005
R1111 drain_right.n197 drain_right.n196 9.3005
R1112 drain_right.n199 drain_right.n198 9.3005
R1113 drain_right.n182 drain_right.n181 9.3005
R1114 drain_right.n205 drain_right.n204 9.3005
R1115 drain_right.n207 drain_right.n206 9.3005
R1116 drain_right.n179 drain_right.n176 9.3005
R1117 drain_right.n238 drain_right.n237 9.3005
R1118 drain_right.n240 drain_right.n239 9.3005
R1119 drain_right.n161 drain_right.n160 9.3005
R1120 drain_right.n246 drain_right.n245 9.3005
R1121 drain_right.n248 drain_right.n247 9.3005
R1122 drain_right.n156 drain_right.n155 9.3005
R1123 drain_right.n254 drain_right.n253 9.3005
R1124 drain_right.n256 drain_right.n255 9.3005
R1125 drain_right.n279 drain_right.n278 9.3005
R1126 drain_right.n144 drain_right.n143 9.3005
R1127 drain_right.n273 drain_right.n272 9.3005
R1128 drain_right.n271 drain_right.n270 9.3005
R1129 drain_right.n148 drain_right.n147 9.3005
R1130 drain_right.n265 drain_right.n264 9.3005
R1131 drain_right.n263 drain_right.n262 9.3005
R1132 drain_right.n152 drain_right.n151 9.3005
R1133 drain_right.n165 drain_right.n164 9.3005
R1134 drain_right.n232 drain_right.n231 9.3005
R1135 drain_right.n230 drain_right.n229 9.3005
R1136 drain_right.n169 drain_right.n168 9.3005
R1137 drain_right.n224 drain_right.n223 9.3005
R1138 drain_right.n222 drain_right.n221 9.3005
R1139 drain_right.n173 drain_right.n172 9.3005
R1140 drain_right.n216 drain_right.n215 9.3005
R1141 drain_right.n214 drain_right.n213 9.3005
R1142 drain_right.n52 drain_right.n51 8.92171
R1143 drain_right.n85 drain_right.n26 8.92171
R1144 drain_right.n98 drain_right.n18 8.92171
R1145 drain_right.n132 drain_right.n131 8.92171
R1146 drain_right.n274 drain_right.n273 8.92171
R1147 drain_right.n241 drain_right.n161 8.92171
R1148 drain_right.n228 drain_right.n169 8.92171
R1149 drain_right.n196 drain_right.n195 8.92171
R1150 drain_right.n48 drain_right.n42 8.14595
R1151 drain_right.n86 drain_right.n24 8.14595
R1152 drain_right.n97 drain_right.n20 8.14595
R1153 drain_right.n135 drain_right.n2 8.14595
R1154 drain_right.n277 drain_right.n144 8.14595
R1155 drain_right.n240 drain_right.n163 8.14595
R1156 drain_right.n229 drain_right.n167 8.14595
R1157 drain_right.n192 drain_right.n186 8.14595
R1158 drain_right.n47 drain_right.n44 7.3702
R1159 drain_right.n90 drain_right.n89 7.3702
R1160 drain_right.n94 drain_right.n93 7.3702
R1161 drain_right.n136 drain_right.n0 7.3702
R1162 drain_right.n278 drain_right.n142 7.3702
R1163 drain_right.n237 drain_right.n236 7.3702
R1164 drain_right.n233 drain_right.n232 7.3702
R1165 drain_right.n191 drain_right.n188 7.3702
R1166 drain_right.n90 drain_right.n22 6.59444
R1167 drain_right.n93 drain_right.n22 6.59444
R1168 drain_right.n138 drain_right.n0 6.59444
R1169 drain_right.n280 drain_right.n142 6.59444
R1170 drain_right.n236 drain_right.n165 6.59444
R1171 drain_right.n233 drain_right.n165 6.59444
R1172 drain_right drain_right.n281 5.92477
R1173 drain_right.n48 drain_right.n47 5.81868
R1174 drain_right.n89 drain_right.n24 5.81868
R1175 drain_right.n94 drain_right.n20 5.81868
R1176 drain_right.n136 drain_right.n135 5.81868
R1177 drain_right.n278 drain_right.n277 5.81868
R1178 drain_right.n237 drain_right.n163 5.81868
R1179 drain_right.n232 drain_right.n167 5.81868
R1180 drain_right.n192 drain_right.n191 5.81868
R1181 drain_right.n51 drain_right.n42 5.04292
R1182 drain_right.n86 drain_right.n85 5.04292
R1183 drain_right.n98 drain_right.n97 5.04292
R1184 drain_right.n132 drain_right.n2 5.04292
R1185 drain_right.n274 drain_right.n144 5.04292
R1186 drain_right.n241 drain_right.n240 5.04292
R1187 drain_right.n229 drain_right.n228 5.04292
R1188 drain_right.n195 drain_right.n186 5.04292
R1189 drain_right.n52 drain_right.n40 4.26717
R1190 drain_right.n82 drain_right.n26 4.26717
R1191 drain_right.n101 drain_right.n18 4.26717
R1192 drain_right.n131 drain_right.n4 4.26717
R1193 drain_right.n273 drain_right.n146 4.26717
R1194 drain_right.n244 drain_right.n161 4.26717
R1195 drain_right.n225 drain_right.n169 4.26717
R1196 drain_right.n196 drain_right.n184 4.26717
R1197 drain_right.n56 drain_right.n55 3.49141
R1198 drain_right.n81 drain_right.n28 3.49141
R1199 drain_right.n102 drain_right.n16 3.49141
R1200 drain_right.n128 drain_right.n127 3.49141
R1201 drain_right.n270 drain_right.n269 3.49141
R1202 drain_right.n245 drain_right.n159 3.49141
R1203 drain_right.n224 drain_right.n171 3.49141
R1204 drain_right.n200 drain_right.n199 3.49141
R1205 drain_right.n190 drain_right.n189 2.84303
R1206 drain_right.n46 drain_right.n45 2.84303
R1207 drain_right.n59 drain_right.n38 2.71565
R1208 drain_right.n78 drain_right.n77 2.71565
R1209 drain_right.n106 drain_right.n105 2.71565
R1210 drain_right.n124 drain_right.n6 2.71565
R1211 drain_right.n266 drain_right.n148 2.71565
R1212 drain_right.n249 drain_right.n248 2.71565
R1213 drain_right.n221 drain_right.n220 2.71565
R1214 drain_right.n203 drain_right.n182 2.71565
R1215 drain_right.n60 drain_right.n36 1.93989
R1216 drain_right.n74 drain_right.n30 1.93989
R1217 drain_right.n110 drain_right.n14 1.93989
R1218 drain_right.n123 drain_right.n8 1.93989
R1219 drain_right.n265 drain_right.n150 1.93989
R1220 drain_right.n252 drain_right.n156 1.93989
R1221 drain_right.n217 drain_right.n173 1.93989
R1222 drain_right.n204 drain_right.n180 1.93989
R1223 drain_right.n65 drain_right.n63 1.16414
R1224 drain_right.n73 drain_right.n32 1.16414
R1225 drain_right.n111 drain_right.n12 1.16414
R1226 drain_right.n120 drain_right.n119 1.16414
R1227 drain_right.n262 drain_right.n261 1.16414
R1228 drain_right.n253 drain_right.n154 1.16414
R1229 drain_right.n216 drain_right.n175 1.16414
R1230 drain_right.n208 drain_right.n207 1.16414
R1231 drain_right.n139 drain_right.t1 0.7925
R1232 drain_right.n139 drain_right.t4 0.7925
R1233 drain_right.n141 drain_right.t0 0.7925
R1234 drain_right.n141 drain_right.t2 0.7925
R1235 drain_right.n64 drain_right.n34 0.388379
R1236 drain_right.n70 drain_right.n69 0.388379
R1237 drain_right.n115 drain_right.n114 0.388379
R1238 drain_right.n116 drain_right.n10 0.388379
R1239 drain_right.n258 drain_right.n152 0.388379
R1240 drain_right.n257 drain_right.n256 0.388379
R1241 drain_right.n213 drain_right.n212 0.388379
R1242 drain_right.n179 drain_right.n177 0.388379
R1243 drain_right.n46 drain_right.n41 0.155672
R1244 drain_right.n53 drain_right.n41 0.155672
R1245 drain_right.n54 drain_right.n53 0.155672
R1246 drain_right.n54 drain_right.n37 0.155672
R1247 drain_right.n61 drain_right.n37 0.155672
R1248 drain_right.n62 drain_right.n61 0.155672
R1249 drain_right.n62 drain_right.n33 0.155672
R1250 drain_right.n71 drain_right.n33 0.155672
R1251 drain_right.n72 drain_right.n71 0.155672
R1252 drain_right.n72 drain_right.n29 0.155672
R1253 drain_right.n79 drain_right.n29 0.155672
R1254 drain_right.n80 drain_right.n79 0.155672
R1255 drain_right.n80 drain_right.n25 0.155672
R1256 drain_right.n87 drain_right.n25 0.155672
R1257 drain_right.n88 drain_right.n87 0.155672
R1258 drain_right.n88 drain_right.n21 0.155672
R1259 drain_right.n95 drain_right.n21 0.155672
R1260 drain_right.n96 drain_right.n95 0.155672
R1261 drain_right.n96 drain_right.n17 0.155672
R1262 drain_right.n103 drain_right.n17 0.155672
R1263 drain_right.n104 drain_right.n103 0.155672
R1264 drain_right.n104 drain_right.n13 0.155672
R1265 drain_right.n112 drain_right.n13 0.155672
R1266 drain_right.n113 drain_right.n112 0.155672
R1267 drain_right.n113 drain_right.n9 0.155672
R1268 drain_right.n121 drain_right.n9 0.155672
R1269 drain_right.n122 drain_right.n121 0.155672
R1270 drain_right.n122 drain_right.n5 0.155672
R1271 drain_right.n129 drain_right.n5 0.155672
R1272 drain_right.n130 drain_right.n129 0.155672
R1273 drain_right.n130 drain_right.n1 0.155672
R1274 drain_right.n137 drain_right.n1 0.155672
R1275 drain_right.n279 drain_right.n143 0.155672
R1276 drain_right.n272 drain_right.n143 0.155672
R1277 drain_right.n272 drain_right.n271 0.155672
R1278 drain_right.n271 drain_right.n147 0.155672
R1279 drain_right.n264 drain_right.n147 0.155672
R1280 drain_right.n264 drain_right.n263 0.155672
R1281 drain_right.n263 drain_right.n151 0.155672
R1282 drain_right.n255 drain_right.n151 0.155672
R1283 drain_right.n255 drain_right.n254 0.155672
R1284 drain_right.n254 drain_right.n155 0.155672
R1285 drain_right.n247 drain_right.n155 0.155672
R1286 drain_right.n247 drain_right.n246 0.155672
R1287 drain_right.n246 drain_right.n160 0.155672
R1288 drain_right.n239 drain_right.n160 0.155672
R1289 drain_right.n239 drain_right.n238 0.155672
R1290 drain_right.n238 drain_right.n164 0.155672
R1291 drain_right.n231 drain_right.n164 0.155672
R1292 drain_right.n231 drain_right.n230 0.155672
R1293 drain_right.n230 drain_right.n168 0.155672
R1294 drain_right.n223 drain_right.n168 0.155672
R1295 drain_right.n223 drain_right.n222 0.155672
R1296 drain_right.n222 drain_right.n172 0.155672
R1297 drain_right.n215 drain_right.n172 0.155672
R1298 drain_right.n215 drain_right.n214 0.155672
R1299 drain_right.n214 drain_right.n176 0.155672
R1300 drain_right.n206 drain_right.n176 0.155672
R1301 drain_right.n206 drain_right.n205 0.155672
R1302 drain_right.n205 drain_right.n181 0.155672
R1303 drain_right.n198 drain_right.n181 0.155672
R1304 drain_right.n198 drain_right.n197 0.155672
R1305 drain_right.n197 drain_right.n185 0.155672
R1306 drain_right.n190 drain_right.n185 0.155672
R1307 plus.n0 plus.t0 2168.27
R1308 plus.n2 plus.t3 2168.27
R1309 plus.n4 plus.t4 2168.27
R1310 plus.n6 plus.t5 2168.27
R1311 plus.n1 plus.t1 2112.77
R1312 plus.n5 plus.t2 2112.77
R1313 plus.n3 plus.n0 161.489
R1314 plus.n7 plus.n4 161.489
R1315 plus.n3 plus.n2 161.3
R1316 plus.n7 plus.n6 161.3
R1317 plus.n1 plus.n0 36.5157
R1318 plus.n2 plus.n1 36.5157
R1319 plus.n6 plus.n5 36.5157
R1320 plus.n5 plus.n4 36.5157
R1321 plus plus.n7 32.5805
R1322 plus plus.n3 17.1009
R1323 drain_left.n134 drain_left.n0 289.615
R1324 drain_left.n275 drain_left.n141 289.615
R1325 drain_left.n44 drain_left.n43 185
R1326 drain_left.n49 drain_left.n48 185
R1327 drain_left.n51 drain_left.n50 185
R1328 drain_left.n40 drain_left.n39 185
R1329 drain_left.n57 drain_left.n56 185
R1330 drain_left.n59 drain_left.n58 185
R1331 drain_left.n36 drain_left.n35 185
R1332 drain_left.n66 drain_left.n65 185
R1333 drain_left.n67 drain_left.n34 185
R1334 drain_left.n69 drain_left.n68 185
R1335 drain_left.n32 drain_left.n31 185
R1336 drain_left.n75 drain_left.n74 185
R1337 drain_left.n77 drain_left.n76 185
R1338 drain_left.n28 drain_left.n27 185
R1339 drain_left.n83 drain_left.n82 185
R1340 drain_left.n85 drain_left.n84 185
R1341 drain_left.n24 drain_left.n23 185
R1342 drain_left.n91 drain_left.n90 185
R1343 drain_left.n93 drain_left.n92 185
R1344 drain_left.n20 drain_left.n19 185
R1345 drain_left.n99 drain_left.n98 185
R1346 drain_left.n101 drain_left.n100 185
R1347 drain_left.n16 drain_left.n15 185
R1348 drain_left.n107 drain_left.n106 185
R1349 drain_left.n110 drain_left.n109 185
R1350 drain_left.n108 drain_left.n12 185
R1351 drain_left.n115 drain_left.n11 185
R1352 drain_left.n117 drain_left.n116 185
R1353 drain_left.n119 drain_left.n118 185
R1354 drain_left.n8 drain_left.n7 185
R1355 drain_left.n125 drain_left.n124 185
R1356 drain_left.n127 drain_left.n126 185
R1357 drain_left.n4 drain_left.n3 185
R1358 drain_left.n133 drain_left.n132 185
R1359 drain_left.n135 drain_left.n134 185
R1360 drain_left.n276 drain_left.n275 185
R1361 drain_left.n274 drain_left.n273 185
R1362 drain_left.n145 drain_left.n144 185
R1363 drain_left.n268 drain_left.n267 185
R1364 drain_left.n266 drain_left.n265 185
R1365 drain_left.n149 drain_left.n148 185
R1366 drain_left.n260 drain_left.n259 185
R1367 drain_left.n258 drain_left.n257 185
R1368 drain_left.n256 drain_left.n152 185
R1369 drain_left.n156 drain_left.n153 185
R1370 drain_left.n251 drain_left.n250 185
R1371 drain_left.n249 drain_left.n248 185
R1372 drain_left.n158 drain_left.n157 185
R1373 drain_left.n243 drain_left.n242 185
R1374 drain_left.n241 drain_left.n240 185
R1375 drain_left.n162 drain_left.n161 185
R1376 drain_left.n235 drain_left.n234 185
R1377 drain_left.n233 drain_left.n232 185
R1378 drain_left.n166 drain_left.n165 185
R1379 drain_left.n227 drain_left.n226 185
R1380 drain_left.n225 drain_left.n224 185
R1381 drain_left.n170 drain_left.n169 185
R1382 drain_left.n219 drain_left.n218 185
R1383 drain_left.n217 drain_left.n216 185
R1384 drain_left.n174 drain_left.n173 185
R1385 drain_left.n211 drain_left.n210 185
R1386 drain_left.n209 drain_left.n176 185
R1387 drain_left.n208 drain_left.n207 185
R1388 drain_left.n179 drain_left.n177 185
R1389 drain_left.n202 drain_left.n201 185
R1390 drain_left.n200 drain_left.n199 185
R1391 drain_left.n183 drain_left.n182 185
R1392 drain_left.n194 drain_left.n193 185
R1393 drain_left.n192 drain_left.n191 185
R1394 drain_left.n187 drain_left.n186 185
R1395 drain_left.n45 drain_left.t0 149.524
R1396 drain_left.n188 drain_left.t5 149.524
R1397 drain_left.n49 drain_left.n43 104.615
R1398 drain_left.n50 drain_left.n49 104.615
R1399 drain_left.n50 drain_left.n39 104.615
R1400 drain_left.n57 drain_left.n39 104.615
R1401 drain_left.n58 drain_left.n57 104.615
R1402 drain_left.n58 drain_left.n35 104.615
R1403 drain_left.n66 drain_left.n35 104.615
R1404 drain_left.n67 drain_left.n66 104.615
R1405 drain_left.n68 drain_left.n67 104.615
R1406 drain_left.n68 drain_left.n31 104.615
R1407 drain_left.n75 drain_left.n31 104.615
R1408 drain_left.n76 drain_left.n75 104.615
R1409 drain_left.n76 drain_left.n27 104.615
R1410 drain_left.n83 drain_left.n27 104.615
R1411 drain_left.n84 drain_left.n83 104.615
R1412 drain_left.n84 drain_left.n23 104.615
R1413 drain_left.n91 drain_left.n23 104.615
R1414 drain_left.n92 drain_left.n91 104.615
R1415 drain_left.n92 drain_left.n19 104.615
R1416 drain_left.n99 drain_left.n19 104.615
R1417 drain_left.n100 drain_left.n99 104.615
R1418 drain_left.n100 drain_left.n15 104.615
R1419 drain_left.n107 drain_left.n15 104.615
R1420 drain_left.n109 drain_left.n107 104.615
R1421 drain_left.n109 drain_left.n108 104.615
R1422 drain_left.n108 drain_left.n11 104.615
R1423 drain_left.n117 drain_left.n11 104.615
R1424 drain_left.n118 drain_left.n117 104.615
R1425 drain_left.n118 drain_left.n7 104.615
R1426 drain_left.n125 drain_left.n7 104.615
R1427 drain_left.n126 drain_left.n125 104.615
R1428 drain_left.n126 drain_left.n3 104.615
R1429 drain_left.n133 drain_left.n3 104.615
R1430 drain_left.n134 drain_left.n133 104.615
R1431 drain_left.n275 drain_left.n274 104.615
R1432 drain_left.n274 drain_left.n144 104.615
R1433 drain_left.n267 drain_left.n144 104.615
R1434 drain_left.n267 drain_left.n266 104.615
R1435 drain_left.n266 drain_left.n148 104.615
R1436 drain_left.n259 drain_left.n148 104.615
R1437 drain_left.n259 drain_left.n258 104.615
R1438 drain_left.n258 drain_left.n152 104.615
R1439 drain_left.n156 drain_left.n152 104.615
R1440 drain_left.n250 drain_left.n156 104.615
R1441 drain_left.n250 drain_left.n249 104.615
R1442 drain_left.n249 drain_left.n157 104.615
R1443 drain_left.n242 drain_left.n157 104.615
R1444 drain_left.n242 drain_left.n241 104.615
R1445 drain_left.n241 drain_left.n161 104.615
R1446 drain_left.n234 drain_left.n161 104.615
R1447 drain_left.n234 drain_left.n233 104.615
R1448 drain_left.n233 drain_left.n165 104.615
R1449 drain_left.n226 drain_left.n165 104.615
R1450 drain_left.n226 drain_left.n225 104.615
R1451 drain_left.n225 drain_left.n169 104.615
R1452 drain_left.n218 drain_left.n169 104.615
R1453 drain_left.n218 drain_left.n217 104.615
R1454 drain_left.n217 drain_left.n173 104.615
R1455 drain_left.n210 drain_left.n173 104.615
R1456 drain_left.n210 drain_left.n209 104.615
R1457 drain_left.n209 drain_left.n208 104.615
R1458 drain_left.n208 drain_left.n177 104.615
R1459 drain_left.n201 drain_left.n177 104.615
R1460 drain_left.n201 drain_left.n200 104.615
R1461 drain_left.n200 drain_left.n182 104.615
R1462 drain_left.n193 drain_left.n182 104.615
R1463 drain_left.n193 drain_left.n192 104.615
R1464 drain_left.n192 drain_left.n186 104.615
R1465 drain_left.n140 drain_left.n139 58.7959
R1466 drain_left.n281 drain_left.n280 58.7153
R1467 drain_left.t0 drain_left.n43 52.3082
R1468 drain_left.t5 drain_left.n186 52.3082
R1469 drain_left.n281 drain_left.n279 47.8557
R1470 drain_left.n140 drain_left.n138 47.6646
R1471 drain_left drain_left.n140 38.7091
R1472 drain_left.n69 drain_left.n34 13.1884
R1473 drain_left.n116 drain_left.n115 13.1884
R1474 drain_left.n257 drain_left.n256 13.1884
R1475 drain_left.n211 drain_left.n176 13.1884
R1476 drain_left.n65 drain_left.n64 12.8005
R1477 drain_left.n70 drain_left.n32 12.8005
R1478 drain_left.n114 drain_left.n12 12.8005
R1479 drain_left.n119 drain_left.n10 12.8005
R1480 drain_left.n260 drain_left.n151 12.8005
R1481 drain_left.n255 drain_left.n153 12.8005
R1482 drain_left.n212 drain_left.n174 12.8005
R1483 drain_left.n207 drain_left.n178 12.8005
R1484 drain_left.n63 drain_left.n36 12.0247
R1485 drain_left.n74 drain_left.n73 12.0247
R1486 drain_left.n111 drain_left.n110 12.0247
R1487 drain_left.n120 drain_left.n8 12.0247
R1488 drain_left.n261 drain_left.n149 12.0247
R1489 drain_left.n252 drain_left.n251 12.0247
R1490 drain_left.n216 drain_left.n215 12.0247
R1491 drain_left.n206 drain_left.n179 12.0247
R1492 drain_left.n60 drain_left.n59 11.249
R1493 drain_left.n77 drain_left.n30 11.249
R1494 drain_left.n106 drain_left.n14 11.249
R1495 drain_left.n124 drain_left.n123 11.249
R1496 drain_left.n265 drain_left.n264 11.249
R1497 drain_left.n248 drain_left.n155 11.249
R1498 drain_left.n219 drain_left.n172 11.249
R1499 drain_left.n203 drain_left.n202 11.249
R1500 drain_left.n56 drain_left.n38 10.4732
R1501 drain_left.n78 drain_left.n28 10.4732
R1502 drain_left.n105 drain_left.n16 10.4732
R1503 drain_left.n127 drain_left.n6 10.4732
R1504 drain_left.n268 drain_left.n147 10.4732
R1505 drain_left.n247 drain_left.n158 10.4732
R1506 drain_left.n220 drain_left.n170 10.4732
R1507 drain_left.n199 drain_left.n181 10.4732
R1508 drain_left.n45 drain_left.n44 10.2747
R1509 drain_left.n188 drain_left.n187 10.2747
R1510 drain_left.n55 drain_left.n40 9.69747
R1511 drain_left.n82 drain_left.n81 9.69747
R1512 drain_left.n102 drain_left.n101 9.69747
R1513 drain_left.n128 drain_left.n4 9.69747
R1514 drain_left.n269 drain_left.n145 9.69747
R1515 drain_left.n244 drain_left.n243 9.69747
R1516 drain_left.n224 drain_left.n223 9.69747
R1517 drain_left.n198 drain_left.n183 9.69747
R1518 drain_left.n138 drain_left.n137 9.45567
R1519 drain_left.n279 drain_left.n278 9.45567
R1520 drain_left.n2 drain_left.n1 9.3005
R1521 drain_left.n131 drain_left.n130 9.3005
R1522 drain_left.n129 drain_left.n128 9.3005
R1523 drain_left.n6 drain_left.n5 9.3005
R1524 drain_left.n123 drain_left.n122 9.3005
R1525 drain_left.n121 drain_left.n120 9.3005
R1526 drain_left.n10 drain_left.n9 9.3005
R1527 drain_left.n89 drain_left.n88 9.3005
R1528 drain_left.n87 drain_left.n86 9.3005
R1529 drain_left.n26 drain_left.n25 9.3005
R1530 drain_left.n81 drain_left.n80 9.3005
R1531 drain_left.n79 drain_left.n78 9.3005
R1532 drain_left.n30 drain_left.n29 9.3005
R1533 drain_left.n73 drain_left.n72 9.3005
R1534 drain_left.n71 drain_left.n70 9.3005
R1535 drain_left.n47 drain_left.n46 9.3005
R1536 drain_left.n42 drain_left.n41 9.3005
R1537 drain_left.n53 drain_left.n52 9.3005
R1538 drain_left.n55 drain_left.n54 9.3005
R1539 drain_left.n38 drain_left.n37 9.3005
R1540 drain_left.n61 drain_left.n60 9.3005
R1541 drain_left.n63 drain_left.n62 9.3005
R1542 drain_left.n64 drain_left.n33 9.3005
R1543 drain_left.n22 drain_left.n21 9.3005
R1544 drain_left.n95 drain_left.n94 9.3005
R1545 drain_left.n97 drain_left.n96 9.3005
R1546 drain_left.n18 drain_left.n17 9.3005
R1547 drain_left.n103 drain_left.n102 9.3005
R1548 drain_left.n105 drain_left.n104 9.3005
R1549 drain_left.n14 drain_left.n13 9.3005
R1550 drain_left.n112 drain_left.n111 9.3005
R1551 drain_left.n114 drain_left.n113 9.3005
R1552 drain_left.n137 drain_left.n136 9.3005
R1553 drain_left.n190 drain_left.n189 9.3005
R1554 drain_left.n185 drain_left.n184 9.3005
R1555 drain_left.n196 drain_left.n195 9.3005
R1556 drain_left.n198 drain_left.n197 9.3005
R1557 drain_left.n181 drain_left.n180 9.3005
R1558 drain_left.n204 drain_left.n203 9.3005
R1559 drain_left.n206 drain_left.n205 9.3005
R1560 drain_left.n178 drain_left.n175 9.3005
R1561 drain_left.n237 drain_left.n236 9.3005
R1562 drain_left.n239 drain_left.n238 9.3005
R1563 drain_left.n160 drain_left.n159 9.3005
R1564 drain_left.n245 drain_left.n244 9.3005
R1565 drain_left.n247 drain_left.n246 9.3005
R1566 drain_left.n155 drain_left.n154 9.3005
R1567 drain_left.n253 drain_left.n252 9.3005
R1568 drain_left.n255 drain_left.n254 9.3005
R1569 drain_left.n278 drain_left.n277 9.3005
R1570 drain_left.n143 drain_left.n142 9.3005
R1571 drain_left.n272 drain_left.n271 9.3005
R1572 drain_left.n270 drain_left.n269 9.3005
R1573 drain_left.n147 drain_left.n146 9.3005
R1574 drain_left.n264 drain_left.n263 9.3005
R1575 drain_left.n262 drain_left.n261 9.3005
R1576 drain_left.n151 drain_left.n150 9.3005
R1577 drain_left.n164 drain_left.n163 9.3005
R1578 drain_left.n231 drain_left.n230 9.3005
R1579 drain_left.n229 drain_left.n228 9.3005
R1580 drain_left.n168 drain_left.n167 9.3005
R1581 drain_left.n223 drain_left.n222 9.3005
R1582 drain_left.n221 drain_left.n220 9.3005
R1583 drain_left.n172 drain_left.n171 9.3005
R1584 drain_left.n215 drain_left.n214 9.3005
R1585 drain_left.n213 drain_left.n212 9.3005
R1586 drain_left.n52 drain_left.n51 8.92171
R1587 drain_left.n85 drain_left.n26 8.92171
R1588 drain_left.n98 drain_left.n18 8.92171
R1589 drain_left.n132 drain_left.n131 8.92171
R1590 drain_left.n273 drain_left.n272 8.92171
R1591 drain_left.n240 drain_left.n160 8.92171
R1592 drain_left.n227 drain_left.n168 8.92171
R1593 drain_left.n195 drain_left.n194 8.92171
R1594 drain_left.n48 drain_left.n42 8.14595
R1595 drain_left.n86 drain_left.n24 8.14595
R1596 drain_left.n97 drain_left.n20 8.14595
R1597 drain_left.n135 drain_left.n2 8.14595
R1598 drain_left.n276 drain_left.n143 8.14595
R1599 drain_left.n239 drain_left.n162 8.14595
R1600 drain_left.n228 drain_left.n166 8.14595
R1601 drain_left.n191 drain_left.n185 8.14595
R1602 drain_left.n47 drain_left.n44 7.3702
R1603 drain_left.n90 drain_left.n89 7.3702
R1604 drain_left.n94 drain_left.n93 7.3702
R1605 drain_left.n136 drain_left.n0 7.3702
R1606 drain_left.n277 drain_left.n141 7.3702
R1607 drain_left.n236 drain_left.n235 7.3702
R1608 drain_left.n232 drain_left.n231 7.3702
R1609 drain_left.n190 drain_left.n187 7.3702
R1610 drain_left.n90 drain_left.n22 6.59444
R1611 drain_left.n93 drain_left.n22 6.59444
R1612 drain_left.n138 drain_left.n0 6.59444
R1613 drain_left.n279 drain_left.n141 6.59444
R1614 drain_left.n235 drain_left.n164 6.59444
R1615 drain_left.n232 drain_left.n164 6.59444
R1616 drain_left drain_left.n281 6.19632
R1617 drain_left.n48 drain_left.n47 5.81868
R1618 drain_left.n89 drain_left.n24 5.81868
R1619 drain_left.n94 drain_left.n20 5.81868
R1620 drain_left.n136 drain_left.n135 5.81868
R1621 drain_left.n277 drain_left.n276 5.81868
R1622 drain_left.n236 drain_left.n162 5.81868
R1623 drain_left.n231 drain_left.n166 5.81868
R1624 drain_left.n191 drain_left.n190 5.81868
R1625 drain_left.n51 drain_left.n42 5.04292
R1626 drain_left.n86 drain_left.n85 5.04292
R1627 drain_left.n98 drain_left.n97 5.04292
R1628 drain_left.n132 drain_left.n2 5.04292
R1629 drain_left.n273 drain_left.n143 5.04292
R1630 drain_left.n240 drain_left.n239 5.04292
R1631 drain_left.n228 drain_left.n227 5.04292
R1632 drain_left.n194 drain_left.n185 5.04292
R1633 drain_left.n52 drain_left.n40 4.26717
R1634 drain_left.n82 drain_left.n26 4.26717
R1635 drain_left.n101 drain_left.n18 4.26717
R1636 drain_left.n131 drain_left.n4 4.26717
R1637 drain_left.n272 drain_left.n145 4.26717
R1638 drain_left.n243 drain_left.n160 4.26717
R1639 drain_left.n224 drain_left.n168 4.26717
R1640 drain_left.n195 drain_left.n183 4.26717
R1641 drain_left.n56 drain_left.n55 3.49141
R1642 drain_left.n81 drain_left.n28 3.49141
R1643 drain_left.n102 drain_left.n16 3.49141
R1644 drain_left.n128 drain_left.n127 3.49141
R1645 drain_left.n269 drain_left.n268 3.49141
R1646 drain_left.n244 drain_left.n158 3.49141
R1647 drain_left.n223 drain_left.n170 3.49141
R1648 drain_left.n199 drain_left.n198 3.49141
R1649 drain_left.n189 drain_left.n188 2.84303
R1650 drain_left.n46 drain_left.n45 2.84303
R1651 drain_left.n59 drain_left.n38 2.71565
R1652 drain_left.n78 drain_left.n77 2.71565
R1653 drain_left.n106 drain_left.n105 2.71565
R1654 drain_left.n124 drain_left.n6 2.71565
R1655 drain_left.n265 drain_left.n147 2.71565
R1656 drain_left.n248 drain_left.n247 2.71565
R1657 drain_left.n220 drain_left.n219 2.71565
R1658 drain_left.n202 drain_left.n181 2.71565
R1659 drain_left.n60 drain_left.n36 1.93989
R1660 drain_left.n74 drain_left.n30 1.93989
R1661 drain_left.n110 drain_left.n14 1.93989
R1662 drain_left.n123 drain_left.n8 1.93989
R1663 drain_left.n264 drain_left.n149 1.93989
R1664 drain_left.n251 drain_left.n155 1.93989
R1665 drain_left.n216 drain_left.n172 1.93989
R1666 drain_left.n203 drain_left.n179 1.93989
R1667 drain_left.n65 drain_left.n63 1.16414
R1668 drain_left.n73 drain_left.n32 1.16414
R1669 drain_left.n111 drain_left.n12 1.16414
R1670 drain_left.n120 drain_left.n119 1.16414
R1671 drain_left.n261 drain_left.n260 1.16414
R1672 drain_left.n252 drain_left.n153 1.16414
R1673 drain_left.n215 drain_left.n174 1.16414
R1674 drain_left.n207 drain_left.n206 1.16414
R1675 drain_left.n139 drain_left.t3 0.7925
R1676 drain_left.n139 drain_left.t1 0.7925
R1677 drain_left.n280 drain_left.t4 0.7925
R1678 drain_left.n280 drain_left.t2 0.7925
R1679 drain_left.n64 drain_left.n34 0.388379
R1680 drain_left.n70 drain_left.n69 0.388379
R1681 drain_left.n115 drain_left.n114 0.388379
R1682 drain_left.n116 drain_left.n10 0.388379
R1683 drain_left.n257 drain_left.n151 0.388379
R1684 drain_left.n256 drain_left.n255 0.388379
R1685 drain_left.n212 drain_left.n211 0.388379
R1686 drain_left.n178 drain_left.n176 0.388379
R1687 drain_left.n46 drain_left.n41 0.155672
R1688 drain_left.n53 drain_left.n41 0.155672
R1689 drain_left.n54 drain_left.n53 0.155672
R1690 drain_left.n54 drain_left.n37 0.155672
R1691 drain_left.n61 drain_left.n37 0.155672
R1692 drain_left.n62 drain_left.n61 0.155672
R1693 drain_left.n62 drain_left.n33 0.155672
R1694 drain_left.n71 drain_left.n33 0.155672
R1695 drain_left.n72 drain_left.n71 0.155672
R1696 drain_left.n72 drain_left.n29 0.155672
R1697 drain_left.n79 drain_left.n29 0.155672
R1698 drain_left.n80 drain_left.n79 0.155672
R1699 drain_left.n80 drain_left.n25 0.155672
R1700 drain_left.n87 drain_left.n25 0.155672
R1701 drain_left.n88 drain_left.n87 0.155672
R1702 drain_left.n88 drain_left.n21 0.155672
R1703 drain_left.n95 drain_left.n21 0.155672
R1704 drain_left.n96 drain_left.n95 0.155672
R1705 drain_left.n96 drain_left.n17 0.155672
R1706 drain_left.n103 drain_left.n17 0.155672
R1707 drain_left.n104 drain_left.n103 0.155672
R1708 drain_left.n104 drain_left.n13 0.155672
R1709 drain_left.n112 drain_left.n13 0.155672
R1710 drain_left.n113 drain_left.n112 0.155672
R1711 drain_left.n113 drain_left.n9 0.155672
R1712 drain_left.n121 drain_left.n9 0.155672
R1713 drain_left.n122 drain_left.n121 0.155672
R1714 drain_left.n122 drain_left.n5 0.155672
R1715 drain_left.n129 drain_left.n5 0.155672
R1716 drain_left.n130 drain_left.n129 0.155672
R1717 drain_left.n130 drain_left.n1 0.155672
R1718 drain_left.n137 drain_left.n1 0.155672
R1719 drain_left.n278 drain_left.n142 0.155672
R1720 drain_left.n271 drain_left.n142 0.155672
R1721 drain_left.n271 drain_left.n270 0.155672
R1722 drain_left.n270 drain_left.n146 0.155672
R1723 drain_left.n263 drain_left.n146 0.155672
R1724 drain_left.n263 drain_left.n262 0.155672
R1725 drain_left.n262 drain_left.n150 0.155672
R1726 drain_left.n254 drain_left.n150 0.155672
R1727 drain_left.n254 drain_left.n253 0.155672
R1728 drain_left.n253 drain_left.n154 0.155672
R1729 drain_left.n246 drain_left.n154 0.155672
R1730 drain_left.n246 drain_left.n245 0.155672
R1731 drain_left.n245 drain_left.n159 0.155672
R1732 drain_left.n238 drain_left.n159 0.155672
R1733 drain_left.n238 drain_left.n237 0.155672
R1734 drain_left.n237 drain_left.n163 0.155672
R1735 drain_left.n230 drain_left.n163 0.155672
R1736 drain_left.n230 drain_left.n229 0.155672
R1737 drain_left.n229 drain_left.n167 0.155672
R1738 drain_left.n222 drain_left.n167 0.155672
R1739 drain_left.n222 drain_left.n221 0.155672
R1740 drain_left.n221 drain_left.n171 0.155672
R1741 drain_left.n214 drain_left.n171 0.155672
R1742 drain_left.n214 drain_left.n213 0.155672
R1743 drain_left.n213 drain_left.n175 0.155672
R1744 drain_left.n205 drain_left.n175 0.155672
R1745 drain_left.n205 drain_left.n204 0.155672
R1746 drain_left.n204 drain_left.n180 0.155672
R1747 drain_left.n197 drain_left.n180 0.155672
R1748 drain_left.n197 drain_left.n196 0.155672
R1749 drain_left.n196 drain_left.n184 0.155672
R1750 drain_left.n189 drain_left.n184 0.155672
C0 source drain_right 27.529099f
C1 minus plus 7.0757f
C2 minus source 4.30867f
C3 plus source 4.324069f
C4 drain_left drain_right 0.574239f
C5 minus drain_left 0.17071f
C6 plus drain_left 5.46359f
C7 source drain_left 27.5513f
C8 minus drain_right 5.35531f
C9 plus drain_right 0.272105f
C10 drain_right a_n1220_n5888# 10.09813f
C11 drain_left a_n1220_n5888# 10.2974f
C12 source a_n1220_n5888# 10.704732f
C13 minus a_n1220_n5888# 5.536969f
C14 plus a_n1220_n5888# 8.587561f
C15 drain_left.n0 a_n1220_n5888# 0.03855f
C16 drain_left.n1 a_n1220_n5888# 0.027963f
C17 drain_left.n2 a_n1220_n5888# 0.015026f
C18 drain_left.n3 a_n1220_n5888# 0.035516f
C19 drain_left.n4 a_n1220_n5888# 0.01591f
C20 drain_left.n5 a_n1220_n5888# 0.027963f
C21 drain_left.n6 a_n1220_n5888# 0.015026f
C22 drain_left.n7 a_n1220_n5888# 0.035516f
C23 drain_left.n8 a_n1220_n5888# 0.01591f
C24 drain_left.n9 a_n1220_n5888# 0.027963f
C25 drain_left.n10 a_n1220_n5888# 0.015026f
C26 drain_left.n11 a_n1220_n5888# 0.035516f
C27 drain_left.n12 a_n1220_n5888# 0.01591f
C28 drain_left.n13 a_n1220_n5888# 0.027963f
C29 drain_left.n14 a_n1220_n5888# 0.015026f
C30 drain_left.n15 a_n1220_n5888# 0.035516f
C31 drain_left.n16 a_n1220_n5888# 0.01591f
C32 drain_left.n17 a_n1220_n5888# 0.027963f
C33 drain_left.n18 a_n1220_n5888# 0.015026f
C34 drain_left.n19 a_n1220_n5888# 0.035516f
C35 drain_left.n20 a_n1220_n5888# 0.01591f
C36 drain_left.n21 a_n1220_n5888# 0.027963f
C37 drain_left.n22 a_n1220_n5888# 0.015026f
C38 drain_left.n23 a_n1220_n5888# 0.035516f
C39 drain_left.n24 a_n1220_n5888# 0.01591f
C40 drain_left.n25 a_n1220_n5888# 0.027963f
C41 drain_left.n26 a_n1220_n5888# 0.015026f
C42 drain_left.n27 a_n1220_n5888# 0.035516f
C43 drain_left.n28 a_n1220_n5888# 0.01591f
C44 drain_left.n29 a_n1220_n5888# 0.027963f
C45 drain_left.n30 a_n1220_n5888# 0.015026f
C46 drain_left.n31 a_n1220_n5888# 0.035516f
C47 drain_left.n32 a_n1220_n5888# 0.01591f
C48 drain_left.n33 a_n1220_n5888# 0.027963f
C49 drain_left.n34 a_n1220_n5888# 0.015468f
C50 drain_left.n35 a_n1220_n5888# 0.035516f
C51 drain_left.n36 a_n1220_n5888# 0.01591f
C52 drain_left.n37 a_n1220_n5888# 0.027963f
C53 drain_left.n38 a_n1220_n5888# 0.015026f
C54 drain_left.n39 a_n1220_n5888# 0.035516f
C55 drain_left.n40 a_n1220_n5888# 0.01591f
C56 drain_left.n41 a_n1220_n5888# 0.027963f
C57 drain_left.n42 a_n1220_n5888# 0.015026f
C58 drain_left.n43 a_n1220_n5888# 0.026637f
C59 drain_left.n44 a_n1220_n5888# 0.025107f
C60 drain_left.t0 a_n1220_n5888# 0.061942f
C61 drain_left.n45 a_n1220_n5888# 0.34117f
C62 drain_left.n46 a_n1220_n5888# 3.02755f
C63 drain_left.n47 a_n1220_n5888# 0.015026f
C64 drain_left.n48 a_n1220_n5888# 0.01591f
C65 drain_left.n49 a_n1220_n5888# 0.035516f
C66 drain_left.n50 a_n1220_n5888# 0.035516f
C67 drain_left.n51 a_n1220_n5888# 0.01591f
C68 drain_left.n52 a_n1220_n5888# 0.015026f
C69 drain_left.n53 a_n1220_n5888# 0.027963f
C70 drain_left.n54 a_n1220_n5888# 0.027963f
C71 drain_left.n55 a_n1220_n5888# 0.015026f
C72 drain_left.n56 a_n1220_n5888# 0.01591f
C73 drain_left.n57 a_n1220_n5888# 0.035516f
C74 drain_left.n58 a_n1220_n5888# 0.035516f
C75 drain_left.n59 a_n1220_n5888# 0.01591f
C76 drain_left.n60 a_n1220_n5888# 0.015026f
C77 drain_left.n61 a_n1220_n5888# 0.027963f
C78 drain_left.n62 a_n1220_n5888# 0.027963f
C79 drain_left.n63 a_n1220_n5888# 0.015026f
C80 drain_left.n64 a_n1220_n5888# 0.015026f
C81 drain_left.n65 a_n1220_n5888# 0.01591f
C82 drain_left.n66 a_n1220_n5888# 0.035516f
C83 drain_left.n67 a_n1220_n5888# 0.035516f
C84 drain_left.n68 a_n1220_n5888# 0.035516f
C85 drain_left.n69 a_n1220_n5888# 0.015468f
C86 drain_left.n70 a_n1220_n5888# 0.015026f
C87 drain_left.n71 a_n1220_n5888# 0.027963f
C88 drain_left.n72 a_n1220_n5888# 0.027963f
C89 drain_left.n73 a_n1220_n5888# 0.015026f
C90 drain_left.n74 a_n1220_n5888# 0.01591f
C91 drain_left.n75 a_n1220_n5888# 0.035516f
C92 drain_left.n76 a_n1220_n5888# 0.035516f
C93 drain_left.n77 a_n1220_n5888# 0.01591f
C94 drain_left.n78 a_n1220_n5888# 0.015026f
C95 drain_left.n79 a_n1220_n5888# 0.027963f
C96 drain_left.n80 a_n1220_n5888# 0.027963f
C97 drain_left.n81 a_n1220_n5888# 0.015026f
C98 drain_left.n82 a_n1220_n5888# 0.01591f
C99 drain_left.n83 a_n1220_n5888# 0.035516f
C100 drain_left.n84 a_n1220_n5888# 0.035516f
C101 drain_left.n85 a_n1220_n5888# 0.01591f
C102 drain_left.n86 a_n1220_n5888# 0.015026f
C103 drain_left.n87 a_n1220_n5888# 0.027963f
C104 drain_left.n88 a_n1220_n5888# 0.027963f
C105 drain_left.n89 a_n1220_n5888# 0.015026f
C106 drain_left.n90 a_n1220_n5888# 0.01591f
C107 drain_left.n91 a_n1220_n5888# 0.035516f
C108 drain_left.n92 a_n1220_n5888# 0.035516f
C109 drain_left.n93 a_n1220_n5888# 0.01591f
C110 drain_left.n94 a_n1220_n5888# 0.015026f
C111 drain_left.n95 a_n1220_n5888# 0.027963f
C112 drain_left.n96 a_n1220_n5888# 0.027963f
C113 drain_left.n97 a_n1220_n5888# 0.015026f
C114 drain_left.n98 a_n1220_n5888# 0.01591f
C115 drain_left.n99 a_n1220_n5888# 0.035516f
C116 drain_left.n100 a_n1220_n5888# 0.035516f
C117 drain_left.n101 a_n1220_n5888# 0.01591f
C118 drain_left.n102 a_n1220_n5888# 0.015026f
C119 drain_left.n103 a_n1220_n5888# 0.027963f
C120 drain_left.n104 a_n1220_n5888# 0.027963f
C121 drain_left.n105 a_n1220_n5888# 0.015026f
C122 drain_left.n106 a_n1220_n5888# 0.01591f
C123 drain_left.n107 a_n1220_n5888# 0.035516f
C124 drain_left.n108 a_n1220_n5888# 0.035516f
C125 drain_left.n109 a_n1220_n5888# 0.035516f
C126 drain_left.n110 a_n1220_n5888# 0.01591f
C127 drain_left.n111 a_n1220_n5888# 0.015026f
C128 drain_left.n112 a_n1220_n5888# 0.027963f
C129 drain_left.n113 a_n1220_n5888# 0.027963f
C130 drain_left.n114 a_n1220_n5888# 0.015026f
C131 drain_left.n115 a_n1220_n5888# 0.015468f
C132 drain_left.n116 a_n1220_n5888# 0.015468f
C133 drain_left.n117 a_n1220_n5888# 0.035516f
C134 drain_left.n118 a_n1220_n5888# 0.035516f
C135 drain_left.n119 a_n1220_n5888# 0.01591f
C136 drain_left.n120 a_n1220_n5888# 0.015026f
C137 drain_left.n121 a_n1220_n5888# 0.027963f
C138 drain_left.n122 a_n1220_n5888# 0.027963f
C139 drain_left.n123 a_n1220_n5888# 0.015026f
C140 drain_left.n124 a_n1220_n5888# 0.01591f
C141 drain_left.n125 a_n1220_n5888# 0.035516f
C142 drain_left.n126 a_n1220_n5888# 0.035516f
C143 drain_left.n127 a_n1220_n5888# 0.01591f
C144 drain_left.n128 a_n1220_n5888# 0.015026f
C145 drain_left.n129 a_n1220_n5888# 0.027963f
C146 drain_left.n130 a_n1220_n5888# 0.027963f
C147 drain_left.n131 a_n1220_n5888# 0.015026f
C148 drain_left.n132 a_n1220_n5888# 0.01591f
C149 drain_left.n133 a_n1220_n5888# 0.035516f
C150 drain_left.n134 a_n1220_n5888# 0.075552f
C151 drain_left.n135 a_n1220_n5888# 0.01591f
C152 drain_left.n136 a_n1220_n5888# 0.015026f
C153 drain_left.n137 a_n1220_n5888# 0.061579f
C154 drain_left.n138 a_n1220_n5888# 0.062007f
C155 drain_left.t3 a_n1220_n5888# 0.552427f
C156 drain_left.t1 a_n1220_n5888# 0.552427f
C157 drain_left.n139 a_n1220_n5888# 5.09164f
C158 drain_left.n140 a_n1220_n5888# 2.49836f
C159 drain_left.n141 a_n1220_n5888# 0.03855f
C160 drain_left.n142 a_n1220_n5888# 0.027963f
C161 drain_left.n143 a_n1220_n5888# 0.015026f
C162 drain_left.n144 a_n1220_n5888# 0.035516f
C163 drain_left.n145 a_n1220_n5888# 0.01591f
C164 drain_left.n146 a_n1220_n5888# 0.027963f
C165 drain_left.n147 a_n1220_n5888# 0.015026f
C166 drain_left.n148 a_n1220_n5888# 0.035516f
C167 drain_left.n149 a_n1220_n5888# 0.01591f
C168 drain_left.n150 a_n1220_n5888# 0.027963f
C169 drain_left.n151 a_n1220_n5888# 0.015026f
C170 drain_left.n152 a_n1220_n5888# 0.035516f
C171 drain_left.n153 a_n1220_n5888# 0.01591f
C172 drain_left.n154 a_n1220_n5888# 0.027963f
C173 drain_left.n155 a_n1220_n5888# 0.015026f
C174 drain_left.n156 a_n1220_n5888# 0.035516f
C175 drain_left.n157 a_n1220_n5888# 0.035516f
C176 drain_left.n158 a_n1220_n5888# 0.01591f
C177 drain_left.n159 a_n1220_n5888# 0.027963f
C178 drain_left.n160 a_n1220_n5888# 0.015026f
C179 drain_left.n161 a_n1220_n5888# 0.035516f
C180 drain_left.n162 a_n1220_n5888# 0.01591f
C181 drain_left.n163 a_n1220_n5888# 0.027963f
C182 drain_left.n164 a_n1220_n5888# 0.015026f
C183 drain_left.n165 a_n1220_n5888# 0.035516f
C184 drain_left.n166 a_n1220_n5888# 0.01591f
C185 drain_left.n167 a_n1220_n5888# 0.027963f
C186 drain_left.n168 a_n1220_n5888# 0.015026f
C187 drain_left.n169 a_n1220_n5888# 0.035516f
C188 drain_left.n170 a_n1220_n5888# 0.01591f
C189 drain_left.n171 a_n1220_n5888# 0.027963f
C190 drain_left.n172 a_n1220_n5888# 0.015026f
C191 drain_left.n173 a_n1220_n5888# 0.035516f
C192 drain_left.n174 a_n1220_n5888# 0.01591f
C193 drain_left.n175 a_n1220_n5888# 0.027963f
C194 drain_left.n176 a_n1220_n5888# 0.015468f
C195 drain_left.n177 a_n1220_n5888# 0.035516f
C196 drain_left.n178 a_n1220_n5888# 0.015026f
C197 drain_left.n179 a_n1220_n5888# 0.01591f
C198 drain_left.n180 a_n1220_n5888# 0.027963f
C199 drain_left.n181 a_n1220_n5888# 0.015026f
C200 drain_left.n182 a_n1220_n5888# 0.035516f
C201 drain_left.n183 a_n1220_n5888# 0.01591f
C202 drain_left.n184 a_n1220_n5888# 0.027963f
C203 drain_left.n185 a_n1220_n5888# 0.015026f
C204 drain_left.n186 a_n1220_n5888# 0.026637f
C205 drain_left.n187 a_n1220_n5888# 0.025107f
C206 drain_left.t5 a_n1220_n5888# 0.061942f
C207 drain_left.n188 a_n1220_n5888# 0.34117f
C208 drain_left.n189 a_n1220_n5888# 3.02755f
C209 drain_left.n190 a_n1220_n5888# 0.015026f
C210 drain_left.n191 a_n1220_n5888# 0.01591f
C211 drain_left.n192 a_n1220_n5888# 0.035516f
C212 drain_left.n193 a_n1220_n5888# 0.035516f
C213 drain_left.n194 a_n1220_n5888# 0.01591f
C214 drain_left.n195 a_n1220_n5888# 0.015026f
C215 drain_left.n196 a_n1220_n5888# 0.027963f
C216 drain_left.n197 a_n1220_n5888# 0.027963f
C217 drain_left.n198 a_n1220_n5888# 0.015026f
C218 drain_left.n199 a_n1220_n5888# 0.01591f
C219 drain_left.n200 a_n1220_n5888# 0.035516f
C220 drain_left.n201 a_n1220_n5888# 0.035516f
C221 drain_left.n202 a_n1220_n5888# 0.01591f
C222 drain_left.n203 a_n1220_n5888# 0.015026f
C223 drain_left.n204 a_n1220_n5888# 0.027963f
C224 drain_left.n205 a_n1220_n5888# 0.027963f
C225 drain_left.n206 a_n1220_n5888# 0.015026f
C226 drain_left.n207 a_n1220_n5888# 0.01591f
C227 drain_left.n208 a_n1220_n5888# 0.035516f
C228 drain_left.n209 a_n1220_n5888# 0.035516f
C229 drain_left.n210 a_n1220_n5888# 0.035516f
C230 drain_left.n211 a_n1220_n5888# 0.015468f
C231 drain_left.n212 a_n1220_n5888# 0.015026f
C232 drain_left.n213 a_n1220_n5888# 0.027963f
C233 drain_left.n214 a_n1220_n5888# 0.027963f
C234 drain_left.n215 a_n1220_n5888# 0.015026f
C235 drain_left.n216 a_n1220_n5888# 0.01591f
C236 drain_left.n217 a_n1220_n5888# 0.035516f
C237 drain_left.n218 a_n1220_n5888# 0.035516f
C238 drain_left.n219 a_n1220_n5888# 0.01591f
C239 drain_left.n220 a_n1220_n5888# 0.015026f
C240 drain_left.n221 a_n1220_n5888# 0.027963f
C241 drain_left.n222 a_n1220_n5888# 0.027963f
C242 drain_left.n223 a_n1220_n5888# 0.015026f
C243 drain_left.n224 a_n1220_n5888# 0.01591f
C244 drain_left.n225 a_n1220_n5888# 0.035516f
C245 drain_left.n226 a_n1220_n5888# 0.035516f
C246 drain_left.n227 a_n1220_n5888# 0.01591f
C247 drain_left.n228 a_n1220_n5888# 0.015026f
C248 drain_left.n229 a_n1220_n5888# 0.027963f
C249 drain_left.n230 a_n1220_n5888# 0.027963f
C250 drain_left.n231 a_n1220_n5888# 0.015026f
C251 drain_left.n232 a_n1220_n5888# 0.01591f
C252 drain_left.n233 a_n1220_n5888# 0.035516f
C253 drain_left.n234 a_n1220_n5888# 0.035516f
C254 drain_left.n235 a_n1220_n5888# 0.01591f
C255 drain_left.n236 a_n1220_n5888# 0.015026f
C256 drain_left.n237 a_n1220_n5888# 0.027963f
C257 drain_left.n238 a_n1220_n5888# 0.027963f
C258 drain_left.n239 a_n1220_n5888# 0.015026f
C259 drain_left.n240 a_n1220_n5888# 0.01591f
C260 drain_left.n241 a_n1220_n5888# 0.035516f
C261 drain_left.n242 a_n1220_n5888# 0.035516f
C262 drain_left.n243 a_n1220_n5888# 0.01591f
C263 drain_left.n244 a_n1220_n5888# 0.015026f
C264 drain_left.n245 a_n1220_n5888# 0.027963f
C265 drain_left.n246 a_n1220_n5888# 0.027963f
C266 drain_left.n247 a_n1220_n5888# 0.015026f
C267 drain_left.n248 a_n1220_n5888# 0.01591f
C268 drain_left.n249 a_n1220_n5888# 0.035516f
C269 drain_left.n250 a_n1220_n5888# 0.035516f
C270 drain_left.n251 a_n1220_n5888# 0.01591f
C271 drain_left.n252 a_n1220_n5888# 0.015026f
C272 drain_left.n253 a_n1220_n5888# 0.027963f
C273 drain_left.n254 a_n1220_n5888# 0.027963f
C274 drain_left.n255 a_n1220_n5888# 0.015026f
C275 drain_left.n256 a_n1220_n5888# 0.015468f
C276 drain_left.n257 a_n1220_n5888# 0.015468f
C277 drain_left.n258 a_n1220_n5888# 0.035516f
C278 drain_left.n259 a_n1220_n5888# 0.035516f
C279 drain_left.n260 a_n1220_n5888# 0.01591f
C280 drain_left.n261 a_n1220_n5888# 0.015026f
C281 drain_left.n262 a_n1220_n5888# 0.027963f
C282 drain_left.n263 a_n1220_n5888# 0.027963f
C283 drain_left.n264 a_n1220_n5888# 0.015026f
C284 drain_left.n265 a_n1220_n5888# 0.01591f
C285 drain_left.n266 a_n1220_n5888# 0.035516f
C286 drain_left.n267 a_n1220_n5888# 0.035516f
C287 drain_left.n268 a_n1220_n5888# 0.01591f
C288 drain_left.n269 a_n1220_n5888# 0.015026f
C289 drain_left.n270 a_n1220_n5888# 0.027963f
C290 drain_left.n271 a_n1220_n5888# 0.027963f
C291 drain_left.n272 a_n1220_n5888# 0.015026f
C292 drain_left.n273 a_n1220_n5888# 0.01591f
C293 drain_left.n274 a_n1220_n5888# 0.035516f
C294 drain_left.n275 a_n1220_n5888# 0.075552f
C295 drain_left.n276 a_n1220_n5888# 0.01591f
C296 drain_left.n277 a_n1220_n5888# 0.015026f
C297 drain_left.n278 a_n1220_n5888# 0.061579f
C298 drain_left.n279 a_n1220_n5888# 0.062521f
C299 drain_left.t4 a_n1220_n5888# 0.552427f
C300 drain_left.t2 a_n1220_n5888# 0.552427f
C301 drain_left.n280 a_n1220_n5888# 5.0912f
C302 drain_left.n281 a_n1220_n5888# 0.666884f
C303 plus.t0 a_n1220_n5888# 1.26226f
C304 plus.n0 a_n1220_n5888# 0.474269f
C305 plus.t1 a_n1220_n5888# 1.25044f
C306 plus.n1 a_n1220_n5888# 0.455009f
C307 plus.t3 a_n1220_n5888# 1.26226f
C308 plus.n2 a_n1220_n5888# 0.474176f
C309 plus.n3 a_n1220_n5888# 1.14172f
C310 plus.t4 a_n1220_n5888# 1.26226f
C311 plus.n4 a_n1220_n5888# 0.474269f
C312 plus.t5 a_n1220_n5888# 1.26226f
C313 plus.t2 a_n1220_n5888# 1.25044f
C314 plus.n5 a_n1220_n5888# 0.455009f
C315 plus.n6 a_n1220_n5888# 0.474176f
C316 plus.n7 a_n1220_n5888# 2.18183f
C317 drain_right.n0 a_n1220_n5888# 0.038444f
C318 drain_right.n1 a_n1220_n5888# 0.027886f
C319 drain_right.n2 a_n1220_n5888# 0.014985f
C320 drain_right.n3 a_n1220_n5888# 0.035418f
C321 drain_right.n4 a_n1220_n5888# 0.015866f
C322 drain_right.n5 a_n1220_n5888# 0.027886f
C323 drain_right.n6 a_n1220_n5888# 0.014985f
C324 drain_right.n7 a_n1220_n5888# 0.035418f
C325 drain_right.n8 a_n1220_n5888# 0.015866f
C326 drain_right.n9 a_n1220_n5888# 0.027886f
C327 drain_right.n10 a_n1220_n5888# 0.014985f
C328 drain_right.n11 a_n1220_n5888# 0.035418f
C329 drain_right.n12 a_n1220_n5888# 0.015866f
C330 drain_right.n13 a_n1220_n5888# 0.027886f
C331 drain_right.n14 a_n1220_n5888# 0.014985f
C332 drain_right.n15 a_n1220_n5888# 0.035418f
C333 drain_right.n16 a_n1220_n5888# 0.015866f
C334 drain_right.n17 a_n1220_n5888# 0.027886f
C335 drain_right.n18 a_n1220_n5888# 0.014985f
C336 drain_right.n19 a_n1220_n5888# 0.035418f
C337 drain_right.n20 a_n1220_n5888# 0.015866f
C338 drain_right.n21 a_n1220_n5888# 0.027886f
C339 drain_right.n22 a_n1220_n5888# 0.014985f
C340 drain_right.n23 a_n1220_n5888# 0.035418f
C341 drain_right.n24 a_n1220_n5888# 0.015866f
C342 drain_right.n25 a_n1220_n5888# 0.027886f
C343 drain_right.n26 a_n1220_n5888# 0.014985f
C344 drain_right.n27 a_n1220_n5888# 0.035418f
C345 drain_right.n28 a_n1220_n5888# 0.015866f
C346 drain_right.n29 a_n1220_n5888# 0.027886f
C347 drain_right.n30 a_n1220_n5888# 0.014985f
C348 drain_right.n31 a_n1220_n5888# 0.035418f
C349 drain_right.n32 a_n1220_n5888# 0.015866f
C350 drain_right.n33 a_n1220_n5888# 0.027886f
C351 drain_right.n34 a_n1220_n5888# 0.015426f
C352 drain_right.n35 a_n1220_n5888# 0.035418f
C353 drain_right.n36 a_n1220_n5888# 0.015866f
C354 drain_right.n37 a_n1220_n5888# 0.027886f
C355 drain_right.n38 a_n1220_n5888# 0.014985f
C356 drain_right.n39 a_n1220_n5888# 0.035418f
C357 drain_right.n40 a_n1220_n5888# 0.015866f
C358 drain_right.n41 a_n1220_n5888# 0.027886f
C359 drain_right.n42 a_n1220_n5888# 0.014985f
C360 drain_right.n43 a_n1220_n5888# 0.026564f
C361 drain_right.n44 a_n1220_n5888# 0.025038f
C362 drain_right.t3 a_n1220_n5888# 0.061772f
C363 drain_right.n45 a_n1220_n5888# 0.340233f
C364 drain_right.n46 a_n1220_n5888# 3.01923f
C365 drain_right.n47 a_n1220_n5888# 0.014985f
C366 drain_right.n48 a_n1220_n5888# 0.015866f
C367 drain_right.n49 a_n1220_n5888# 0.035418f
C368 drain_right.n50 a_n1220_n5888# 0.035418f
C369 drain_right.n51 a_n1220_n5888# 0.015866f
C370 drain_right.n52 a_n1220_n5888# 0.014985f
C371 drain_right.n53 a_n1220_n5888# 0.027886f
C372 drain_right.n54 a_n1220_n5888# 0.027886f
C373 drain_right.n55 a_n1220_n5888# 0.014985f
C374 drain_right.n56 a_n1220_n5888# 0.015866f
C375 drain_right.n57 a_n1220_n5888# 0.035418f
C376 drain_right.n58 a_n1220_n5888# 0.035418f
C377 drain_right.n59 a_n1220_n5888# 0.015866f
C378 drain_right.n60 a_n1220_n5888# 0.014985f
C379 drain_right.n61 a_n1220_n5888# 0.027886f
C380 drain_right.n62 a_n1220_n5888# 0.027886f
C381 drain_right.n63 a_n1220_n5888# 0.014985f
C382 drain_right.n64 a_n1220_n5888# 0.014985f
C383 drain_right.n65 a_n1220_n5888# 0.015866f
C384 drain_right.n66 a_n1220_n5888# 0.035418f
C385 drain_right.n67 a_n1220_n5888# 0.035418f
C386 drain_right.n68 a_n1220_n5888# 0.035418f
C387 drain_right.n69 a_n1220_n5888# 0.015426f
C388 drain_right.n70 a_n1220_n5888# 0.014985f
C389 drain_right.n71 a_n1220_n5888# 0.027886f
C390 drain_right.n72 a_n1220_n5888# 0.027886f
C391 drain_right.n73 a_n1220_n5888# 0.014985f
C392 drain_right.n74 a_n1220_n5888# 0.015866f
C393 drain_right.n75 a_n1220_n5888# 0.035418f
C394 drain_right.n76 a_n1220_n5888# 0.035418f
C395 drain_right.n77 a_n1220_n5888# 0.015866f
C396 drain_right.n78 a_n1220_n5888# 0.014985f
C397 drain_right.n79 a_n1220_n5888# 0.027886f
C398 drain_right.n80 a_n1220_n5888# 0.027886f
C399 drain_right.n81 a_n1220_n5888# 0.014985f
C400 drain_right.n82 a_n1220_n5888# 0.015866f
C401 drain_right.n83 a_n1220_n5888# 0.035418f
C402 drain_right.n84 a_n1220_n5888# 0.035418f
C403 drain_right.n85 a_n1220_n5888# 0.015866f
C404 drain_right.n86 a_n1220_n5888# 0.014985f
C405 drain_right.n87 a_n1220_n5888# 0.027886f
C406 drain_right.n88 a_n1220_n5888# 0.027886f
C407 drain_right.n89 a_n1220_n5888# 0.014985f
C408 drain_right.n90 a_n1220_n5888# 0.015866f
C409 drain_right.n91 a_n1220_n5888# 0.035418f
C410 drain_right.n92 a_n1220_n5888# 0.035418f
C411 drain_right.n93 a_n1220_n5888# 0.015866f
C412 drain_right.n94 a_n1220_n5888# 0.014985f
C413 drain_right.n95 a_n1220_n5888# 0.027886f
C414 drain_right.n96 a_n1220_n5888# 0.027886f
C415 drain_right.n97 a_n1220_n5888# 0.014985f
C416 drain_right.n98 a_n1220_n5888# 0.015866f
C417 drain_right.n99 a_n1220_n5888# 0.035418f
C418 drain_right.n100 a_n1220_n5888# 0.035418f
C419 drain_right.n101 a_n1220_n5888# 0.015866f
C420 drain_right.n102 a_n1220_n5888# 0.014985f
C421 drain_right.n103 a_n1220_n5888# 0.027886f
C422 drain_right.n104 a_n1220_n5888# 0.027886f
C423 drain_right.n105 a_n1220_n5888# 0.014985f
C424 drain_right.n106 a_n1220_n5888# 0.015866f
C425 drain_right.n107 a_n1220_n5888# 0.035418f
C426 drain_right.n108 a_n1220_n5888# 0.035418f
C427 drain_right.n109 a_n1220_n5888# 0.035418f
C428 drain_right.n110 a_n1220_n5888# 0.015866f
C429 drain_right.n111 a_n1220_n5888# 0.014985f
C430 drain_right.n112 a_n1220_n5888# 0.027886f
C431 drain_right.n113 a_n1220_n5888# 0.027886f
C432 drain_right.n114 a_n1220_n5888# 0.014985f
C433 drain_right.n115 a_n1220_n5888# 0.015426f
C434 drain_right.n116 a_n1220_n5888# 0.015426f
C435 drain_right.n117 a_n1220_n5888# 0.035418f
C436 drain_right.n118 a_n1220_n5888# 0.035418f
C437 drain_right.n119 a_n1220_n5888# 0.015866f
C438 drain_right.n120 a_n1220_n5888# 0.014985f
C439 drain_right.n121 a_n1220_n5888# 0.027886f
C440 drain_right.n122 a_n1220_n5888# 0.027886f
C441 drain_right.n123 a_n1220_n5888# 0.014985f
C442 drain_right.n124 a_n1220_n5888# 0.015866f
C443 drain_right.n125 a_n1220_n5888# 0.035418f
C444 drain_right.n126 a_n1220_n5888# 0.035418f
C445 drain_right.n127 a_n1220_n5888# 0.015866f
C446 drain_right.n128 a_n1220_n5888# 0.014985f
C447 drain_right.n129 a_n1220_n5888# 0.027886f
C448 drain_right.n130 a_n1220_n5888# 0.027886f
C449 drain_right.n131 a_n1220_n5888# 0.014985f
C450 drain_right.n132 a_n1220_n5888# 0.015866f
C451 drain_right.n133 a_n1220_n5888# 0.035418f
C452 drain_right.n134 a_n1220_n5888# 0.075344f
C453 drain_right.n135 a_n1220_n5888# 0.015866f
C454 drain_right.n136 a_n1220_n5888# 0.014985f
C455 drain_right.n137 a_n1220_n5888# 0.06141f
C456 drain_right.n138 a_n1220_n5888# 0.061836f
C457 drain_right.t1 a_n1220_n5888# 0.550909f
C458 drain_right.t4 a_n1220_n5888# 0.550909f
C459 drain_right.n139 a_n1220_n5888# 5.07765f
C460 drain_right.n140 a_n1220_n5888# 2.4332f
C461 drain_right.t0 a_n1220_n5888# 0.550909f
C462 drain_right.t2 a_n1220_n5888# 0.550909f
C463 drain_right.n141 a_n1220_n5888# 5.08037f
C464 drain_right.n142 a_n1220_n5888# 0.038444f
C465 drain_right.n143 a_n1220_n5888# 0.027886f
C466 drain_right.n144 a_n1220_n5888# 0.014985f
C467 drain_right.n145 a_n1220_n5888# 0.035418f
C468 drain_right.n146 a_n1220_n5888# 0.015866f
C469 drain_right.n147 a_n1220_n5888# 0.027886f
C470 drain_right.n148 a_n1220_n5888# 0.014985f
C471 drain_right.n149 a_n1220_n5888# 0.035418f
C472 drain_right.n150 a_n1220_n5888# 0.015866f
C473 drain_right.n151 a_n1220_n5888# 0.027886f
C474 drain_right.n152 a_n1220_n5888# 0.014985f
C475 drain_right.n153 a_n1220_n5888# 0.035418f
C476 drain_right.n154 a_n1220_n5888# 0.015866f
C477 drain_right.n155 a_n1220_n5888# 0.027886f
C478 drain_right.n156 a_n1220_n5888# 0.014985f
C479 drain_right.n157 a_n1220_n5888# 0.035418f
C480 drain_right.n158 a_n1220_n5888# 0.035418f
C481 drain_right.n159 a_n1220_n5888# 0.015866f
C482 drain_right.n160 a_n1220_n5888# 0.027886f
C483 drain_right.n161 a_n1220_n5888# 0.014985f
C484 drain_right.n162 a_n1220_n5888# 0.035418f
C485 drain_right.n163 a_n1220_n5888# 0.015866f
C486 drain_right.n164 a_n1220_n5888# 0.027886f
C487 drain_right.n165 a_n1220_n5888# 0.014985f
C488 drain_right.n166 a_n1220_n5888# 0.035418f
C489 drain_right.n167 a_n1220_n5888# 0.015866f
C490 drain_right.n168 a_n1220_n5888# 0.027886f
C491 drain_right.n169 a_n1220_n5888# 0.014985f
C492 drain_right.n170 a_n1220_n5888# 0.035418f
C493 drain_right.n171 a_n1220_n5888# 0.015866f
C494 drain_right.n172 a_n1220_n5888# 0.027886f
C495 drain_right.n173 a_n1220_n5888# 0.014985f
C496 drain_right.n174 a_n1220_n5888# 0.035418f
C497 drain_right.n175 a_n1220_n5888# 0.015866f
C498 drain_right.n176 a_n1220_n5888# 0.027886f
C499 drain_right.n177 a_n1220_n5888# 0.015426f
C500 drain_right.n178 a_n1220_n5888# 0.035418f
C501 drain_right.n179 a_n1220_n5888# 0.014985f
C502 drain_right.n180 a_n1220_n5888# 0.015866f
C503 drain_right.n181 a_n1220_n5888# 0.027886f
C504 drain_right.n182 a_n1220_n5888# 0.014985f
C505 drain_right.n183 a_n1220_n5888# 0.035418f
C506 drain_right.n184 a_n1220_n5888# 0.015866f
C507 drain_right.n185 a_n1220_n5888# 0.027886f
C508 drain_right.n186 a_n1220_n5888# 0.014985f
C509 drain_right.n187 a_n1220_n5888# 0.026564f
C510 drain_right.n188 a_n1220_n5888# 0.025038f
C511 drain_right.t5 a_n1220_n5888# 0.061772f
C512 drain_right.n189 a_n1220_n5888# 0.340233f
C513 drain_right.n190 a_n1220_n5888# 3.01923f
C514 drain_right.n191 a_n1220_n5888# 0.014985f
C515 drain_right.n192 a_n1220_n5888# 0.015866f
C516 drain_right.n193 a_n1220_n5888# 0.035418f
C517 drain_right.n194 a_n1220_n5888# 0.035418f
C518 drain_right.n195 a_n1220_n5888# 0.015866f
C519 drain_right.n196 a_n1220_n5888# 0.014985f
C520 drain_right.n197 a_n1220_n5888# 0.027886f
C521 drain_right.n198 a_n1220_n5888# 0.027886f
C522 drain_right.n199 a_n1220_n5888# 0.014985f
C523 drain_right.n200 a_n1220_n5888# 0.015866f
C524 drain_right.n201 a_n1220_n5888# 0.035418f
C525 drain_right.n202 a_n1220_n5888# 0.035418f
C526 drain_right.n203 a_n1220_n5888# 0.015866f
C527 drain_right.n204 a_n1220_n5888# 0.014985f
C528 drain_right.n205 a_n1220_n5888# 0.027886f
C529 drain_right.n206 a_n1220_n5888# 0.027886f
C530 drain_right.n207 a_n1220_n5888# 0.014985f
C531 drain_right.n208 a_n1220_n5888# 0.015866f
C532 drain_right.n209 a_n1220_n5888# 0.035418f
C533 drain_right.n210 a_n1220_n5888# 0.035418f
C534 drain_right.n211 a_n1220_n5888# 0.035418f
C535 drain_right.n212 a_n1220_n5888# 0.015426f
C536 drain_right.n213 a_n1220_n5888# 0.014985f
C537 drain_right.n214 a_n1220_n5888# 0.027886f
C538 drain_right.n215 a_n1220_n5888# 0.027886f
C539 drain_right.n216 a_n1220_n5888# 0.014985f
C540 drain_right.n217 a_n1220_n5888# 0.015866f
C541 drain_right.n218 a_n1220_n5888# 0.035418f
C542 drain_right.n219 a_n1220_n5888# 0.035418f
C543 drain_right.n220 a_n1220_n5888# 0.015866f
C544 drain_right.n221 a_n1220_n5888# 0.014985f
C545 drain_right.n222 a_n1220_n5888# 0.027886f
C546 drain_right.n223 a_n1220_n5888# 0.027886f
C547 drain_right.n224 a_n1220_n5888# 0.014985f
C548 drain_right.n225 a_n1220_n5888# 0.015866f
C549 drain_right.n226 a_n1220_n5888# 0.035418f
C550 drain_right.n227 a_n1220_n5888# 0.035418f
C551 drain_right.n228 a_n1220_n5888# 0.015866f
C552 drain_right.n229 a_n1220_n5888# 0.014985f
C553 drain_right.n230 a_n1220_n5888# 0.027886f
C554 drain_right.n231 a_n1220_n5888# 0.027886f
C555 drain_right.n232 a_n1220_n5888# 0.014985f
C556 drain_right.n233 a_n1220_n5888# 0.015866f
C557 drain_right.n234 a_n1220_n5888# 0.035418f
C558 drain_right.n235 a_n1220_n5888# 0.035418f
C559 drain_right.n236 a_n1220_n5888# 0.015866f
C560 drain_right.n237 a_n1220_n5888# 0.014985f
C561 drain_right.n238 a_n1220_n5888# 0.027886f
C562 drain_right.n239 a_n1220_n5888# 0.027886f
C563 drain_right.n240 a_n1220_n5888# 0.014985f
C564 drain_right.n241 a_n1220_n5888# 0.015866f
C565 drain_right.n242 a_n1220_n5888# 0.035418f
C566 drain_right.n243 a_n1220_n5888# 0.035418f
C567 drain_right.n244 a_n1220_n5888# 0.015866f
C568 drain_right.n245 a_n1220_n5888# 0.014985f
C569 drain_right.n246 a_n1220_n5888# 0.027886f
C570 drain_right.n247 a_n1220_n5888# 0.027886f
C571 drain_right.n248 a_n1220_n5888# 0.014985f
C572 drain_right.n249 a_n1220_n5888# 0.015866f
C573 drain_right.n250 a_n1220_n5888# 0.035418f
C574 drain_right.n251 a_n1220_n5888# 0.035418f
C575 drain_right.n252 a_n1220_n5888# 0.015866f
C576 drain_right.n253 a_n1220_n5888# 0.014985f
C577 drain_right.n254 a_n1220_n5888# 0.027886f
C578 drain_right.n255 a_n1220_n5888# 0.027886f
C579 drain_right.n256 a_n1220_n5888# 0.014985f
C580 drain_right.n257 a_n1220_n5888# 0.015426f
C581 drain_right.n258 a_n1220_n5888# 0.015426f
C582 drain_right.n259 a_n1220_n5888# 0.035418f
C583 drain_right.n260 a_n1220_n5888# 0.035418f
C584 drain_right.n261 a_n1220_n5888# 0.015866f
C585 drain_right.n262 a_n1220_n5888# 0.014985f
C586 drain_right.n263 a_n1220_n5888# 0.027886f
C587 drain_right.n264 a_n1220_n5888# 0.027886f
C588 drain_right.n265 a_n1220_n5888# 0.014985f
C589 drain_right.n266 a_n1220_n5888# 0.015866f
C590 drain_right.n267 a_n1220_n5888# 0.035418f
C591 drain_right.n268 a_n1220_n5888# 0.035418f
C592 drain_right.n269 a_n1220_n5888# 0.015866f
C593 drain_right.n270 a_n1220_n5888# 0.014985f
C594 drain_right.n271 a_n1220_n5888# 0.027886f
C595 drain_right.n272 a_n1220_n5888# 0.027886f
C596 drain_right.n273 a_n1220_n5888# 0.014985f
C597 drain_right.n274 a_n1220_n5888# 0.015866f
C598 drain_right.n275 a_n1220_n5888# 0.035418f
C599 drain_right.n276 a_n1220_n5888# 0.075344f
C600 drain_right.n277 a_n1220_n5888# 0.015866f
C601 drain_right.n278 a_n1220_n5888# 0.014985f
C602 drain_right.n279 a_n1220_n5888# 0.06141f
C603 drain_right.n280 a_n1220_n5888# 0.061206f
C604 drain_right.n281 a_n1220_n5888# 0.674796f
C605 source.n0 a_n1220_n5888# 0.038272f
C606 source.n1 a_n1220_n5888# 0.027762f
C607 source.n2 a_n1220_n5888# 0.014918f
C608 source.n3 a_n1220_n5888# 0.035261f
C609 source.n4 a_n1220_n5888# 0.015796f
C610 source.n5 a_n1220_n5888# 0.027762f
C611 source.n6 a_n1220_n5888# 0.014918f
C612 source.n7 a_n1220_n5888# 0.035261f
C613 source.n8 a_n1220_n5888# 0.015796f
C614 source.n9 a_n1220_n5888# 0.027762f
C615 source.n10 a_n1220_n5888# 0.014918f
C616 source.n11 a_n1220_n5888# 0.035261f
C617 source.n12 a_n1220_n5888# 0.015796f
C618 source.n13 a_n1220_n5888# 0.027762f
C619 source.n14 a_n1220_n5888# 0.014918f
C620 source.n15 a_n1220_n5888# 0.035261f
C621 source.n16 a_n1220_n5888# 0.035261f
C622 source.n17 a_n1220_n5888# 0.015796f
C623 source.n18 a_n1220_n5888# 0.027762f
C624 source.n19 a_n1220_n5888# 0.014918f
C625 source.n20 a_n1220_n5888# 0.035261f
C626 source.n21 a_n1220_n5888# 0.015796f
C627 source.n22 a_n1220_n5888# 0.027762f
C628 source.n23 a_n1220_n5888# 0.014918f
C629 source.n24 a_n1220_n5888# 0.035261f
C630 source.n25 a_n1220_n5888# 0.015796f
C631 source.n26 a_n1220_n5888# 0.027762f
C632 source.n27 a_n1220_n5888# 0.014918f
C633 source.n28 a_n1220_n5888# 0.035261f
C634 source.n29 a_n1220_n5888# 0.015796f
C635 source.n30 a_n1220_n5888# 0.027762f
C636 source.n31 a_n1220_n5888# 0.014918f
C637 source.n32 a_n1220_n5888# 0.035261f
C638 source.n33 a_n1220_n5888# 0.015796f
C639 source.n34 a_n1220_n5888# 0.027762f
C640 source.n35 a_n1220_n5888# 0.015357f
C641 source.n36 a_n1220_n5888# 0.035261f
C642 source.n37 a_n1220_n5888# 0.014918f
C643 source.n38 a_n1220_n5888# 0.015796f
C644 source.n39 a_n1220_n5888# 0.027762f
C645 source.n40 a_n1220_n5888# 0.014918f
C646 source.n41 a_n1220_n5888# 0.035261f
C647 source.n42 a_n1220_n5888# 0.015796f
C648 source.n43 a_n1220_n5888# 0.027762f
C649 source.n44 a_n1220_n5888# 0.014918f
C650 source.n45 a_n1220_n5888# 0.026445f
C651 source.n46 a_n1220_n5888# 0.024927f
C652 source.t4 a_n1220_n5888# 0.061497f
C653 source.n47 a_n1220_n5888# 0.338716f
C654 source.n48 a_n1220_n5888# 3.00578f
C655 source.n49 a_n1220_n5888# 0.014918f
C656 source.n50 a_n1220_n5888# 0.015796f
C657 source.n51 a_n1220_n5888# 0.035261f
C658 source.n52 a_n1220_n5888# 0.035261f
C659 source.n53 a_n1220_n5888# 0.015796f
C660 source.n54 a_n1220_n5888# 0.014918f
C661 source.n55 a_n1220_n5888# 0.027762f
C662 source.n56 a_n1220_n5888# 0.027762f
C663 source.n57 a_n1220_n5888# 0.014918f
C664 source.n58 a_n1220_n5888# 0.015796f
C665 source.n59 a_n1220_n5888# 0.035261f
C666 source.n60 a_n1220_n5888# 0.035261f
C667 source.n61 a_n1220_n5888# 0.015796f
C668 source.n62 a_n1220_n5888# 0.014918f
C669 source.n63 a_n1220_n5888# 0.027762f
C670 source.n64 a_n1220_n5888# 0.027762f
C671 source.n65 a_n1220_n5888# 0.014918f
C672 source.n66 a_n1220_n5888# 0.015796f
C673 source.n67 a_n1220_n5888# 0.035261f
C674 source.n68 a_n1220_n5888# 0.035261f
C675 source.n69 a_n1220_n5888# 0.035261f
C676 source.n70 a_n1220_n5888# 0.015357f
C677 source.n71 a_n1220_n5888# 0.014918f
C678 source.n72 a_n1220_n5888# 0.027762f
C679 source.n73 a_n1220_n5888# 0.027762f
C680 source.n74 a_n1220_n5888# 0.014918f
C681 source.n75 a_n1220_n5888# 0.015796f
C682 source.n76 a_n1220_n5888# 0.035261f
C683 source.n77 a_n1220_n5888# 0.035261f
C684 source.n78 a_n1220_n5888# 0.015796f
C685 source.n79 a_n1220_n5888# 0.014918f
C686 source.n80 a_n1220_n5888# 0.027762f
C687 source.n81 a_n1220_n5888# 0.027762f
C688 source.n82 a_n1220_n5888# 0.014918f
C689 source.n83 a_n1220_n5888# 0.015796f
C690 source.n84 a_n1220_n5888# 0.035261f
C691 source.n85 a_n1220_n5888# 0.035261f
C692 source.n86 a_n1220_n5888# 0.015796f
C693 source.n87 a_n1220_n5888# 0.014918f
C694 source.n88 a_n1220_n5888# 0.027762f
C695 source.n89 a_n1220_n5888# 0.027762f
C696 source.n90 a_n1220_n5888# 0.014918f
C697 source.n91 a_n1220_n5888# 0.015796f
C698 source.n92 a_n1220_n5888# 0.035261f
C699 source.n93 a_n1220_n5888# 0.035261f
C700 source.n94 a_n1220_n5888# 0.015796f
C701 source.n95 a_n1220_n5888# 0.014918f
C702 source.n96 a_n1220_n5888# 0.027762f
C703 source.n97 a_n1220_n5888# 0.027762f
C704 source.n98 a_n1220_n5888# 0.014918f
C705 source.n99 a_n1220_n5888# 0.015796f
C706 source.n100 a_n1220_n5888# 0.035261f
C707 source.n101 a_n1220_n5888# 0.035261f
C708 source.n102 a_n1220_n5888# 0.015796f
C709 source.n103 a_n1220_n5888# 0.014918f
C710 source.n104 a_n1220_n5888# 0.027762f
C711 source.n105 a_n1220_n5888# 0.027762f
C712 source.n106 a_n1220_n5888# 0.014918f
C713 source.n107 a_n1220_n5888# 0.015796f
C714 source.n108 a_n1220_n5888# 0.035261f
C715 source.n109 a_n1220_n5888# 0.035261f
C716 source.n110 a_n1220_n5888# 0.015796f
C717 source.n111 a_n1220_n5888# 0.014918f
C718 source.n112 a_n1220_n5888# 0.027762f
C719 source.n113 a_n1220_n5888# 0.027762f
C720 source.n114 a_n1220_n5888# 0.014918f
C721 source.n115 a_n1220_n5888# 0.015357f
C722 source.n116 a_n1220_n5888# 0.015357f
C723 source.n117 a_n1220_n5888# 0.035261f
C724 source.n118 a_n1220_n5888# 0.035261f
C725 source.n119 a_n1220_n5888# 0.015796f
C726 source.n120 a_n1220_n5888# 0.014918f
C727 source.n121 a_n1220_n5888# 0.027762f
C728 source.n122 a_n1220_n5888# 0.027762f
C729 source.n123 a_n1220_n5888# 0.014918f
C730 source.n124 a_n1220_n5888# 0.015796f
C731 source.n125 a_n1220_n5888# 0.035261f
C732 source.n126 a_n1220_n5888# 0.035261f
C733 source.n127 a_n1220_n5888# 0.015796f
C734 source.n128 a_n1220_n5888# 0.014918f
C735 source.n129 a_n1220_n5888# 0.027762f
C736 source.n130 a_n1220_n5888# 0.027762f
C737 source.n131 a_n1220_n5888# 0.014918f
C738 source.n132 a_n1220_n5888# 0.015796f
C739 source.n133 a_n1220_n5888# 0.035261f
C740 source.n134 a_n1220_n5888# 0.075008f
C741 source.n135 a_n1220_n5888# 0.015796f
C742 source.n136 a_n1220_n5888# 0.014918f
C743 source.n137 a_n1220_n5888# 0.061136f
C744 source.n138 a_n1220_n5888# 0.041738f
C745 source.n139 a_n1220_n5888# 2.18185f
C746 source.t3 a_n1220_n5888# 0.548454f
C747 source.t0 a_n1220_n5888# 0.548454f
C748 source.n140 a_n1220_n5888# 4.96358f
C749 source.n141 a_n1220_n5888# 0.402847f
C750 source.n142 a_n1220_n5888# 0.038272f
C751 source.n143 a_n1220_n5888# 0.027762f
C752 source.n144 a_n1220_n5888# 0.014918f
C753 source.n145 a_n1220_n5888# 0.035261f
C754 source.n146 a_n1220_n5888# 0.015796f
C755 source.n147 a_n1220_n5888# 0.027762f
C756 source.n148 a_n1220_n5888# 0.014918f
C757 source.n149 a_n1220_n5888# 0.035261f
C758 source.n150 a_n1220_n5888# 0.015796f
C759 source.n151 a_n1220_n5888# 0.027762f
C760 source.n152 a_n1220_n5888# 0.014918f
C761 source.n153 a_n1220_n5888# 0.035261f
C762 source.n154 a_n1220_n5888# 0.015796f
C763 source.n155 a_n1220_n5888# 0.027762f
C764 source.n156 a_n1220_n5888# 0.014918f
C765 source.n157 a_n1220_n5888# 0.035261f
C766 source.n158 a_n1220_n5888# 0.035261f
C767 source.n159 a_n1220_n5888# 0.015796f
C768 source.n160 a_n1220_n5888# 0.027762f
C769 source.n161 a_n1220_n5888# 0.014918f
C770 source.n162 a_n1220_n5888# 0.035261f
C771 source.n163 a_n1220_n5888# 0.015796f
C772 source.n164 a_n1220_n5888# 0.027762f
C773 source.n165 a_n1220_n5888# 0.014918f
C774 source.n166 a_n1220_n5888# 0.035261f
C775 source.n167 a_n1220_n5888# 0.015796f
C776 source.n168 a_n1220_n5888# 0.027762f
C777 source.n169 a_n1220_n5888# 0.014918f
C778 source.n170 a_n1220_n5888# 0.035261f
C779 source.n171 a_n1220_n5888# 0.015796f
C780 source.n172 a_n1220_n5888# 0.027762f
C781 source.n173 a_n1220_n5888# 0.014918f
C782 source.n174 a_n1220_n5888# 0.035261f
C783 source.n175 a_n1220_n5888# 0.015796f
C784 source.n176 a_n1220_n5888# 0.027762f
C785 source.n177 a_n1220_n5888# 0.015357f
C786 source.n178 a_n1220_n5888# 0.035261f
C787 source.n179 a_n1220_n5888# 0.014918f
C788 source.n180 a_n1220_n5888# 0.015796f
C789 source.n181 a_n1220_n5888# 0.027762f
C790 source.n182 a_n1220_n5888# 0.014918f
C791 source.n183 a_n1220_n5888# 0.035261f
C792 source.n184 a_n1220_n5888# 0.015796f
C793 source.n185 a_n1220_n5888# 0.027762f
C794 source.n186 a_n1220_n5888# 0.014918f
C795 source.n187 a_n1220_n5888# 0.026445f
C796 source.n188 a_n1220_n5888# 0.024927f
C797 source.t10 a_n1220_n5888# 0.061497f
C798 source.n189 a_n1220_n5888# 0.338716f
C799 source.n190 a_n1220_n5888# 3.00578f
C800 source.n191 a_n1220_n5888# 0.014918f
C801 source.n192 a_n1220_n5888# 0.015796f
C802 source.n193 a_n1220_n5888# 0.035261f
C803 source.n194 a_n1220_n5888# 0.035261f
C804 source.n195 a_n1220_n5888# 0.015796f
C805 source.n196 a_n1220_n5888# 0.014918f
C806 source.n197 a_n1220_n5888# 0.027762f
C807 source.n198 a_n1220_n5888# 0.027762f
C808 source.n199 a_n1220_n5888# 0.014918f
C809 source.n200 a_n1220_n5888# 0.015796f
C810 source.n201 a_n1220_n5888# 0.035261f
C811 source.n202 a_n1220_n5888# 0.035261f
C812 source.n203 a_n1220_n5888# 0.015796f
C813 source.n204 a_n1220_n5888# 0.014918f
C814 source.n205 a_n1220_n5888# 0.027762f
C815 source.n206 a_n1220_n5888# 0.027762f
C816 source.n207 a_n1220_n5888# 0.014918f
C817 source.n208 a_n1220_n5888# 0.015796f
C818 source.n209 a_n1220_n5888# 0.035261f
C819 source.n210 a_n1220_n5888# 0.035261f
C820 source.n211 a_n1220_n5888# 0.035261f
C821 source.n212 a_n1220_n5888# 0.015357f
C822 source.n213 a_n1220_n5888# 0.014918f
C823 source.n214 a_n1220_n5888# 0.027762f
C824 source.n215 a_n1220_n5888# 0.027762f
C825 source.n216 a_n1220_n5888# 0.014918f
C826 source.n217 a_n1220_n5888# 0.015796f
C827 source.n218 a_n1220_n5888# 0.035261f
C828 source.n219 a_n1220_n5888# 0.035261f
C829 source.n220 a_n1220_n5888# 0.015796f
C830 source.n221 a_n1220_n5888# 0.014918f
C831 source.n222 a_n1220_n5888# 0.027762f
C832 source.n223 a_n1220_n5888# 0.027762f
C833 source.n224 a_n1220_n5888# 0.014918f
C834 source.n225 a_n1220_n5888# 0.015796f
C835 source.n226 a_n1220_n5888# 0.035261f
C836 source.n227 a_n1220_n5888# 0.035261f
C837 source.n228 a_n1220_n5888# 0.015796f
C838 source.n229 a_n1220_n5888# 0.014918f
C839 source.n230 a_n1220_n5888# 0.027762f
C840 source.n231 a_n1220_n5888# 0.027762f
C841 source.n232 a_n1220_n5888# 0.014918f
C842 source.n233 a_n1220_n5888# 0.015796f
C843 source.n234 a_n1220_n5888# 0.035261f
C844 source.n235 a_n1220_n5888# 0.035261f
C845 source.n236 a_n1220_n5888# 0.015796f
C846 source.n237 a_n1220_n5888# 0.014918f
C847 source.n238 a_n1220_n5888# 0.027762f
C848 source.n239 a_n1220_n5888# 0.027762f
C849 source.n240 a_n1220_n5888# 0.014918f
C850 source.n241 a_n1220_n5888# 0.015796f
C851 source.n242 a_n1220_n5888# 0.035261f
C852 source.n243 a_n1220_n5888# 0.035261f
C853 source.n244 a_n1220_n5888# 0.015796f
C854 source.n245 a_n1220_n5888# 0.014918f
C855 source.n246 a_n1220_n5888# 0.027762f
C856 source.n247 a_n1220_n5888# 0.027762f
C857 source.n248 a_n1220_n5888# 0.014918f
C858 source.n249 a_n1220_n5888# 0.015796f
C859 source.n250 a_n1220_n5888# 0.035261f
C860 source.n251 a_n1220_n5888# 0.035261f
C861 source.n252 a_n1220_n5888# 0.015796f
C862 source.n253 a_n1220_n5888# 0.014918f
C863 source.n254 a_n1220_n5888# 0.027762f
C864 source.n255 a_n1220_n5888# 0.027762f
C865 source.n256 a_n1220_n5888# 0.014918f
C866 source.n257 a_n1220_n5888# 0.015357f
C867 source.n258 a_n1220_n5888# 0.015357f
C868 source.n259 a_n1220_n5888# 0.035261f
C869 source.n260 a_n1220_n5888# 0.035261f
C870 source.n261 a_n1220_n5888# 0.015796f
C871 source.n262 a_n1220_n5888# 0.014918f
C872 source.n263 a_n1220_n5888# 0.027762f
C873 source.n264 a_n1220_n5888# 0.027762f
C874 source.n265 a_n1220_n5888# 0.014918f
C875 source.n266 a_n1220_n5888# 0.015796f
C876 source.n267 a_n1220_n5888# 0.035261f
C877 source.n268 a_n1220_n5888# 0.035261f
C878 source.n269 a_n1220_n5888# 0.015796f
C879 source.n270 a_n1220_n5888# 0.014918f
C880 source.n271 a_n1220_n5888# 0.027762f
C881 source.n272 a_n1220_n5888# 0.027762f
C882 source.n273 a_n1220_n5888# 0.014918f
C883 source.n274 a_n1220_n5888# 0.015796f
C884 source.n275 a_n1220_n5888# 0.035261f
C885 source.n276 a_n1220_n5888# 0.075008f
C886 source.n277 a_n1220_n5888# 0.015796f
C887 source.n278 a_n1220_n5888# 0.014918f
C888 source.n279 a_n1220_n5888# 0.061136f
C889 source.n280 a_n1220_n5888# 0.041738f
C890 source.n281 a_n1220_n5888# 0.136903f
C891 source.t8 a_n1220_n5888# 0.548454f
C892 source.t9 a_n1220_n5888# 0.548454f
C893 source.n282 a_n1220_n5888# 4.96358f
C894 source.n283 a_n1220_n5888# 3.00996f
C895 source.t2 a_n1220_n5888# 0.548454f
C896 source.t11 a_n1220_n5888# 0.548454f
C897 source.n284 a_n1220_n5888# 4.96358f
C898 source.n285 a_n1220_n5888# 3.00997f
C899 source.n286 a_n1220_n5888# 0.038272f
C900 source.n287 a_n1220_n5888# 0.027762f
C901 source.n288 a_n1220_n5888# 0.014918f
C902 source.n289 a_n1220_n5888# 0.035261f
C903 source.n290 a_n1220_n5888# 0.015796f
C904 source.n291 a_n1220_n5888# 0.027762f
C905 source.n292 a_n1220_n5888# 0.014918f
C906 source.n293 a_n1220_n5888# 0.035261f
C907 source.n294 a_n1220_n5888# 0.015796f
C908 source.n295 a_n1220_n5888# 0.027762f
C909 source.n296 a_n1220_n5888# 0.014918f
C910 source.n297 a_n1220_n5888# 0.035261f
C911 source.n298 a_n1220_n5888# 0.015796f
C912 source.n299 a_n1220_n5888# 0.027762f
C913 source.n300 a_n1220_n5888# 0.014918f
C914 source.n301 a_n1220_n5888# 0.035261f
C915 source.n302 a_n1220_n5888# 0.015796f
C916 source.n303 a_n1220_n5888# 0.027762f
C917 source.n304 a_n1220_n5888# 0.014918f
C918 source.n305 a_n1220_n5888# 0.035261f
C919 source.n306 a_n1220_n5888# 0.015796f
C920 source.n307 a_n1220_n5888# 0.027762f
C921 source.n308 a_n1220_n5888# 0.014918f
C922 source.n309 a_n1220_n5888# 0.035261f
C923 source.n310 a_n1220_n5888# 0.015796f
C924 source.n311 a_n1220_n5888# 0.027762f
C925 source.n312 a_n1220_n5888# 0.014918f
C926 source.n313 a_n1220_n5888# 0.035261f
C927 source.n314 a_n1220_n5888# 0.015796f
C928 source.n315 a_n1220_n5888# 0.027762f
C929 source.n316 a_n1220_n5888# 0.014918f
C930 source.n317 a_n1220_n5888# 0.035261f
C931 source.n318 a_n1220_n5888# 0.015796f
C932 source.n319 a_n1220_n5888# 0.027762f
C933 source.n320 a_n1220_n5888# 0.015357f
C934 source.n321 a_n1220_n5888# 0.035261f
C935 source.n322 a_n1220_n5888# 0.015796f
C936 source.n323 a_n1220_n5888# 0.027762f
C937 source.n324 a_n1220_n5888# 0.014918f
C938 source.n325 a_n1220_n5888# 0.035261f
C939 source.n326 a_n1220_n5888# 0.015796f
C940 source.n327 a_n1220_n5888# 0.027762f
C941 source.n328 a_n1220_n5888# 0.014918f
C942 source.n329 a_n1220_n5888# 0.026445f
C943 source.n330 a_n1220_n5888# 0.024927f
C944 source.t1 a_n1220_n5888# 0.061497f
C945 source.n331 a_n1220_n5888# 0.338716f
C946 source.n332 a_n1220_n5888# 3.00578f
C947 source.n333 a_n1220_n5888# 0.014918f
C948 source.n334 a_n1220_n5888# 0.015796f
C949 source.n335 a_n1220_n5888# 0.035261f
C950 source.n336 a_n1220_n5888# 0.035261f
C951 source.n337 a_n1220_n5888# 0.015796f
C952 source.n338 a_n1220_n5888# 0.014918f
C953 source.n339 a_n1220_n5888# 0.027762f
C954 source.n340 a_n1220_n5888# 0.027762f
C955 source.n341 a_n1220_n5888# 0.014918f
C956 source.n342 a_n1220_n5888# 0.015796f
C957 source.n343 a_n1220_n5888# 0.035261f
C958 source.n344 a_n1220_n5888# 0.035261f
C959 source.n345 a_n1220_n5888# 0.015796f
C960 source.n346 a_n1220_n5888# 0.014918f
C961 source.n347 a_n1220_n5888# 0.027762f
C962 source.n348 a_n1220_n5888# 0.027762f
C963 source.n349 a_n1220_n5888# 0.014918f
C964 source.n350 a_n1220_n5888# 0.014918f
C965 source.n351 a_n1220_n5888# 0.015796f
C966 source.n352 a_n1220_n5888# 0.035261f
C967 source.n353 a_n1220_n5888# 0.035261f
C968 source.n354 a_n1220_n5888# 0.035261f
C969 source.n355 a_n1220_n5888# 0.015357f
C970 source.n356 a_n1220_n5888# 0.014918f
C971 source.n357 a_n1220_n5888# 0.027762f
C972 source.n358 a_n1220_n5888# 0.027762f
C973 source.n359 a_n1220_n5888# 0.014918f
C974 source.n360 a_n1220_n5888# 0.015796f
C975 source.n361 a_n1220_n5888# 0.035261f
C976 source.n362 a_n1220_n5888# 0.035261f
C977 source.n363 a_n1220_n5888# 0.015796f
C978 source.n364 a_n1220_n5888# 0.014918f
C979 source.n365 a_n1220_n5888# 0.027762f
C980 source.n366 a_n1220_n5888# 0.027762f
C981 source.n367 a_n1220_n5888# 0.014918f
C982 source.n368 a_n1220_n5888# 0.015796f
C983 source.n369 a_n1220_n5888# 0.035261f
C984 source.n370 a_n1220_n5888# 0.035261f
C985 source.n371 a_n1220_n5888# 0.015796f
C986 source.n372 a_n1220_n5888# 0.014918f
C987 source.n373 a_n1220_n5888# 0.027762f
C988 source.n374 a_n1220_n5888# 0.027762f
C989 source.n375 a_n1220_n5888# 0.014918f
C990 source.n376 a_n1220_n5888# 0.015796f
C991 source.n377 a_n1220_n5888# 0.035261f
C992 source.n378 a_n1220_n5888# 0.035261f
C993 source.n379 a_n1220_n5888# 0.015796f
C994 source.n380 a_n1220_n5888# 0.014918f
C995 source.n381 a_n1220_n5888# 0.027762f
C996 source.n382 a_n1220_n5888# 0.027762f
C997 source.n383 a_n1220_n5888# 0.014918f
C998 source.n384 a_n1220_n5888# 0.015796f
C999 source.n385 a_n1220_n5888# 0.035261f
C1000 source.n386 a_n1220_n5888# 0.035261f
C1001 source.n387 a_n1220_n5888# 0.015796f
C1002 source.n388 a_n1220_n5888# 0.014918f
C1003 source.n389 a_n1220_n5888# 0.027762f
C1004 source.n390 a_n1220_n5888# 0.027762f
C1005 source.n391 a_n1220_n5888# 0.014918f
C1006 source.n392 a_n1220_n5888# 0.015796f
C1007 source.n393 a_n1220_n5888# 0.035261f
C1008 source.n394 a_n1220_n5888# 0.035261f
C1009 source.n395 a_n1220_n5888# 0.035261f
C1010 source.n396 a_n1220_n5888# 0.015796f
C1011 source.n397 a_n1220_n5888# 0.014918f
C1012 source.n398 a_n1220_n5888# 0.027762f
C1013 source.n399 a_n1220_n5888# 0.027762f
C1014 source.n400 a_n1220_n5888# 0.014918f
C1015 source.n401 a_n1220_n5888# 0.015357f
C1016 source.n402 a_n1220_n5888# 0.015357f
C1017 source.n403 a_n1220_n5888# 0.035261f
C1018 source.n404 a_n1220_n5888# 0.035261f
C1019 source.n405 a_n1220_n5888# 0.015796f
C1020 source.n406 a_n1220_n5888# 0.014918f
C1021 source.n407 a_n1220_n5888# 0.027762f
C1022 source.n408 a_n1220_n5888# 0.027762f
C1023 source.n409 a_n1220_n5888# 0.014918f
C1024 source.n410 a_n1220_n5888# 0.015796f
C1025 source.n411 a_n1220_n5888# 0.035261f
C1026 source.n412 a_n1220_n5888# 0.035261f
C1027 source.n413 a_n1220_n5888# 0.015796f
C1028 source.n414 a_n1220_n5888# 0.014918f
C1029 source.n415 a_n1220_n5888# 0.027762f
C1030 source.n416 a_n1220_n5888# 0.027762f
C1031 source.n417 a_n1220_n5888# 0.014918f
C1032 source.n418 a_n1220_n5888# 0.015796f
C1033 source.n419 a_n1220_n5888# 0.035261f
C1034 source.n420 a_n1220_n5888# 0.075008f
C1035 source.n421 a_n1220_n5888# 0.015796f
C1036 source.n422 a_n1220_n5888# 0.014918f
C1037 source.n423 a_n1220_n5888# 0.061136f
C1038 source.n424 a_n1220_n5888# 0.041738f
C1039 source.n425 a_n1220_n5888# 0.136903f
C1040 source.t6 a_n1220_n5888# 0.548454f
C1041 source.t5 a_n1220_n5888# 0.548454f
C1042 source.n426 a_n1220_n5888# 4.96358f
C1043 source.n427 a_n1220_n5888# 0.402849f
C1044 source.n428 a_n1220_n5888# 0.038272f
C1045 source.n429 a_n1220_n5888# 0.027762f
C1046 source.n430 a_n1220_n5888# 0.014918f
C1047 source.n431 a_n1220_n5888# 0.035261f
C1048 source.n432 a_n1220_n5888# 0.015796f
C1049 source.n433 a_n1220_n5888# 0.027762f
C1050 source.n434 a_n1220_n5888# 0.014918f
C1051 source.n435 a_n1220_n5888# 0.035261f
C1052 source.n436 a_n1220_n5888# 0.015796f
C1053 source.n437 a_n1220_n5888# 0.027762f
C1054 source.n438 a_n1220_n5888# 0.014918f
C1055 source.n439 a_n1220_n5888# 0.035261f
C1056 source.n440 a_n1220_n5888# 0.015796f
C1057 source.n441 a_n1220_n5888# 0.027762f
C1058 source.n442 a_n1220_n5888# 0.014918f
C1059 source.n443 a_n1220_n5888# 0.035261f
C1060 source.n444 a_n1220_n5888# 0.015796f
C1061 source.n445 a_n1220_n5888# 0.027762f
C1062 source.n446 a_n1220_n5888# 0.014918f
C1063 source.n447 a_n1220_n5888# 0.035261f
C1064 source.n448 a_n1220_n5888# 0.015796f
C1065 source.n449 a_n1220_n5888# 0.027762f
C1066 source.n450 a_n1220_n5888# 0.014918f
C1067 source.n451 a_n1220_n5888# 0.035261f
C1068 source.n452 a_n1220_n5888# 0.015796f
C1069 source.n453 a_n1220_n5888# 0.027762f
C1070 source.n454 a_n1220_n5888# 0.014918f
C1071 source.n455 a_n1220_n5888# 0.035261f
C1072 source.n456 a_n1220_n5888# 0.015796f
C1073 source.n457 a_n1220_n5888# 0.027762f
C1074 source.n458 a_n1220_n5888# 0.014918f
C1075 source.n459 a_n1220_n5888# 0.035261f
C1076 source.n460 a_n1220_n5888# 0.015796f
C1077 source.n461 a_n1220_n5888# 0.027762f
C1078 source.n462 a_n1220_n5888# 0.015357f
C1079 source.n463 a_n1220_n5888# 0.035261f
C1080 source.n464 a_n1220_n5888# 0.015796f
C1081 source.n465 a_n1220_n5888# 0.027762f
C1082 source.n466 a_n1220_n5888# 0.014918f
C1083 source.n467 a_n1220_n5888# 0.035261f
C1084 source.n468 a_n1220_n5888# 0.015796f
C1085 source.n469 a_n1220_n5888# 0.027762f
C1086 source.n470 a_n1220_n5888# 0.014918f
C1087 source.n471 a_n1220_n5888# 0.026445f
C1088 source.n472 a_n1220_n5888# 0.024927f
C1089 source.t7 a_n1220_n5888# 0.061497f
C1090 source.n473 a_n1220_n5888# 0.338716f
C1091 source.n474 a_n1220_n5888# 3.00578f
C1092 source.n475 a_n1220_n5888# 0.014918f
C1093 source.n476 a_n1220_n5888# 0.015796f
C1094 source.n477 a_n1220_n5888# 0.035261f
C1095 source.n478 a_n1220_n5888# 0.035261f
C1096 source.n479 a_n1220_n5888# 0.015796f
C1097 source.n480 a_n1220_n5888# 0.014918f
C1098 source.n481 a_n1220_n5888# 0.027762f
C1099 source.n482 a_n1220_n5888# 0.027762f
C1100 source.n483 a_n1220_n5888# 0.014918f
C1101 source.n484 a_n1220_n5888# 0.015796f
C1102 source.n485 a_n1220_n5888# 0.035261f
C1103 source.n486 a_n1220_n5888# 0.035261f
C1104 source.n487 a_n1220_n5888# 0.015796f
C1105 source.n488 a_n1220_n5888# 0.014918f
C1106 source.n489 a_n1220_n5888# 0.027762f
C1107 source.n490 a_n1220_n5888# 0.027762f
C1108 source.n491 a_n1220_n5888# 0.014918f
C1109 source.n492 a_n1220_n5888# 0.014918f
C1110 source.n493 a_n1220_n5888# 0.015796f
C1111 source.n494 a_n1220_n5888# 0.035261f
C1112 source.n495 a_n1220_n5888# 0.035261f
C1113 source.n496 a_n1220_n5888# 0.035261f
C1114 source.n497 a_n1220_n5888# 0.015357f
C1115 source.n498 a_n1220_n5888# 0.014918f
C1116 source.n499 a_n1220_n5888# 0.027762f
C1117 source.n500 a_n1220_n5888# 0.027762f
C1118 source.n501 a_n1220_n5888# 0.014918f
C1119 source.n502 a_n1220_n5888# 0.015796f
C1120 source.n503 a_n1220_n5888# 0.035261f
C1121 source.n504 a_n1220_n5888# 0.035261f
C1122 source.n505 a_n1220_n5888# 0.015796f
C1123 source.n506 a_n1220_n5888# 0.014918f
C1124 source.n507 a_n1220_n5888# 0.027762f
C1125 source.n508 a_n1220_n5888# 0.027762f
C1126 source.n509 a_n1220_n5888# 0.014918f
C1127 source.n510 a_n1220_n5888# 0.015796f
C1128 source.n511 a_n1220_n5888# 0.035261f
C1129 source.n512 a_n1220_n5888# 0.035261f
C1130 source.n513 a_n1220_n5888# 0.015796f
C1131 source.n514 a_n1220_n5888# 0.014918f
C1132 source.n515 a_n1220_n5888# 0.027762f
C1133 source.n516 a_n1220_n5888# 0.027762f
C1134 source.n517 a_n1220_n5888# 0.014918f
C1135 source.n518 a_n1220_n5888# 0.015796f
C1136 source.n519 a_n1220_n5888# 0.035261f
C1137 source.n520 a_n1220_n5888# 0.035261f
C1138 source.n521 a_n1220_n5888# 0.015796f
C1139 source.n522 a_n1220_n5888# 0.014918f
C1140 source.n523 a_n1220_n5888# 0.027762f
C1141 source.n524 a_n1220_n5888# 0.027762f
C1142 source.n525 a_n1220_n5888# 0.014918f
C1143 source.n526 a_n1220_n5888# 0.015796f
C1144 source.n527 a_n1220_n5888# 0.035261f
C1145 source.n528 a_n1220_n5888# 0.035261f
C1146 source.n529 a_n1220_n5888# 0.015796f
C1147 source.n530 a_n1220_n5888# 0.014918f
C1148 source.n531 a_n1220_n5888# 0.027762f
C1149 source.n532 a_n1220_n5888# 0.027762f
C1150 source.n533 a_n1220_n5888# 0.014918f
C1151 source.n534 a_n1220_n5888# 0.015796f
C1152 source.n535 a_n1220_n5888# 0.035261f
C1153 source.n536 a_n1220_n5888# 0.035261f
C1154 source.n537 a_n1220_n5888# 0.035261f
C1155 source.n538 a_n1220_n5888# 0.015796f
C1156 source.n539 a_n1220_n5888# 0.014918f
C1157 source.n540 a_n1220_n5888# 0.027762f
C1158 source.n541 a_n1220_n5888# 0.027762f
C1159 source.n542 a_n1220_n5888# 0.014918f
C1160 source.n543 a_n1220_n5888# 0.015357f
C1161 source.n544 a_n1220_n5888# 0.015357f
C1162 source.n545 a_n1220_n5888# 0.035261f
C1163 source.n546 a_n1220_n5888# 0.035261f
C1164 source.n547 a_n1220_n5888# 0.015796f
C1165 source.n548 a_n1220_n5888# 0.014918f
C1166 source.n549 a_n1220_n5888# 0.027762f
C1167 source.n550 a_n1220_n5888# 0.027762f
C1168 source.n551 a_n1220_n5888# 0.014918f
C1169 source.n552 a_n1220_n5888# 0.015796f
C1170 source.n553 a_n1220_n5888# 0.035261f
C1171 source.n554 a_n1220_n5888# 0.035261f
C1172 source.n555 a_n1220_n5888# 0.015796f
C1173 source.n556 a_n1220_n5888# 0.014918f
C1174 source.n557 a_n1220_n5888# 0.027762f
C1175 source.n558 a_n1220_n5888# 0.027762f
C1176 source.n559 a_n1220_n5888# 0.014918f
C1177 source.n560 a_n1220_n5888# 0.015796f
C1178 source.n561 a_n1220_n5888# 0.035261f
C1179 source.n562 a_n1220_n5888# 0.075008f
C1180 source.n563 a_n1220_n5888# 0.015796f
C1181 source.n564 a_n1220_n5888# 0.014918f
C1182 source.n565 a_n1220_n5888# 0.061136f
C1183 source.n566 a_n1220_n5888# 0.041738f
C1184 source.n567 a_n1220_n5888# 0.269326f
C1185 source.n568 a_n1220_n5888# 2.95944f
C1186 minus.t3 a_n1220_n5888# 1.24596f
C1187 minus.n0 a_n1220_n5888# 0.468143f
C1188 minus.t0 a_n1220_n5888# 1.24596f
C1189 minus.t5 a_n1220_n5888# 1.23429f
C1190 minus.n1 a_n1220_n5888# 0.449132f
C1191 minus.n2 a_n1220_n5888# 0.468051f
C1192 minus.n3 a_n1220_n5888# 2.81785f
C1193 minus.t2 a_n1220_n5888# 1.24596f
C1194 minus.n4 a_n1220_n5888# 0.468143f
C1195 minus.t4 a_n1220_n5888# 1.23429f
C1196 minus.n5 a_n1220_n5888# 0.449132f
C1197 minus.t1 a_n1220_n5888# 1.24596f
C1198 minus.n6 a_n1220_n5888# 0.468051f
C1199 minus.n7 a_n1220_n5888# 0.465484f
C1200 minus.n8 a_n1220_n5888# 3.25519f
.ends

