* NGSPICE file created from diffpair480.ext - technology: sky130A

.subckt diffpair480 minus drain_right drain_left source plus
X0 drain_right minus source a_n976_n3892# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=7.125 ps=30.95 w=15 l=0.15
X1 a_n976_n3892# a_n976_n3892# a_n976_n3892# a_n976_n3892# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=57 ps=247.6 w=15 l=0.15
X2 drain_left plus source a_n976_n3892# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=7.125 ps=30.95 w=15 l=0.15
X3 drain_left plus source a_n976_n3892# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=7.125 ps=30.95 w=15 l=0.15
X4 a_n976_n3892# a_n976_n3892# a_n976_n3892# a_n976_n3892# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X5 drain_right minus source a_n976_n3892# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=7.125 ps=30.95 w=15 l=0.15
X6 a_n976_n3892# a_n976_n3892# a_n976_n3892# a_n976_n3892# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
X7 a_n976_n3892# a_n976_n3892# a_n976_n3892# a_n976_n3892# sky130_fd_pr__nfet_01v8 ad=7.125 pd=30.95 as=0 ps=0 w=15 l=0.15
.ends

