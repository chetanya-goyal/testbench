* NGSPICE file created from diffpair438.ext - technology: sky130A

.subckt diffpair438 minus drain_right drain_left source plus
X0 source.t37 minus.t0 drain_right.t10 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X1 source.t36 minus.t1 drain_right.t11 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X2 drain_left.t19 plus.t0 source.t8 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X3 source.t35 minus.t2 drain_right.t9 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X4 drain_right.t13 minus.t3 source.t34 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X5 drain_right.t12 minus.t4 source.t33 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X6 drain_right.t19 minus.t5 source.t32 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X7 drain_left.t18 plus.t1 source.t1 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X8 drain_left.t17 plus.t2 source.t4 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X9 source.t11 plus.t3 drain_left.t16 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X10 drain_left.t15 plus.t4 source.t13 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X11 drain_right.t16 minus.t6 source.t31 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X12 source.t30 minus.t7 drain_right.t3 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X13 a_n2102_n3288# a_n2102_n3288# a_n2102_n3288# a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=37.44 ps=198.24 w=12 l=0.3
X14 source.t29 minus.t8 drain_right.t15 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X15 source.t28 minus.t9 drain_right.t14 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X16 a_n2102_n3288# a_n2102_n3288# a_n2102_n3288# a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.3
X17 source.t14 plus.t5 drain_left.t14 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X18 source.t9 plus.t6 drain_left.t13 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X19 drain_left.t12 plus.t7 source.t38 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X20 source.t27 minus.t10 drain_right.t5 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X21 source.t39 plus.t8 drain_left.t11 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X22 source.t3 plus.t9 drain_left.t10 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X23 a_n2102_n3288# a_n2102_n3288# a_n2102_n3288# a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.3
X24 source.t0 plus.t10 drain_left.t9 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X25 drain_right.t18 minus.t11 source.t26 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X26 a_n2102_n3288# a_n2102_n3288# a_n2102_n3288# a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=0.3
X27 drain_left.t8 plus.t11 source.t2 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X28 drain_right.t8 minus.t12 source.t25 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X29 drain_right.t4 minus.t13 source.t24 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X30 source.t23 minus.t14 drain_right.t1 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X31 source.t16 plus.t12 drain_left.t7 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X32 drain_right.t2 minus.t15 source.t22 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X33 source.t10 plus.t13 drain_left.t6 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X34 drain_right.t7 minus.t16 source.t21 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X35 source.t6 plus.t14 drain_left.t5 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=0.3
X36 drain_left.t4 plus.t15 source.t12 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X37 drain_right.t0 minus.t17 source.t20 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X38 drain_left.t3 plus.t16 source.t15 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=0.3
X39 drain_left.t2 plus.t17 source.t5 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X40 source.t19 minus.t18 drain_right.t17 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X41 source.t18 minus.t19 drain_right.t6 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X42 source.t7 plus.t18 drain_left.t1 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
X43 drain_left.t0 plus.t19 source.t17 a_n2102_n3288# sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=0.3
R0 minus.n27 minus.t7 1117.36
R1 minus.n7 minus.t11 1117.36
R2 minus.n56 minus.t3 1117.36
R3 minus.n35 minus.t1 1117.36
R4 minus.n26 minus.t5 1068.43
R5 minus.n24 minus.t19 1068.43
R6 minus.n3 minus.t6 1068.43
R7 minus.n18 minus.t2 1068.43
R8 minus.n16 minus.t17 1068.43
R9 minus.n4 minus.t10 1068.43
R10 minus.n10 minus.t4 1068.43
R11 minus.n6 minus.t18 1068.43
R12 minus.n55 minus.t14 1068.43
R13 minus.n53 minus.t15 1068.43
R14 minus.n47 minus.t8 1068.43
R15 minus.n46 minus.t16 1068.43
R16 minus.n44 minus.t9 1068.43
R17 minus.n32 minus.t12 1068.43
R18 minus.n38 minus.t0 1068.43
R19 minus.n34 minus.t13 1068.43
R20 minus.n8 minus.n7 161.489
R21 minus.n36 minus.n35 161.489
R22 minus.n28 minus.n27 161.3
R23 minus.n25 minus.n0 161.3
R24 minus.n23 minus.n22 161.3
R25 minus.n21 minus.n1 161.3
R26 minus.n20 minus.n19 161.3
R27 minus.n17 minus.n2 161.3
R28 minus.n15 minus.n14 161.3
R29 minus.n13 minus.n12 161.3
R30 minus.n11 minus.n5 161.3
R31 minus.n9 minus.n8 161.3
R32 minus.n57 minus.n56 161.3
R33 minus.n54 minus.n29 161.3
R34 minus.n52 minus.n51 161.3
R35 minus.n50 minus.n30 161.3
R36 minus.n49 minus.n48 161.3
R37 minus.n45 minus.n31 161.3
R38 minus.n43 minus.n42 161.3
R39 minus.n41 minus.n40 161.3
R40 minus.n39 minus.n33 161.3
R41 minus.n37 minus.n36 161.3
R42 minus.n23 minus.n1 73.0308
R43 minus.n12 minus.n11 73.0308
R44 minus.n40 minus.n39 73.0308
R45 minus.n52 minus.n30 73.0308
R46 minus.n19 minus.n3 64.9975
R47 minus.n15 minus.n4 64.9975
R48 minus.n43 minus.n32 64.9975
R49 minus.n48 minus.n47 64.9975
R50 minus.n25 minus.n24 62.0763
R51 minus.n10 minus.n9 62.0763
R52 minus.n38 minus.n37 62.0763
R53 minus.n54 minus.n53 62.0763
R54 minus.n18 minus.n17 46.0096
R55 minus.n17 minus.n16 46.0096
R56 minus.n45 minus.n44 46.0096
R57 minus.n46 minus.n45 46.0096
R58 minus.n27 minus.n26 43.0884
R59 minus.n7 minus.n6 43.0884
R60 minus.n35 minus.n34 43.0884
R61 minus.n56 minus.n55 43.0884
R62 minus.n58 minus.n28 37.099
R63 minus.n26 minus.n25 29.9429
R64 minus.n9 minus.n6 29.9429
R65 minus.n37 minus.n34 29.9429
R66 minus.n55 minus.n54 29.9429
R67 minus.n19 minus.n18 27.0217
R68 minus.n16 minus.n15 27.0217
R69 minus.n44 minus.n43 27.0217
R70 minus.n48 minus.n46 27.0217
R71 minus.n24 minus.n23 10.955
R72 minus.n11 minus.n10 10.955
R73 minus.n39 minus.n38 10.955
R74 minus.n53 minus.n52 10.955
R75 minus.n3 minus.n1 8.03383
R76 minus.n12 minus.n4 8.03383
R77 minus.n40 minus.n32 8.03383
R78 minus.n47 minus.n30 8.03383
R79 minus.n58 minus.n57 6.51565
R80 minus.n28 minus.n0 0.189894
R81 minus.n22 minus.n0 0.189894
R82 minus.n22 minus.n21 0.189894
R83 minus.n21 minus.n20 0.189894
R84 minus.n20 minus.n2 0.189894
R85 minus.n14 minus.n2 0.189894
R86 minus.n14 minus.n13 0.189894
R87 minus.n13 minus.n5 0.189894
R88 minus.n8 minus.n5 0.189894
R89 minus.n36 minus.n33 0.189894
R90 minus.n41 minus.n33 0.189894
R91 minus.n42 minus.n41 0.189894
R92 minus.n42 minus.n31 0.189894
R93 minus.n49 minus.n31 0.189894
R94 minus.n50 minus.n49 0.189894
R95 minus.n51 minus.n50 0.189894
R96 minus.n51 minus.n29 0.189894
R97 minus.n57 minus.n29 0.189894
R98 minus minus.n58 0.188
R99 drain_right.n6 drain_right.n4 60.0956
R100 drain_right.n2 drain_right.n0 60.0956
R101 drain_right.n10 drain_right.n8 60.0956
R102 drain_right.n10 drain_right.n9 59.5527
R103 drain_right.n12 drain_right.n11 59.5527
R104 drain_right.n14 drain_right.n13 59.5527
R105 drain_right.n16 drain_right.n15 59.5527
R106 drain_right.n7 drain_right.n3 59.5525
R107 drain_right.n6 drain_right.n5 59.5525
R108 drain_right.n2 drain_right.n1 59.5525
R109 drain_right drain_right.n7 31.1587
R110 drain_right drain_right.n16 6.19632
R111 drain_right.n3 drain_right.t14 1.6505
R112 drain_right.n3 drain_right.t7 1.6505
R113 drain_right.n4 drain_right.t1 1.6505
R114 drain_right.n4 drain_right.t13 1.6505
R115 drain_right.n5 drain_right.t15 1.6505
R116 drain_right.n5 drain_right.t2 1.6505
R117 drain_right.n1 drain_right.t10 1.6505
R118 drain_right.n1 drain_right.t8 1.6505
R119 drain_right.n0 drain_right.t11 1.6505
R120 drain_right.n0 drain_right.t4 1.6505
R121 drain_right.n8 drain_right.t17 1.6505
R122 drain_right.n8 drain_right.t18 1.6505
R123 drain_right.n9 drain_right.t5 1.6505
R124 drain_right.n9 drain_right.t12 1.6505
R125 drain_right.n11 drain_right.t9 1.6505
R126 drain_right.n11 drain_right.t0 1.6505
R127 drain_right.n13 drain_right.t6 1.6505
R128 drain_right.n13 drain_right.t16 1.6505
R129 drain_right.n15 drain_right.t3 1.6505
R130 drain_right.n15 drain_right.t19 1.6505
R131 drain_right.n16 drain_right.n14 0.543603
R132 drain_right.n14 drain_right.n12 0.543603
R133 drain_right.n12 drain_right.n10 0.543603
R134 drain_right.n7 drain_right.n6 0.488257
R135 drain_right.n7 drain_right.n2 0.488257
R136 source.n554 source.n494 289.615
R137 source.n480 source.n420 289.615
R138 source.n414 source.n354 289.615
R139 source.n340 source.n280 289.615
R140 source.n60 source.n0 289.615
R141 source.n134 source.n74 289.615
R142 source.n200 source.n140 289.615
R143 source.n274 source.n214 289.615
R144 source.n514 source.n513 185
R145 source.n519 source.n518 185
R146 source.n521 source.n520 185
R147 source.n510 source.n509 185
R148 source.n527 source.n526 185
R149 source.n529 source.n528 185
R150 source.n506 source.n505 185
R151 source.n536 source.n535 185
R152 source.n537 source.n504 185
R153 source.n539 source.n538 185
R154 source.n502 source.n501 185
R155 source.n545 source.n544 185
R156 source.n547 source.n546 185
R157 source.n498 source.n497 185
R158 source.n553 source.n552 185
R159 source.n555 source.n554 185
R160 source.n440 source.n439 185
R161 source.n445 source.n444 185
R162 source.n447 source.n446 185
R163 source.n436 source.n435 185
R164 source.n453 source.n452 185
R165 source.n455 source.n454 185
R166 source.n432 source.n431 185
R167 source.n462 source.n461 185
R168 source.n463 source.n430 185
R169 source.n465 source.n464 185
R170 source.n428 source.n427 185
R171 source.n471 source.n470 185
R172 source.n473 source.n472 185
R173 source.n424 source.n423 185
R174 source.n479 source.n478 185
R175 source.n481 source.n480 185
R176 source.n374 source.n373 185
R177 source.n379 source.n378 185
R178 source.n381 source.n380 185
R179 source.n370 source.n369 185
R180 source.n387 source.n386 185
R181 source.n389 source.n388 185
R182 source.n366 source.n365 185
R183 source.n396 source.n395 185
R184 source.n397 source.n364 185
R185 source.n399 source.n398 185
R186 source.n362 source.n361 185
R187 source.n405 source.n404 185
R188 source.n407 source.n406 185
R189 source.n358 source.n357 185
R190 source.n413 source.n412 185
R191 source.n415 source.n414 185
R192 source.n300 source.n299 185
R193 source.n305 source.n304 185
R194 source.n307 source.n306 185
R195 source.n296 source.n295 185
R196 source.n313 source.n312 185
R197 source.n315 source.n314 185
R198 source.n292 source.n291 185
R199 source.n322 source.n321 185
R200 source.n323 source.n290 185
R201 source.n325 source.n324 185
R202 source.n288 source.n287 185
R203 source.n331 source.n330 185
R204 source.n333 source.n332 185
R205 source.n284 source.n283 185
R206 source.n339 source.n338 185
R207 source.n341 source.n340 185
R208 source.n61 source.n60 185
R209 source.n59 source.n58 185
R210 source.n4 source.n3 185
R211 source.n53 source.n52 185
R212 source.n51 source.n50 185
R213 source.n8 source.n7 185
R214 source.n45 source.n44 185
R215 source.n43 source.n10 185
R216 source.n42 source.n41 185
R217 source.n13 source.n11 185
R218 source.n36 source.n35 185
R219 source.n34 source.n33 185
R220 source.n17 source.n16 185
R221 source.n28 source.n27 185
R222 source.n26 source.n25 185
R223 source.n21 source.n20 185
R224 source.n135 source.n134 185
R225 source.n133 source.n132 185
R226 source.n78 source.n77 185
R227 source.n127 source.n126 185
R228 source.n125 source.n124 185
R229 source.n82 source.n81 185
R230 source.n119 source.n118 185
R231 source.n117 source.n84 185
R232 source.n116 source.n115 185
R233 source.n87 source.n85 185
R234 source.n110 source.n109 185
R235 source.n108 source.n107 185
R236 source.n91 source.n90 185
R237 source.n102 source.n101 185
R238 source.n100 source.n99 185
R239 source.n95 source.n94 185
R240 source.n201 source.n200 185
R241 source.n199 source.n198 185
R242 source.n144 source.n143 185
R243 source.n193 source.n192 185
R244 source.n191 source.n190 185
R245 source.n148 source.n147 185
R246 source.n185 source.n184 185
R247 source.n183 source.n150 185
R248 source.n182 source.n181 185
R249 source.n153 source.n151 185
R250 source.n176 source.n175 185
R251 source.n174 source.n173 185
R252 source.n157 source.n156 185
R253 source.n168 source.n167 185
R254 source.n166 source.n165 185
R255 source.n161 source.n160 185
R256 source.n275 source.n274 185
R257 source.n273 source.n272 185
R258 source.n218 source.n217 185
R259 source.n267 source.n266 185
R260 source.n265 source.n264 185
R261 source.n222 source.n221 185
R262 source.n259 source.n258 185
R263 source.n257 source.n224 185
R264 source.n256 source.n255 185
R265 source.n227 source.n225 185
R266 source.n250 source.n249 185
R267 source.n248 source.n247 185
R268 source.n231 source.n230 185
R269 source.n242 source.n241 185
R270 source.n240 source.n239 185
R271 source.n235 source.n234 185
R272 source.n515 source.t34 149.524
R273 source.n441 source.t36 149.524
R274 source.n375 source.t15 149.524
R275 source.n301 source.t6 149.524
R276 source.n22 source.t12 149.524
R277 source.n96 source.t11 149.524
R278 source.n162 source.t26 149.524
R279 source.n236 source.t30 149.524
R280 source.n519 source.n513 104.615
R281 source.n520 source.n519 104.615
R282 source.n520 source.n509 104.615
R283 source.n527 source.n509 104.615
R284 source.n528 source.n527 104.615
R285 source.n528 source.n505 104.615
R286 source.n536 source.n505 104.615
R287 source.n537 source.n536 104.615
R288 source.n538 source.n537 104.615
R289 source.n538 source.n501 104.615
R290 source.n545 source.n501 104.615
R291 source.n546 source.n545 104.615
R292 source.n546 source.n497 104.615
R293 source.n553 source.n497 104.615
R294 source.n554 source.n553 104.615
R295 source.n445 source.n439 104.615
R296 source.n446 source.n445 104.615
R297 source.n446 source.n435 104.615
R298 source.n453 source.n435 104.615
R299 source.n454 source.n453 104.615
R300 source.n454 source.n431 104.615
R301 source.n462 source.n431 104.615
R302 source.n463 source.n462 104.615
R303 source.n464 source.n463 104.615
R304 source.n464 source.n427 104.615
R305 source.n471 source.n427 104.615
R306 source.n472 source.n471 104.615
R307 source.n472 source.n423 104.615
R308 source.n479 source.n423 104.615
R309 source.n480 source.n479 104.615
R310 source.n379 source.n373 104.615
R311 source.n380 source.n379 104.615
R312 source.n380 source.n369 104.615
R313 source.n387 source.n369 104.615
R314 source.n388 source.n387 104.615
R315 source.n388 source.n365 104.615
R316 source.n396 source.n365 104.615
R317 source.n397 source.n396 104.615
R318 source.n398 source.n397 104.615
R319 source.n398 source.n361 104.615
R320 source.n405 source.n361 104.615
R321 source.n406 source.n405 104.615
R322 source.n406 source.n357 104.615
R323 source.n413 source.n357 104.615
R324 source.n414 source.n413 104.615
R325 source.n305 source.n299 104.615
R326 source.n306 source.n305 104.615
R327 source.n306 source.n295 104.615
R328 source.n313 source.n295 104.615
R329 source.n314 source.n313 104.615
R330 source.n314 source.n291 104.615
R331 source.n322 source.n291 104.615
R332 source.n323 source.n322 104.615
R333 source.n324 source.n323 104.615
R334 source.n324 source.n287 104.615
R335 source.n331 source.n287 104.615
R336 source.n332 source.n331 104.615
R337 source.n332 source.n283 104.615
R338 source.n339 source.n283 104.615
R339 source.n340 source.n339 104.615
R340 source.n60 source.n59 104.615
R341 source.n59 source.n3 104.615
R342 source.n52 source.n3 104.615
R343 source.n52 source.n51 104.615
R344 source.n51 source.n7 104.615
R345 source.n44 source.n7 104.615
R346 source.n44 source.n43 104.615
R347 source.n43 source.n42 104.615
R348 source.n42 source.n11 104.615
R349 source.n35 source.n11 104.615
R350 source.n35 source.n34 104.615
R351 source.n34 source.n16 104.615
R352 source.n27 source.n16 104.615
R353 source.n27 source.n26 104.615
R354 source.n26 source.n20 104.615
R355 source.n134 source.n133 104.615
R356 source.n133 source.n77 104.615
R357 source.n126 source.n77 104.615
R358 source.n126 source.n125 104.615
R359 source.n125 source.n81 104.615
R360 source.n118 source.n81 104.615
R361 source.n118 source.n117 104.615
R362 source.n117 source.n116 104.615
R363 source.n116 source.n85 104.615
R364 source.n109 source.n85 104.615
R365 source.n109 source.n108 104.615
R366 source.n108 source.n90 104.615
R367 source.n101 source.n90 104.615
R368 source.n101 source.n100 104.615
R369 source.n100 source.n94 104.615
R370 source.n200 source.n199 104.615
R371 source.n199 source.n143 104.615
R372 source.n192 source.n143 104.615
R373 source.n192 source.n191 104.615
R374 source.n191 source.n147 104.615
R375 source.n184 source.n147 104.615
R376 source.n184 source.n183 104.615
R377 source.n183 source.n182 104.615
R378 source.n182 source.n151 104.615
R379 source.n175 source.n151 104.615
R380 source.n175 source.n174 104.615
R381 source.n174 source.n156 104.615
R382 source.n167 source.n156 104.615
R383 source.n167 source.n166 104.615
R384 source.n166 source.n160 104.615
R385 source.n274 source.n273 104.615
R386 source.n273 source.n217 104.615
R387 source.n266 source.n217 104.615
R388 source.n266 source.n265 104.615
R389 source.n265 source.n221 104.615
R390 source.n258 source.n221 104.615
R391 source.n258 source.n257 104.615
R392 source.n257 source.n256 104.615
R393 source.n256 source.n225 104.615
R394 source.n249 source.n225 104.615
R395 source.n249 source.n248 104.615
R396 source.n248 source.n230 104.615
R397 source.n241 source.n230 104.615
R398 source.n241 source.n240 104.615
R399 source.n240 source.n234 104.615
R400 source.t34 source.n513 52.3082
R401 source.t36 source.n439 52.3082
R402 source.t15 source.n373 52.3082
R403 source.t6 source.n299 52.3082
R404 source.t12 source.n20 52.3082
R405 source.t11 source.n94 52.3082
R406 source.t26 source.n160 52.3082
R407 source.t30 source.n234 52.3082
R408 source.n67 source.n66 42.8739
R409 source.n69 source.n68 42.8739
R410 source.n71 source.n70 42.8739
R411 source.n73 source.n72 42.8739
R412 source.n207 source.n206 42.8739
R413 source.n209 source.n208 42.8739
R414 source.n211 source.n210 42.8739
R415 source.n213 source.n212 42.8739
R416 source.n493 source.n492 42.8737
R417 source.n491 source.n490 42.8737
R418 source.n489 source.n488 42.8737
R419 source.n487 source.n486 42.8737
R420 source.n353 source.n352 42.8737
R421 source.n351 source.n350 42.8737
R422 source.n349 source.n348 42.8737
R423 source.n347 source.n346 42.8737
R424 source.n559 source.n558 29.8581
R425 source.n485 source.n484 29.8581
R426 source.n419 source.n418 29.8581
R427 source.n345 source.n344 29.8581
R428 source.n65 source.n64 29.8581
R429 source.n139 source.n138 29.8581
R430 source.n205 source.n204 29.8581
R431 source.n279 source.n278 29.8581
R432 source.n345 source.n279 21.8308
R433 source.n560 source.n65 16.2963
R434 source.n539 source.n504 13.1884
R435 source.n465 source.n430 13.1884
R436 source.n399 source.n364 13.1884
R437 source.n325 source.n290 13.1884
R438 source.n45 source.n10 13.1884
R439 source.n119 source.n84 13.1884
R440 source.n185 source.n150 13.1884
R441 source.n259 source.n224 13.1884
R442 source.n535 source.n534 12.8005
R443 source.n540 source.n502 12.8005
R444 source.n461 source.n460 12.8005
R445 source.n466 source.n428 12.8005
R446 source.n395 source.n394 12.8005
R447 source.n400 source.n362 12.8005
R448 source.n321 source.n320 12.8005
R449 source.n326 source.n288 12.8005
R450 source.n46 source.n8 12.8005
R451 source.n41 source.n12 12.8005
R452 source.n120 source.n82 12.8005
R453 source.n115 source.n86 12.8005
R454 source.n186 source.n148 12.8005
R455 source.n181 source.n152 12.8005
R456 source.n260 source.n222 12.8005
R457 source.n255 source.n226 12.8005
R458 source.n533 source.n506 12.0247
R459 source.n544 source.n543 12.0247
R460 source.n459 source.n432 12.0247
R461 source.n470 source.n469 12.0247
R462 source.n393 source.n366 12.0247
R463 source.n404 source.n403 12.0247
R464 source.n319 source.n292 12.0247
R465 source.n330 source.n329 12.0247
R466 source.n50 source.n49 12.0247
R467 source.n40 source.n13 12.0247
R468 source.n124 source.n123 12.0247
R469 source.n114 source.n87 12.0247
R470 source.n190 source.n189 12.0247
R471 source.n180 source.n153 12.0247
R472 source.n264 source.n263 12.0247
R473 source.n254 source.n227 12.0247
R474 source.n530 source.n529 11.249
R475 source.n547 source.n500 11.249
R476 source.n456 source.n455 11.249
R477 source.n473 source.n426 11.249
R478 source.n390 source.n389 11.249
R479 source.n407 source.n360 11.249
R480 source.n316 source.n315 11.249
R481 source.n333 source.n286 11.249
R482 source.n53 source.n6 11.249
R483 source.n37 source.n36 11.249
R484 source.n127 source.n80 11.249
R485 source.n111 source.n110 11.249
R486 source.n193 source.n146 11.249
R487 source.n177 source.n176 11.249
R488 source.n267 source.n220 11.249
R489 source.n251 source.n250 11.249
R490 source.n526 source.n508 10.4732
R491 source.n548 source.n498 10.4732
R492 source.n452 source.n434 10.4732
R493 source.n474 source.n424 10.4732
R494 source.n386 source.n368 10.4732
R495 source.n408 source.n358 10.4732
R496 source.n312 source.n294 10.4732
R497 source.n334 source.n284 10.4732
R498 source.n54 source.n4 10.4732
R499 source.n33 source.n15 10.4732
R500 source.n128 source.n78 10.4732
R501 source.n107 source.n89 10.4732
R502 source.n194 source.n144 10.4732
R503 source.n173 source.n155 10.4732
R504 source.n268 source.n218 10.4732
R505 source.n247 source.n229 10.4732
R506 source.n515 source.n514 10.2747
R507 source.n441 source.n440 10.2747
R508 source.n375 source.n374 10.2747
R509 source.n301 source.n300 10.2747
R510 source.n22 source.n21 10.2747
R511 source.n96 source.n95 10.2747
R512 source.n162 source.n161 10.2747
R513 source.n236 source.n235 10.2747
R514 source.n525 source.n510 9.69747
R515 source.n552 source.n551 9.69747
R516 source.n451 source.n436 9.69747
R517 source.n478 source.n477 9.69747
R518 source.n385 source.n370 9.69747
R519 source.n412 source.n411 9.69747
R520 source.n311 source.n296 9.69747
R521 source.n338 source.n337 9.69747
R522 source.n58 source.n57 9.69747
R523 source.n32 source.n17 9.69747
R524 source.n132 source.n131 9.69747
R525 source.n106 source.n91 9.69747
R526 source.n198 source.n197 9.69747
R527 source.n172 source.n157 9.69747
R528 source.n272 source.n271 9.69747
R529 source.n246 source.n231 9.69747
R530 source.n558 source.n557 9.45567
R531 source.n484 source.n483 9.45567
R532 source.n418 source.n417 9.45567
R533 source.n344 source.n343 9.45567
R534 source.n64 source.n63 9.45567
R535 source.n138 source.n137 9.45567
R536 source.n204 source.n203 9.45567
R537 source.n278 source.n277 9.45567
R538 source.n557 source.n556 9.3005
R539 source.n496 source.n495 9.3005
R540 source.n551 source.n550 9.3005
R541 source.n549 source.n548 9.3005
R542 source.n500 source.n499 9.3005
R543 source.n543 source.n542 9.3005
R544 source.n541 source.n540 9.3005
R545 source.n517 source.n516 9.3005
R546 source.n512 source.n511 9.3005
R547 source.n523 source.n522 9.3005
R548 source.n525 source.n524 9.3005
R549 source.n508 source.n507 9.3005
R550 source.n531 source.n530 9.3005
R551 source.n533 source.n532 9.3005
R552 source.n534 source.n503 9.3005
R553 source.n483 source.n482 9.3005
R554 source.n422 source.n421 9.3005
R555 source.n477 source.n476 9.3005
R556 source.n475 source.n474 9.3005
R557 source.n426 source.n425 9.3005
R558 source.n469 source.n468 9.3005
R559 source.n467 source.n466 9.3005
R560 source.n443 source.n442 9.3005
R561 source.n438 source.n437 9.3005
R562 source.n449 source.n448 9.3005
R563 source.n451 source.n450 9.3005
R564 source.n434 source.n433 9.3005
R565 source.n457 source.n456 9.3005
R566 source.n459 source.n458 9.3005
R567 source.n460 source.n429 9.3005
R568 source.n417 source.n416 9.3005
R569 source.n356 source.n355 9.3005
R570 source.n411 source.n410 9.3005
R571 source.n409 source.n408 9.3005
R572 source.n360 source.n359 9.3005
R573 source.n403 source.n402 9.3005
R574 source.n401 source.n400 9.3005
R575 source.n377 source.n376 9.3005
R576 source.n372 source.n371 9.3005
R577 source.n383 source.n382 9.3005
R578 source.n385 source.n384 9.3005
R579 source.n368 source.n367 9.3005
R580 source.n391 source.n390 9.3005
R581 source.n393 source.n392 9.3005
R582 source.n394 source.n363 9.3005
R583 source.n343 source.n342 9.3005
R584 source.n282 source.n281 9.3005
R585 source.n337 source.n336 9.3005
R586 source.n335 source.n334 9.3005
R587 source.n286 source.n285 9.3005
R588 source.n329 source.n328 9.3005
R589 source.n327 source.n326 9.3005
R590 source.n303 source.n302 9.3005
R591 source.n298 source.n297 9.3005
R592 source.n309 source.n308 9.3005
R593 source.n311 source.n310 9.3005
R594 source.n294 source.n293 9.3005
R595 source.n317 source.n316 9.3005
R596 source.n319 source.n318 9.3005
R597 source.n320 source.n289 9.3005
R598 source.n24 source.n23 9.3005
R599 source.n19 source.n18 9.3005
R600 source.n30 source.n29 9.3005
R601 source.n32 source.n31 9.3005
R602 source.n15 source.n14 9.3005
R603 source.n38 source.n37 9.3005
R604 source.n40 source.n39 9.3005
R605 source.n12 source.n9 9.3005
R606 source.n63 source.n62 9.3005
R607 source.n2 source.n1 9.3005
R608 source.n57 source.n56 9.3005
R609 source.n55 source.n54 9.3005
R610 source.n6 source.n5 9.3005
R611 source.n49 source.n48 9.3005
R612 source.n47 source.n46 9.3005
R613 source.n98 source.n97 9.3005
R614 source.n93 source.n92 9.3005
R615 source.n104 source.n103 9.3005
R616 source.n106 source.n105 9.3005
R617 source.n89 source.n88 9.3005
R618 source.n112 source.n111 9.3005
R619 source.n114 source.n113 9.3005
R620 source.n86 source.n83 9.3005
R621 source.n137 source.n136 9.3005
R622 source.n76 source.n75 9.3005
R623 source.n131 source.n130 9.3005
R624 source.n129 source.n128 9.3005
R625 source.n80 source.n79 9.3005
R626 source.n123 source.n122 9.3005
R627 source.n121 source.n120 9.3005
R628 source.n164 source.n163 9.3005
R629 source.n159 source.n158 9.3005
R630 source.n170 source.n169 9.3005
R631 source.n172 source.n171 9.3005
R632 source.n155 source.n154 9.3005
R633 source.n178 source.n177 9.3005
R634 source.n180 source.n179 9.3005
R635 source.n152 source.n149 9.3005
R636 source.n203 source.n202 9.3005
R637 source.n142 source.n141 9.3005
R638 source.n197 source.n196 9.3005
R639 source.n195 source.n194 9.3005
R640 source.n146 source.n145 9.3005
R641 source.n189 source.n188 9.3005
R642 source.n187 source.n186 9.3005
R643 source.n238 source.n237 9.3005
R644 source.n233 source.n232 9.3005
R645 source.n244 source.n243 9.3005
R646 source.n246 source.n245 9.3005
R647 source.n229 source.n228 9.3005
R648 source.n252 source.n251 9.3005
R649 source.n254 source.n253 9.3005
R650 source.n226 source.n223 9.3005
R651 source.n277 source.n276 9.3005
R652 source.n216 source.n215 9.3005
R653 source.n271 source.n270 9.3005
R654 source.n269 source.n268 9.3005
R655 source.n220 source.n219 9.3005
R656 source.n263 source.n262 9.3005
R657 source.n261 source.n260 9.3005
R658 source.n522 source.n521 8.92171
R659 source.n555 source.n496 8.92171
R660 source.n448 source.n447 8.92171
R661 source.n481 source.n422 8.92171
R662 source.n382 source.n381 8.92171
R663 source.n415 source.n356 8.92171
R664 source.n308 source.n307 8.92171
R665 source.n341 source.n282 8.92171
R666 source.n61 source.n2 8.92171
R667 source.n29 source.n28 8.92171
R668 source.n135 source.n76 8.92171
R669 source.n103 source.n102 8.92171
R670 source.n201 source.n142 8.92171
R671 source.n169 source.n168 8.92171
R672 source.n275 source.n216 8.92171
R673 source.n243 source.n242 8.92171
R674 source.n518 source.n512 8.14595
R675 source.n556 source.n494 8.14595
R676 source.n444 source.n438 8.14595
R677 source.n482 source.n420 8.14595
R678 source.n378 source.n372 8.14595
R679 source.n416 source.n354 8.14595
R680 source.n304 source.n298 8.14595
R681 source.n342 source.n280 8.14595
R682 source.n62 source.n0 8.14595
R683 source.n25 source.n19 8.14595
R684 source.n136 source.n74 8.14595
R685 source.n99 source.n93 8.14595
R686 source.n202 source.n140 8.14595
R687 source.n165 source.n159 8.14595
R688 source.n276 source.n214 8.14595
R689 source.n239 source.n233 8.14595
R690 source.n517 source.n514 7.3702
R691 source.n443 source.n440 7.3702
R692 source.n377 source.n374 7.3702
R693 source.n303 source.n300 7.3702
R694 source.n24 source.n21 7.3702
R695 source.n98 source.n95 7.3702
R696 source.n164 source.n161 7.3702
R697 source.n238 source.n235 7.3702
R698 source.n518 source.n517 5.81868
R699 source.n558 source.n494 5.81868
R700 source.n444 source.n443 5.81868
R701 source.n484 source.n420 5.81868
R702 source.n378 source.n377 5.81868
R703 source.n418 source.n354 5.81868
R704 source.n304 source.n303 5.81868
R705 source.n344 source.n280 5.81868
R706 source.n64 source.n0 5.81868
R707 source.n25 source.n24 5.81868
R708 source.n138 source.n74 5.81868
R709 source.n99 source.n98 5.81868
R710 source.n204 source.n140 5.81868
R711 source.n165 source.n164 5.81868
R712 source.n278 source.n214 5.81868
R713 source.n239 source.n238 5.81868
R714 source.n560 source.n559 5.53498
R715 source.n521 source.n512 5.04292
R716 source.n556 source.n555 5.04292
R717 source.n447 source.n438 5.04292
R718 source.n482 source.n481 5.04292
R719 source.n381 source.n372 5.04292
R720 source.n416 source.n415 5.04292
R721 source.n307 source.n298 5.04292
R722 source.n342 source.n341 5.04292
R723 source.n62 source.n61 5.04292
R724 source.n28 source.n19 5.04292
R725 source.n136 source.n135 5.04292
R726 source.n102 source.n93 5.04292
R727 source.n202 source.n201 5.04292
R728 source.n168 source.n159 5.04292
R729 source.n276 source.n275 5.04292
R730 source.n242 source.n233 5.04292
R731 source.n522 source.n510 4.26717
R732 source.n552 source.n496 4.26717
R733 source.n448 source.n436 4.26717
R734 source.n478 source.n422 4.26717
R735 source.n382 source.n370 4.26717
R736 source.n412 source.n356 4.26717
R737 source.n308 source.n296 4.26717
R738 source.n338 source.n282 4.26717
R739 source.n58 source.n2 4.26717
R740 source.n29 source.n17 4.26717
R741 source.n132 source.n76 4.26717
R742 source.n103 source.n91 4.26717
R743 source.n198 source.n142 4.26717
R744 source.n169 source.n157 4.26717
R745 source.n272 source.n216 4.26717
R746 source.n243 source.n231 4.26717
R747 source.n526 source.n525 3.49141
R748 source.n551 source.n498 3.49141
R749 source.n452 source.n451 3.49141
R750 source.n477 source.n424 3.49141
R751 source.n386 source.n385 3.49141
R752 source.n411 source.n358 3.49141
R753 source.n312 source.n311 3.49141
R754 source.n337 source.n284 3.49141
R755 source.n57 source.n4 3.49141
R756 source.n33 source.n32 3.49141
R757 source.n131 source.n78 3.49141
R758 source.n107 source.n106 3.49141
R759 source.n197 source.n144 3.49141
R760 source.n173 source.n172 3.49141
R761 source.n271 source.n218 3.49141
R762 source.n247 source.n246 3.49141
R763 source.n516 source.n515 2.84303
R764 source.n442 source.n441 2.84303
R765 source.n376 source.n375 2.84303
R766 source.n302 source.n301 2.84303
R767 source.n23 source.n22 2.84303
R768 source.n97 source.n96 2.84303
R769 source.n163 source.n162 2.84303
R770 source.n237 source.n236 2.84303
R771 source.n529 source.n508 2.71565
R772 source.n548 source.n547 2.71565
R773 source.n455 source.n434 2.71565
R774 source.n474 source.n473 2.71565
R775 source.n389 source.n368 2.71565
R776 source.n408 source.n407 2.71565
R777 source.n315 source.n294 2.71565
R778 source.n334 source.n333 2.71565
R779 source.n54 source.n53 2.71565
R780 source.n36 source.n15 2.71565
R781 source.n128 source.n127 2.71565
R782 source.n110 source.n89 2.71565
R783 source.n194 source.n193 2.71565
R784 source.n176 source.n155 2.71565
R785 source.n268 source.n267 2.71565
R786 source.n250 source.n229 2.71565
R787 source.n530 source.n506 1.93989
R788 source.n544 source.n500 1.93989
R789 source.n456 source.n432 1.93989
R790 source.n470 source.n426 1.93989
R791 source.n390 source.n366 1.93989
R792 source.n404 source.n360 1.93989
R793 source.n316 source.n292 1.93989
R794 source.n330 source.n286 1.93989
R795 source.n50 source.n6 1.93989
R796 source.n37 source.n13 1.93989
R797 source.n124 source.n80 1.93989
R798 source.n111 source.n87 1.93989
R799 source.n190 source.n146 1.93989
R800 source.n177 source.n153 1.93989
R801 source.n264 source.n220 1.93989
R802 source.n251 source.n227 1.93989
R803 source.n492 source.t22 1.6505
R804 source.n492 source.t23 1.6505
R805 source.n490 source.t21 1.6505
R806 source.n490 source.t29 1.6505
R807 source.n488 source.t25 1.6505
R808 source.n488 source.t28 1.6505
R809 source.n486 source.t24 1.6505
R810 source.n486 source.t37 1.6505
R811 source.n352 source.t5 1.6505
R812 source.n352 source.t9 1.6505
R813 source.n350 source.t4 1.6505
R814 source.n350 source.t39 1.6505
R815 source.n348 source.t13 1.6505
R816 source.n348 source.t3 1.6505
R817 source.n346 source.t1 1.6505
R818 source.n346 source.t10 1.6505
R819 source.n66 source.t8 1.6505
R820 source.n66 source.t0 1.6505
R821 source.n68 source.t2 1.6505
R822 source.n68 source.t7 1.6505
R823 source.n70 source.t17 1.6505
R824 source.n70 source.t14 1.6505
R825 source.n72 source.t38 1.6505
R826 source.n72 source.t16 1.6505
R827 source.n206 source.t33 1.6505
R828 source.n206 source.t19 1.6505
R829 source.n208 source.t20 1.6505
R830 source.n208 source.t27 1.6505
R831 source.n210 source.t31 1.6505
R832 source.n210 source.t35 1.6505
R833 source.n212 source.t32 1.6505
R834 source.n212 source.t18 1.6505
R835 source.n535 source.n533 1.16414
R836 source.n543 source.n502 1.16414
R837 source.n461 source.n459 1.16414
R838 source.n469 source.n428 1.16414
R839 source.n395 source.n393 1.16414
R840 source.n403 source.n362 1.16414
R841 source.n321 source.n319 1.16414
R842 source.n329 source.n288 1.16414
R843 source.n49 source.n8 1.16414
R844 source.n41 source.n40 1.16414
R845 source.n123 source.n82 1.16414
R846 source.n115 source.n114 1.16414
R847 source.n189 source.n148 1.16414
R848 source.n181 source.n180 1.16414
R849 source.n263 source.n222 1.16414
R850 source.n255 source.n254 1.16414
R851 source.n279 source.n213 0.543603
R852 source.n213 source.n211 0.543603
R853 source.n211 source.n209 0.543603
R854 source.n209 source.n207 0.543603
R855 source.n207 source.n205 0.543603
R856 source.n139 source.n73 0.543603
R857 source.n73 source.n71 0.543603
R858 source.n71 source.n69 0.543603
R859 source.n69 source.n67 0.543603
R860 source.n67 source.n65 0.543603
R861 source.n347 source.n345 0.543603
R862 source.n349 source.n347 0.543603
R863 source.n351 source.n349 0.543603
R864 source.n353 source.n351 0.543603
R865 source.n419 source.n353 0.543603
R866 source.n487 source.n485 0.543603
R867 source.n489 source.n487 0.543603
R868 source.n491 source.n489 0.543603
R869 source.n493 source.n491 0.543603
R870 source.n559 source.n493 0.543603
R871 source.n205 source.n139 0.470328
R872 source.n485 source.n419 0.470328
R873 source.n534 source.n504 0.388379
R874 source.n540 source.n539 0.388379
R875 source.n460 source.n430 0.388379
R876 source.n466 source.n465 0.388379
R877 source.n394 source.n364 0.388379
R878 source.n400 source.n399 0.388379
R879 source.n320 source.n290 0.388379
R880 source.n326 source.n325 0.388379
R881 source.n46 source.n45 0.388379
R882 source.n12 source.n10 0.388379
R883 source.n120 source.n119 0.388379
R884 source.n86 source.n84 0.388379
R885 source.n186 source.n185 0.388379
R886 source.n152 source.n150 0.388379
R887 source.n260 source.n259 0.388379
R888 source.n226 source.n224 0.388379
R889 source source.n560 0.188
R890 source.n516 source.n511 0.155672
R891 source.n523 source.n511 0.155672
R892 source.n524 source.n523 0.155672
R893 source.n524 source.n507 0.155672
R894 source.n531 source.n507 0.155672
R895 source.n532 source.n531 0.155672
R896 source.n532 source.n503 0.155672
R897 source.n541 source.n503 0.155672
R898 source.n542 source.n541 0.155672
R899 source.n542 source.n499 0.155672
R900 source.n549 source.n499 0.155672
R901 source.n550 source.n549 0.155672
R902 source.n550 source.n495 0.155672
R903 source.n557 source.n495 0.155672
R904 source.n442 source.n437 0.155672
R905 source.n449 source.n437 0.155672
R906 source.n450 source.n449 0.155672
R907 source.n450 source.n433 0.155672
R908 source.n457 source.n433 0.155672
R909 source.n458 source.n457 0.155672
R910 source.n458 source.n429 0.155672
R911 source.n467 source.n429 0.155672
R912 source.n468 source.n467 0.155672
R913 source.n468 source.n425 0.155672
R914 source.n475 source.n425 0.155672
R915 source.n476 source.n475 0.155672
R916 source.n476 source.n421 0.155672
R917 source.n483 source.n421 0.155672
R918 source.n376 source.n371 0.155672
R919 source.n383 source.n371 0.155672
R920 source.n384 source.n383 0.155672
R921 source.n384 source.n367 0.155672
R922 source.n391 source.n367 0.155672
R923 source.n392 source.n391 0.155672
R924 source.n392 source.n363 0.155672
R925 source.n401 source.n363 0.155672
R926 source.n402 source.n401 0.155672
R927 source.n402 source.n359 0.155672
R928 source.n409 source.n359 0.155672
R929 source.n410 source.n409 0.155672
R930 source.n410 source.n355 0.155672
R931 source.n417 source.n355 0.155672
R932 source.n302 source.n297 0.155672
R933 source.n309 source.n297 0.155672
R934 source.n310 source.n309 0.155672
R935 source.n310 source.n293 0.155672
R936 source.n317 source.n293 0.155672
R937 source.n318 source.n317 0.155672
R938 source.n318 source.n289 0.155672
R939 source.n327 source.n289 0.155672
R940 source.n328 source.n327 0.155672
R941 source.n328 source.n285 0.155672
R942 source.n335 source.n285 0.155672
R943 source.n336 source.n335 0.155672
R944 source.n336 source.n281 0.155672
R945 source.n343 source.n281 0.155672
R946 source.n63 source.n1 0.155672
R947 source.n56 source.n1 0.155672
R948 source.n56 source.n55 0.155672
R949 source.n55 source.n5 0.155672
R950 source.n48 source.n5 0.155672
R951 source.n48 source.n47 0.155672
R952 source.n47 source.n9 0.155672
R953 source.n39 source.n9 0.155672
R954 source.n39 source.n38 0.155672
R955 source.n38 source.n14 0.155672
R956 source.n31 source.n14 0.155672
R957 source.n31 source.n30 0.155672
R958 source.n30 source.n18 0.155672
R959 source.n23 source.n18 0.155672
R960 source.n137 source.n75 0.155672
R961 source.n130 source.n75 0.155672
R962 source.n130 source.n129 0.155672
R963 source.n129 source.n79 0.155672
R964 source.n122 source.n79 0.155672
R965 source.n122 source.n121 0.155672
R966 source.n121 source.n83 0.155672
R967 source.n113 source.n83 0.155672
R968 source.n113 source.n112 0.155672
R969 source.n112 source.n88 0.155672
R970 source.n105 source.n88 0.155672
R971 source.n105 source.n104 0.155672
R972 source.n104 source.n92 0.155672
R973 source.n97 source.n92 0.155672
R974 source.n203 source.n141 0.155672
R975 source.n196 source.n141 0.155672
R976 source.n196 source.n195 0.155672
R977 source.n195 source.n145 0.155672
R978 source.n188 source.n145 0.155672
R979 source.n188 source.n187 0.155672
R980 source.n187 source.n149 0.155672
R981 source.n179 source.n149 0.155672
R982 source.n179 source.n178 0.155672
R983 source.n178 source.n154 0.155672
R984 source.n171 source.n154 0.155672
R985 source.n171 source.n170 0.155672
R986 source.n170 source.n158 0.155672
R987 source.n163 source.n158 0.155672
R988 source.n277 source.n215 0.155672
R989 source.n270 source.n215 0.155672
R990 source.n270 source.n269 0.155672
R991 source.n269 source.n219 0.155672
R992 source.n262 source.n219 0.155672
R993 source.n262 source.n261 0.155672
R994 source.n261 source.n223 0.155672
R995 source.n253 source.n223 0.155672
R996 source.n253 source.n252 0.155672
R997 source.n252 source.n228 0.155672
R998 source.n245 source.n228 0.155672
R999 source.n245 source.n244 0.155672
R1000 source.n244 source.n232 0.155672
R1001 source.n237 source.n232 0.155672
R1002 plus.n6 plus.t3 1117.36
R1003 plus.n27 plus.t15 1117.36
R1004 plus.n36 plus.t16 1117.36
R1005 plus.n56 plus.t14 1117.36
R1006 plus.n5 plus.t7 1068.43
R1007 plus.n9 plus.t12 1068.43
R1008 plus.n3 plus.t19 1068.43
R1009 plus.n15 plus.t5 1068.43
R1010 plus.n17 plus.t11 1068.43
R1011 plus.n18 plus.t18 1068.43
R1012 plus.n24 plus.t0 1068.43
R1013 plus.n26 plus.t10 1068.43
R1014 plus.n35 plus.t6 1068.43
R1015 plus.n39 plus.t17 1068.43
R1016 plus.n33 plus.t8 1068.43
R1017 plus.n45 plus.t2 1068.43
R1018 plus.n47 plus.t9 1068.43
R1019 plus.n32 plus.t4 1068.43
R1020 plus.n53 plus.t13 1068.43
R1021 plus.n55 plus.t1 1068.43
R1022 plus.n7 plus.n6 161.489
R1023 plus.n37 plus.n36 161.489
R1024 plus.n8 plus.n7 161.3
R1025 plus.n10 plus.n4 161.3
R1026 plus.n12 plus.n11 161.3
R1027 plus.n14 plus.n13 161.3
R1028 plus.n16 plus.n2 161.3
R1029 plus.n20 plus.n19 161.3
R1030 plus.n21 plus.n1 161.3
R1031 plus.n23 plus.n22 161.3
R1032 plus.n25 plus.n0 161.3
R1033 plus.n28 plus.n27 161.3
R1034 plus.n38 plus.n37 161.3
R1035 plus.n40 plus.n34 161.3
R1036 plus.n42 plus.n41 161.3
R1037 plus.n44 plus.n43 161.3
R1038 plus.n46 plus.n31 161.3
R1039 plus.n49 plus.n48 161.3
R1040 plus.n50 plus.n30 161.3
R1041 plus.n52 plus.n51 161.3
R1042 plus.n54 plus.n29 161.3
R1043 plus.n57 plus.n56 161.3
R1044 plus.n11 plus.n10 73.0308
R1045 plus.n23 plus.n1 73.0308
R1046 plus.n52 plus.n30 73.0308
R1047 plus.n41 plus.n40 73.0308
R1048 plus.n14 plus.n3 64.9975
R1049 plus.n19 plus.n18 64.9975
R1050 plus.n48 plus.n32 64.9975
R1051 plus.n44 plus.n33 64.9975
R1052 plus.n9 plus.n8 62.0763
R1053 plus.n25 plus.n24 62.0763
R1054 plus.n54 plus.n53 62.0763
R1055 plus.n39 plus.n38 62.0763
R1056 plus.n16 plus.n15 46.0096
R1057 plus.n17 plus.n16 46.0096
R1058 plus.n47 plus.n46 46.0096
R1059 plus.n46 plus.n45 46.0096
R1060 plus.n6 plus.n5 43.0884
R1061 plus.n27 plus.n26 43.0884
R1062 plus.n56 plus.n55 43.0884
R1063 plus.n36 plus.n35 43.0884
R1064 plus plus.n57 30.9801
R1065 plus.n8 plus.n5 29.9429
R1066 plus.n26 plus.n25 29.9429
R1067 plus.n55 plus.n54 29.9429
R1068 plus.n38 plus.n35 29.9429
R1069 plus.n15 plus.n14 27.0217
R1070 plus.n19 plus.n17 27.0217
R1071 plus.n48 plus.n47 27.0217
R1072 plus.n45 plus.n44 27.0217
R1073 plus plus.n28 12.1596
R1074 plus.n10 plus.n9 10.955
R1075 plus.n24 plus.n23 10.955
R1076 plus.n53 plus.n52 10.955
R1077 plus.n40 plus.n39 10.955
R1078 plus.n11 plus.n3 8.03383
R1079 plus.n18 plus.n1 8.03383
R1080 plus.n32 plus.n30 8.03383
R1081 plus.n41 plus.n33 8.03383
R1082 plus.n7 plus.n4 0.189894
R1083 plus.n12 plus.n4 0.189894
R1084 plus.n13 plus.n12 0.189894
R1085 plus.n13 plus.n2 0.189894
R1086 plus.n20 plus.n2 0.189894
R1087 plus.n21 plus.n20 0.189894
R1088 plus.n22 plus.n21 0.189894
R1089 plus.n22 plus.n0 0.189894
R1090 plus.n28 plus.n0 0.189894
R1091 plus.n57 plus.n29 0.189894
R1092 plus.n51 plus.n29 0.189894
R1093 plus.n51 plus.n50 0.189894
R1094 plus.n50 plus.n49 0.189894
R1095 plus.n49 plus.n31 0.189894
R1096 plus.n43 plus.n31 0.189894
R1097 plus.n43 plus.n42 0.189894
R1098 plus.n42 plus.n34 0.189894
R1099 plus.n37 plus.n34 0.189894
R1100 drain_left.n10 drain_left.n8 60.0958
R1101 drain_left.n6 drain_left.n4 60.0956
R1102 drain_left.n2 drain_left.n0 60.0956
R1103 drain_left.n14 drain_left.n13 59.5527
R1104 drain_left.n12 drain_left.n11 59.5527
R1105 drain_left.n10 drain_left.n9 59.5527
R1106 drain_left.n7 drain_left.n3 59.5525
R1107 drain_left.n6 drain_left.n5 59.5525
R1108 drain_left.n2 drain_left.n1 59.5525
R1109 drain_left.n16 drain_left.n15 59.5525
R1110 drain_left drain_left.n7 31.7119
R1111 drain_left drain_left.n16 6.19632
R1112 drain_left.n3 drain_left.t10 1.6505
R1113 drain_left.n3 drain_left.t17 1.6505
R1114 drain_left.n4 drain_left.t13 1.6505
R1115 drain_left.n4 drain_left.t3 1.6505
R1116 drain_left.n5 drain_left.t11 1.6505
R1117 drain_left.n5 drain_left.t2 1.6505
R1118 drain_left.n1 drain_left.t6 1.6505
R1119 drain_left.n1 drain_left.t15 1.6505
R1120 drain_left.n0 drain_left.t5 1.6505
R1121 drain_left.n0 drain_left.t18 1.6505
R1122 drain_left.n15 drain_left.t9 1.6505
R1123 drain_left.n15 drain_left.t4 1.6505
R1124 drain_left.n13 drain_left.t1 1.6505
R1125 drain_left.n13 drain_left.t19 1.6505
R1126 drain_left.n11 drain_left.t14 1.6505
R1127 drain_left.n11 drain_left.t8 1.6505
R1128 drain_left.n9 drain_left.t7 1.6505
R1129 drain_left.n9 drain_left.t0 1.6505
R1130 drain_left.n8 drain_left.t16 1.6505
R1131 drain_left.n8 drain_left.t12 1.6505
R1132 drain_left.n12 drain_left.n10 0.543603
R1133 drain_left.n14 drain_left.n12 0.543603
R1134 drain_left.n16 drain_left.n14 0.543603
R1135 drain_left.n7 drain_left.n6 0.488257
R1136 drain_left.n7 drain_left.n2 0.488257
C0 drain_left minus 0.171748f
C1 source drain_left 37.4577f
C2 plus drain_right 0.36079f
C3 plus minus 5.77444f
C4 minus drain_right 7.17712f
C5 plus source 6.93977f
C6 plus drain_left 7.38307f
C7 source drain_right 37.4581f
C8 source minus 6.92573f
C9 drain_left drain_right 1.10832f
C10 drain_right a_n2102_n3288# 6.94922f
C11 drain_left a_n2102_n3288# 7.268641f
C12 source a_n2102_n3288# 8.808213f
C13 minus a_n2102_n3288# 8.245524f
C14 plus a_n2102_n3288# 10.26762f
C15 drain_left.t5 a_n2102_n3288# 0.324295f
C16 drain_left.t18 a_n2102_n3288# 0.324295f
C17 drain_left.n0 a_n2102_n3288# 2.88952f
C18 drain_left.t6 a_n2102_n3288# 0.324295f
C19 drain_left.t15 a_n2102_n3288# 0.324295f
C20 drain_left.n1 a_n2102_n3288# 2.88572f
C21 drain_left.n2 a_n2102_n3288# 0.818912f
C22 drain_left.t10 a_n2102_n3288# 0.324295f
C23 drain_left.t17 a_n2102_n3288# 0.324295f
C24 drain_left.n3 a_n2102_n3288# 2.88572f
C25 drain_left.t13 a_n2102_n3288# 0.324295f
C26 drain_left.t3 a_n2102_n3288# 0.324295f
C27 drain_left.n4 a_n2102_n3288# 2.88952f
C28 drain_left.t11 a_n2102_n3288# 0.324295f
C29 drain_left.t2 a_n2102_n3288# 0.324295f
C30 drain_left.n5 a_n2102_n3288# 2.88572f
C31 drain_left.n6 a_n2102_n3288# 0.818912f
C32 drain_left.n7 a_n2102_n3288# 2.11674f
C33 drain_left.t16 a_n2102_n3288# 0.324295f
C34 drain_left.t12 a_n2102_n3288# 0.324295f
C35 drain_left.n8 a_n2102_n3288# 2.88953f
C36 drain_left.t7 a_n2102_n3288# 0.324295f
C37 drain_left.t0 a_n2102_n3288# 0.324295f
C38 drain_left.n9 a_n2102_n3288# 2.88573f
C39 drain_left.n10 a_n2102_n3288# 0.823362f
C40 drain_left.t14 a_n2102_n3288# 0.324295f
C41 drain_left.t8 a_n2102_n3288# 0.324295f
C42 drain_left.n11 a_n2102_n3288# 2.88573f
C43 drain_left.n12 a_n2102_n3288# 0.406694f
C44 drain_left.t1 a_n2102_n3288# 0.324295f
C45 drain_left.t19 a_n2102_n3288# 0.324295f
C46 drain_left.n13 a_n2102_n3288# 2.88573f
C47 drain_left.n14 a_n2102_n3288# 0.406694f
C48 drain_left.t9 a_n2102_n3288# 0.324295f
C49 drain_left.t4 a_n2102_n3288# 0.324295f
C50 drain_left.n15 a_n2102_n3288# 2.88572f
C51 drain_left.n16 a_n2102_n3288# 0.691359f
C52 plus.n0 a_n2102_n3288# 0.050217f
C53 plus.t10 a_n2102_n3288# 0.510854f
C54 plus.t0 a_n2102_n3288# 0.510854f
C55 plus.n1 a_n2102_n3288# 0.018361f
C56 plus.n2 a_n2102_n3288# 0.050217f
C57 plus.t11 a_n2102_n3288# 0.510854f
C58 plus.t5 a_n2102_n3288# 0.510854f
C59 plus.t19 a_n2102_n3288# 0.510854f
C60 plus.n3 a_n2102_n3288# 0.202653f
C61 plus.n4 a_n2102_n3288# 0.050217f
C62 plus.t12 a_n2102_n3288# 0.510854f
C63 plus.t7 a_n2102_n3288# 0.510854f
C64 plus.n5 a_n2102_n3288# 0.202653f
C65 plus.t3 a_n2102_n3288# 0.519912f
C66 plus.n6 a_n2102_n3288# 0.218535f
C67 plus.n7 a_n2102_n3288# 0.114909f
C68 plus.n8 a_n2102_n3288# 0.020684f
C69 plus.n9 a_n2102_n3288# 0.202653f
C70 plus.n10 a_n2102_n3288# 0.018981f
C71 plus.n11 a_n2102_n3288# 0.018361f
C72 plus.n12 a_n2102_n3288# 0.050217f
C73 plus.n13 a_n2102_n3288# 0.050217f
C74 plus.n14 a_n2102_n3288# 0.020684f
C75 plus.n15 a_n2102_n3288# 0.202653f
C76 plus.n16 a_n2102_n3288# 0.020684f
C77 plus.n17 a_n2102_n3288# 0.202653f
C78 plus.t18 a_n2102_n3288# 0.510854f
C79 plus.n18 a_n2102_n3288# 0.202653f
C80 plus.n19 a_n2102_n3288# 0.020684f
C81 plus.n20 a_n2102_n3288# 0.050217f
C82 plus.n21 a_n2102_n3288# 0.050217f
C83 plus.n22 a_n2102_n3288# 0.050217f
C84 plus.n23 a_n2102_n3288# 0.018981f
C85 plus.n24 a_n2102_n3288# 0.202653f
C86 plus.n25 a_n2102_n3288# 0.020684f
C87 plus.n26 a_n2102_n3288# 0.202653f
C88 plus.t15 a_n2102_n3288# 0.519912f
C89 plus.n27 a_n2102_n3288# 0.218459f
C90 plus.n28 a_n2102_n3288# 0.563729f
C91 plus.n29 a_n2102_n3288# 0.050217f
C92 plus.t14 a_n2102_n3288# 0.519912f
C93 plus.t1 a_n2102_n3288# 0.510854f
C94 plus.t13 a_n2102_n3288# 0.510854f
C95 plus.n30 a_n2102_n3288# 0.018361f
C96 plus.n31 a_n2102_n3288# 0.050217f
C97 plus.t4 a_n2102_n3288# 0.510854f
C98 plus.n32 a_n2102_n3288# 0.202653f
C99 plus.t9 a_n2102_n3288# 0.510854f
C100 plus.t2 a_n2102_n3288# 0.510854f
C101 plus.t8 a_n2102_n3288# 0.510854f
C102 plus.n33 a_n2102_n3288# 0.202653f
C103 plus.n34 a_n2102_n3288# 0.050217f
C104 plus.t17 a_n2102_n3288# 0.510854f
C105 plus.t6 a_n2102_n3288# 0.510854f
C106 plus.n35 a_n2102_n3288# 0.202653f
C107 plus.t16 a_n2102_n3288# 0.519912f
C108 plus.n36 a_n2102_n3288# 0.218535f
C109 plus.n37 a_n2102_n3288# 0.114909f
C110 plus.n38 a_n2102_n3288# 0.020684f
C111 plus.n39 a_n2102_n3288# 0.202653f
C112 plus.n40 a_n2102_n3288# 0.018981f
C113 plus.n41 a_n2102_n3288# 0.018361f
C114 plus.n42 a_n2102_n3288# 0.050217f
C115 plus.n43 a_n2102_n3288# 0.050217f
C116 plus.n44 a_n2102_n3288# 0.020684f
C117 plus.n45 a_n2102_n3288# 0.202653f
C118 plus.n46 a_n2102_n3288# 0.020684f
C119 plus.n47 a_n2102_n3288# 0.202653f
C120 plus.n48 a_n2102_n3288# 0.020684f
C121 plus.n49 a_n2102_n3288# 0.050217f
C122 plus.n50 a_n2102_n3288# 0.050217f
C123 plus.n51 a_n2102_n3288# 0.050217f
C124 plus.n52 a_n2102_n3288# 0.018981f
C125 plus.n53 a_n2102_n3288# 0.202653f
C126 plus.n54 a_n2102_n3288# 0.020684f
C127 plus.n55 a_n2102_n3288# 0.202653f
C128 plus.n56 a_n2102_n3288# 0.218459f
C129 plus.n57 a_n2102_n3288# 1.56364f
C130 source.n0 a_n2102_n3288# 0.039254f
C131 source.n1 a_n2102_n3288# 0.029634f
C132 source.n2 a_n2102_n3288# 0.015924f
C133 source.n3 a_n2102_n3288# 0.037638f
C134 source.n4 a_n2102_n3288# 0.01686f
C135 source.n5 a_n2102_n3288# 0.029634f
C136 source.n6 a_n2102_n3288# 0.015924f
C137 source.n7 a_n2102_n3288# 0.037638f
C138 source.n8 a_n2102_n3288# 0.01686f
C139 source.n9 a_n2102_n3288# 0.029634f
C140 source.n10 a_n2102_n3288# 0.016392f
C141 source.n11 a_n2102_n3288# 0.037638f
C142 source.n12 a_n2102_n3288# 0.015924f
C143 source.n13 a_n2102_n3288# 0.01686f
C144 source.n14 a_n2102_n3288# 0.029634f
C145 source.n15 a_n2102_n3288# 0.015924f
C146 source.n16 a_n2102_n3288# 0.037638f
C147 source.n17 a_n2102_n3288# 0.01686f
C148 source.n18 a_n2102_n3288# 0.029634f
C149 source.n19 a_n2102_n3288# 0.015924f
C150 source.n20 a_n2102_n3288# 0.028229f
C151 source.n21 a_n2102_n3288# 0.026607f
C152 source.t12 a_n2102_n3288# 0.063568f
C153 source.n22 a_n2102_n3288# 0.213655f
C154 source.n23 a_n2102_n3288# 1.49497f
C155 source.n24 a_n2102_n3288# 0.015924f
C156 source.n25 a_n2102_n3288# 0.01686f
C157 source.n26 a_n2102_n3288# 0.037638f
C158 source.n27 a_n2102_n3288# 0.037638f
C159 source.n28 a_n2102_n3288# 0.01686f
C160 source.n29 a_n2102_n3288# 0.015924f
C161 source.n30 a_n2102_n3288# 0.029634f
C162 source.n31 a_n2102_n3288# 0.029634f
C163 source.n32 a_n2102_n3288# 0.015924f
C164 source.n33 a_n2102_n3288# 0.01686f
C165 source.n34 a_n2102_n3288# 0.037638f
C166 source.n35 a_n2102_n3288# 0.037638f
C167 source.n36 a_n2102_n3288# 0.01686f
C168 source.n37 a_n2102_n3288# 0.015924f
C169 source.n38 a_n2102_n3288# 0.029634f
C170 source.n39 a_n2102_n3288# 0.029634f
C171 source.n40 a_n2102_n3288# 0.015924f
C172 source.n41 a_n2102_n3288# 0.01686f
C173 source.n42 a_n2102_n3288# 0.037638f
C174 source.n43 a_n2102_n3288# 0.037638f
C175 source.n44 a_n2102_n3288# 0.037638f
C176 source.n45 a_n2102_n3288# 0.016392f
C177 source.n46 a_n2102_n3288# 0.015924f
C178 source.n47 a_n2102_n3288# 0.029634f
C179 source.n48 a_n2102_n3288# 0.029634f
C180 source.n49 a_n2102_n3288# 0.015924f
C181 source.n50 a_n2102_n3288# 0.01686f
C182 source.n51 a_n2102_n3288# 0.037638f
C183 source.n52 a_n2102_n3288# 0.037638f
C184 source.n53 a_n2102_n3288# 0.01686f
C185 source.n54 a_n2102_n3288# 0.015924f
C186 source.n55 a_n2102_n3288# 0.029634f
C187 source.n56 a_n2102_n3288# 0.029634f
C188 source.n57 a_n2102_n3288# 0.015924f
C189 source.n58 a_n2102_n3288# 0.01686f
C190 source.n59 a_n2102_n3288# 0.037638f
C191 source.n60 a_n2102_n3288# 0.077238f
C192 source.n61 a_n2102_n3288# 0.01686f
C193 source.n62 a_n2102_n3288# 0.015924f
C194 source.n63 a_n2102_n3288# 0.063639f
C195 source.n64 a_n2102_n3288# 0.042627f
C196 source.n65 a_n2102_n3288# 1.19261f
C197 source.t8 a_n2102_n3288# 0.281009f
C198 source.t0 a_n2102_n3288# 0.281009f
C199 source.n66 a_n2102_n3288# 2.406f
C200 source.n67 a_n2102_n3288# 0.406684f
C201 source.t2 a_n2102_n3288# 0.281009f
C202 source.t7 a_n2102_n3288# 0.281009f
C203 source.n68 a_n2102_n3288# 2.406f
C204 source.n69 a_n2102_n3288# 0.406684f
C205 source.t17 a_n2102_n3288# 0.281009f
C206 source.t14 a_n2102_n3288# 0.281009f
C207 source.n70 a_n2102_n3288# 2.406f
C208 source.n71 a_n2102_n3288# 0.406684f
C209 source.t38 a_n2102_n3288# 0.281009f
C210 source.t16 a_n2102_n3288# 0.281009f
C211 source.n72 a_n2102_n3288# 2.406f
C212 source.n73 a_n2102_n3288# 0.406684f
C213 source.n74 a_n2102_n3288# 0.039254f
C214 source.n75 a_n2102_n3288# 0.029634f
C215 source.n76 a_n2102_n3288# 0.015924f
C216 source.n77 a_n2102_n3288# 0.037638f
C217 source.n78 a_n2102_n3288# 0.01686f
C218 source.n79 a_n2102_n3288# 0.029634f
C219 source.n80 a_n2102_n3288# 0.015924f
C220 source.n81 a_n2102_n3288# 0.037638f
C221 source.n82 a_n2102_n3288# 0.01686f
C222 source.n83 a_n2102_n3288# 0.029634f
C223 source.n84 a_n2102_n3288# 0.016392f
C224 source.n85 a_n2102_n3288# 0.037638f
C225 source.n86 a_n2102_n3288# 0.015924f
C226 source.n87 a_n2102_n3288# 0.01686f
C227 source.n88 a_n2102_n3288# 0.029634f
C228 source.n89 a_n2102_n3288# 0.015924f
C229 source.n90 a_n2102_n3288# 0.037638f
C230 source.n91 a_n2102_n3288# 0.01686f
C231 source.n92 a_n2102_n3288# 0.029634f
C232 source.n93 a_n2102_n3288# 0.015924f
C233 source.n94 a_n2102_n3288# 0.028229f
C234 source.n95 a_n2102_n3288# 0.026607f
C235 source.t11 a_n2102_n3288# 0.063568f
C236 source.n96 a_n2102_n3288# 0.213655f
C237 source.n97 a_n2102_n3288# 1.49497f
C238 source.n98 a_n2102_n3288# 0.015924f
C239 source.n99 a_n2102_n3288# 0.01686f
C240 source.n100 a_n2102_n3288# 0.037638f
C241 source.n101 a_n2102_n3288# 0.037638f
C242 source.n102 a_n2102_n3288# 0.01686f
C243 source.n103 a_n2102_n3288# 0.015924f
C244 source.n104 a_n2102_n3288# 0.029634f
C245 source.n105 a_n2102_n3288# 0.029634f
C246 source.n106 a_n2102_n3288# 0.015924f
C247 source.n107 a_n2102_n3288# 0.01686f
C248 source.n108 a_n2102_n3288# 0.037638f
C249 source.n109 a_n2102_n3288# 0.037638f
C250 source.n110 a_n2102_n3288# 0.01686f
C251 source.n111 a_n2102_n3288# 0.015924f
C252 source.n112 a_n2102_n3288# 0.029634f
C253 source.n113 a_n2102_n3288# 0.029634f
C254 source.n114 a_n2102_n3288# 0.015924f
C255 source.n115 a_n2102_n3288# 0.01686f
C256 source.n116 a_n2102_n3288# 0.037638f
C257 source.n117 a_n2102_n3288# 0.037638f
C258 source.n118 a_n2102_n3288# 0.037638f
C259 source.n119 a_n2102_n3288# 0.016392f
C260 source.n120 a_n2102_n3288# 0.015924f
C261 source.n121 a_n2102_n3288# 0.029634f
C262 source.n122 a_n2102_n3288# 0.029634f
C263 source.n123 a_n2102_n3288# 0.015924f
C264 source.n124 a_n2102_n3288# 0.01686f
C265 source.n125 a_n2102_n3288# 0.037638f
C266 source.n126 a_n2102_n3288# 0.037638f
C267 source.n127 a_n2102_n3288# 0.01686f
C268 source.n128 a_n2102_n3288# 0.015924f
C269 source.n129 a_n2102_n3288# 0.029634f
C270 source.n130 a_n2102_n3288# 0.029634f
C271 source.n131 a_n2102_n3288# 0.015924f
C272 source.n132 a_n2102_n3288# 0.01686f
C273 source.n133 a_n2102_n3288# 0.037638f
C274 source.n134 a_n2102_n3288# 0.077238f
C275 source.n135 a_n2102_n3288# 0.01686f
C276 source.n136 a_n2102_n3288# 0.015924f
C277 source.n137 a_n2102_n3288# 0.063639f
C278 source.n138 a_n2102_n3288# 0.042627f
C279 source.n139 a_n2102_n3288# 0.119294f
C280 source.n140 a_n2102_n3288# 0.039254f
C281 source.n141 a_n2102_n3288# 0.029634f
C282 source.n142 a_n2102_n3288# 0.015924f
C283 source.n143 a_n2102_n3288# 0.037638f
C284 source.n144 a_n2102_n3288# 0.01686f
C285 source.n145 a_n2102_n3288# 0.029634f
C286 source.n146 a_n2102_n3288# 0.015924f
C287 source.n147 a_n2102_n3288# 0.037638f
C288 source.n148 a_n2102_n3288# 0.01686f
C289 source.n149 a_n2102_n3288# 0.029634f
C290 source.n150 a_n2102_n3288# 0.016392f
C291 source.n151 a_n2102_n3288# 0.037638f
C292 source.n152 a_n2102_n3288# 0.015924f
C293 source.n153 a_n2102_n3288# 0.01686f
C294 source.n154 a_n2102_n3288# 0.029634f
C295 source.n155 a_n2102_n3288# 0.015924f
C296 source.n156 a_n2102_n3288# 0.037638f
C297 source.n157 a_n2102_n3288# 0.01686f
C298 source.n158 a_n2102_n3288# 0.029634f
C299 source.n159 a_n2102_n3288# 0.015924f
C300 source.n160 a_n2102_n3288# 0.028229f
C301 source.n161 a_n2102_n3288# 0.026607f
C302 source.t26 a_n2102_n3288# 0.063568f
C303 source.n162 a_n2102_n3288# 0.213655f
C304 source.n163 a_n2102_n3288# 1.49497f
C305 source.n164 a_n2102_n3288# 0.015924f
C306 source.n165 a_n2102_n3288# 0.01686f
C307 source.n166 a_n2102_n3288# 0.037638f
C308 source.n167 a_n2102_n3288# 0.037638f
C309 source.n168 a_n2102_n3288# 0.01686f
C310 source.n169 a_n2102_n3288# 0.015924f
C311 source.n170 a_n2102_n3288# 0.029634f
C312 source.n171 a_n2102_n3288# 0.029634f
C313 source.n172 a_n2102_n3288# 0.015924f
C314 source.n173 a_n2102_n3288# 0.01686f
C315 source.n174 a_n2102_n3288# 0.037638f
C316 source.n175 a_n2102_n3288# 0.037638f
C317 source.n176 a_n2102_n3288# 0.01686f
C318 source.n177 a_n2102_n3288# 0.015924f
C319 source.n178 a_n2102_n3288# 0.029634f
C320 source.n179 a_n2102_n3288# 0.029634f
C321 source.n180 a_n2102_n3288# 0.015924f
C322 source.n181 a_n2102_n3288# 0.01686f
C323 source.n182 a_n2102_n3288# 0.037638f
C324 source.n183 a_n2102_n3288# 0.037638f
C325 source.n184 a_n2102_n3288# 0.037638f
C326 source.n185 a_n2102_n3288# 0.016392f
C327 source.n186 a_n2102_n3288# 0.015924f
C328 source.n187 a_n2102_n3288# 0.029634f
C329 source.n188 a_n2102_n3288# 0.029634f
C330 source.n189 a_n2102_n3288# 0.015924f
C331 source.n190 a_n2102_n3288# 0.01686f
C332 source.n191 a_n2102_n3288# 0.037638f
C333 source.n192 a_n2102_n3288# 0.037638f
C334 source.n193 a_n2102_n3288# 0.01686f
C335 source.n194 a_n2102_n3288# 0.015924f
C336 source.n195 a_n2102_n3288# 0.029634f
C337 source.n196 a_n2102_n3288# 0.029634f
C338 source.n197 a_n2102_n3288# 0.015924f
C339 source.n198 a_n2102_n3288# 0.01686f
C340 source.n199 a_n2102_n3288# 0.037638f
C341 source.n200 a_n2102_n3288# 0.077238f
C342 source.n201 a_n2102_n3288# 0.01686f
C343 source.n202 a_n2102_n3288# 0.015924f
C344 source.n203 a_n2102_n3288# 0.063639f
C345 source.n204 a_n2102_n3288# 0.042627f
C346 source.n205 a_n2102_n3288# 0.119294f
C347 source.t33 a_n2102_n3288# 0.281009f
C348 source.t19 a_n2102_n3288# 0.281009f
C349 source.n206 a_n2102_n3288# 2.406f
C350 source.n207 a_n2102_n3288# 0.406684f
C351 source.t20 a_n2102_n3288# 0.281009f
C352 source.t27 a_n2102_n3288# 0.281009f
C353 source.n208 a_n2102_n3288# 2.406f
C354 source.n209 a_n2102_n3288# 0.406684f
C355 source.t31 a_n2102_n3288# 0.281009f
C356 source.t35 a_n2102_n3288# 0.281009f
C357 source.n210 a_n2102_n3288# 2.406f
C358 source.n211 a_n2102_n3288# 0.406684f
C359 source.t32 a_n2102_n3288# 0.281009f
C360 source.t18 a_n2102_n3288# 0.281009f
C361 source.n212 a_n2102_n3288# 2.406f
C362 source.n213 a_n2102_n3288# 0.406684f
C363 source.n214 a_n2102_n3288# 0.039254f
C364 source.n215 a_n2102_n3288# 0.029634f
C365 source.n216 a_n2102_n3288# 0.015924f
C366 source.n217 a_n2102_n3288# 0.037638f
C367 source.n218 a_n2102_n3288# 0.01686f
C368 source.n219 a_n2102_n3288# 0.029634f
C369 source.n220 a_n2102_n3288# 0.015924f
C370 source.n221 a_n2102_n3288# 0.037638f
C371 source.n222 a_n2102_n3288# 0.01686f
C372 source.n223 a_n2102_n3288# 0.029634f
C373 source.n224 a_n2102_n3288# 0.016392f
C374 source.n225 a_n2102_n3288# 0.037638f
C375 source.n226 a_n2102_n3288# 0.015924f
C376 source.n227 a_n2102_n3288# 0.01686f
C377 source.n228 a_n2102_n3288# 0.029634f
C378 source.n229 a_n2102_n3288# 0.015924f
C379 source.n230 a_n2102_n3288# 0.037638f
C380 source.n231 a_n2102_n3288# 0.01686f
C381 source.n232 a_n2102_n3288# 0.029634f
C382 source.n233 a_n2102_n3288# 0.015924f
C383 source.n234 a_n2102_n3288# 0.028229f
C384 source.n235 a_n2102_n3288# 0.026607f
C385 source.t30 a_n2102_n3288# 0.063568f
C386 source.n236 a_n2102_n3288# 0.213655f
C387 source.n237 a_n2102_n3288# 1.49497f
C388 source.n238 a_n2102_n3288# 0.015924f
C389 source.n239 a_n2102_n3288# 0.01686f
C390 source.n240 a_n2102_n3288# 0.037638f
C391 source.n241 a_n2102_n3288# 0.037638f
C392 source.n242 a_n2102_n3288# 0.01686f
C393 source.n243 a_n2102_n3288# 0.015924f
C394 source.n244 a_n2102_n3288# 0.029634f
C395 source.n245 a_n2102_n3288# 0.029634f
C396 source.n246 a_n2102_n3288# 0.015924f
C397 source.n247 a_n2102_n3288# 0.01686f
C398 source.n248 a_n2102_n3288# 0.037638f
C399 source.n249 a_n2102_n3288# 0.037638f
C400 source.n250 a_n2102_n3288# 0.01686f
C401 source.n251 a_n2102_n3288# 0.015924f
C402 source.n252 a_n2102_n3288# 0.029634f
C403 source.n253 a_n2102_n3288# 0.029634f
C404 source.n254 a_n2102_n3288# 0.015924f
C405 source.n255 a_n2102_n3288# 0.01686f
C406 source.n256 a_n2102_n3288# 0.037638f
C407 source.n257 a_n2102_n3288# 0.037638f
C408 source.n258 a_n2102_n3288# 0.037638f
C409 source.n259 a_n2102_n3288# 0.016392f
C410 source.n260 a_n2102_n3288# 0.015924f
C411 source.n261 a_n2102_n3288# 0.029634f
C412 source.n262 a_n2102_n3288# 0.029634f
C413 source.n263 a_n2102_n3288# 0.015924f
C414 source.n264 a_n2102_n3288# 0.01686f
C415 source.n265 a_n2102_n3288# 0.037638f
C416 source.n266 a_n2102_n3288# 0.037638f
C417 source.n267 a_n2102_n3288# 0.01686f
C418 source.n268 a_n2102_n3288# 0.015924f
C419 source.n269 a_n2102_n3288# 0.029634f
C420 source.n270 a_n2102_n3288# 0.029634f
C421 source.n271 a_n2102_n3288# 0.015924f
C422 source.n272 a_n2102_n3288# 0.01686f
C423 source.n273 a_n2102_n3288# 0.037638f
C424 source.n274 a_n2102_n3288# 0.077238f
C425 source.n275 a_n2102_n3288# 0.01686f
C426 source.n276 a_n2102_n3288# 0.015924f
C427 source.n277 a_n2102_n3288# 0.063639f
C428 source.n278 a_n2102_n3288# 0.042627f
C429 source.n279 a_n2102_n3288# 1.65857f
C430 source.n280 a_n2102_n3288# 0.039254f
C431 source.n281 a_n2102_n3288# 0.029634f
C432 source.n282 a_n2102_n3288# 0.015924f
C433 source.n283 a_n2102_n3288# 0.037638f
C434 source.n284 a_n2102_n3288# 0.01686f
C435 source.n285 a_n2102_n3288# 0.029634f
C436 source.n286 a_n2102_n3288# 0.015924f
C437 source.n287 a_n2102_n3288# 0.037638f
C438 source.n288 a_n2102_n3288# 0.01686f
C439 source.n289 a_n2102_n3288# 0.029634f
C440 source.n290 a_n2102_n3288# 0.016392f
C441 source.n291 a_n2102_n3288# 0.037638f
C442 source.n292 a_n2102_n3288# 0.01686f
C443 source.n293 a_n2102_n3288# 0.029634f
C444 source.n294 a_n2102_n3288# 0.015924f
C445 source.n295 a_n2102_n3288# 0.037638f
C446 source.n296 a_n2102_n3288# 0.01686f
C447 source.n297 a_n2102_n3288# 0.029634f
C448 source.n298 a_n2102_n3288# 0.015924f
C449 source.n299 a_n2102_n3288# 0.028229f
C450 source.n300 a_n2102_n3288# 0.026607f
C451 source.t6 a_n2102_n3288# 0.063568f
C452 source.n301 a_n2102_n3288# 0.213655f
C453 source.n302 a_n2102_n3288# 1.49497f
C454 source.n303 a_n2102_n3288# 0.015924f
C455 source.n304 a_n2102_n3288# 0.01686f
C456 source.n305 a_n2102_n3288# 0.037638f
C457 source.n306 a_n2102_n3288# 0.037638f
C458 source.n307 a_n2102_n3288# 0.01686f
C459 source.n308 a_n2102_n3288# 0.015924f
C460 source.n309 a_n2102_n3288# 0.029634f
C461 source.n310 a_n2102_n3288# 0.029634f
C462 source.n311 a_n2102_n3288# 0.015924f
C463 source.n312 a_n2102_n3288# 0.01686f
C464 source.n313 a_n2102_n3288# 0.037638f
C465 source.n314 a_n2102_n3288# 0.037638f
C466 source.n315 a_n2102_n3288# 0.01686f
C467 source.n316 a_n2102_n3288# 0.015924f
C468 source.n317 a_n2102_n3288# 0.029634f
C469 source.n318 a_n2102_n3288# 0.029634f
C470 source.n319 a_n2102_n3288# 0.015924f
C471 source.n320 a_n2102_n3288# 0.015924f
C472 source.n321 a_n2102_n3288# 0.01686f
C473 source.n322 a_n2102_n3288# 0.037638f
C474 source.n323 a_n2102_n3288# 0.037638f
C475 source.n324 a_n2102_n3288# 0.037638f
C476 source.n325 a_n2102_n3288# 0.016392f
C477 source.n326 a_n2102_n3288# 0.015924f
C478 source.n327 a_n2102_n3288# 0.029634f
C479 source.n328 a_n2102_n3288# 0.029634f
C480 source.n329 a_n2102_n3288# 0.015924f
C481 source.n330 a_n2102_n3288# 0.01686f
C482 source.n331 a_n2102_n3288# 0.037638f
C483 source.n332 a_n2102_n3288# 0.037638f
C484 source.n333 a_n2102_n3288# 0.01686f
C485 source.n334 a_n2102_n3288# 0.015924f
C486 source.n335 a_n2102_n3288# 0.029634f
C487 source.n336 a_n2102_n3288# 0.029634f
C488 source.n337 a_n2102_n3288# 0.015924f
C489 source.n338 a_n2102_n3288# 0.01686f
C490 source.n339 a_n2102_n3288# 0.037638f
C491 source.n340 a_n2102_n3288# 0.077238f
C492 source.n341 a_n2102_n3288# 0.01686f
C493 source.n342 a_n2102_n3288# 0.015924f
C494 source.n343 a_n2102_n3288# 0.063639f
C495 source.n344 a_n2102_n3288# 0.042627f
C496 source.n345 a_n2102_n3288# 1.65857f
C497 source.t1 a_n2102_n3288# 0.281009f
C498 source.t10 a_n2102_n3288# 0.281009f
C499 source.n346 a_n2102_n3288# 2.40599f
C500 source.n347 a_n2102_n3288# 0.406699f
C501 source.t13 a_n2102_n3288# 0.281009f
C502 source.t3 a_n2102_n3288# 0.281009f
C503 source.n348 a_n2102_n3288# 2.40599f
C504 source.n349 a_n2102_n3288# 0.406699f
C505 source.t4 a_n2102_n3288# 0.281009f
C506 source.t39 a_n2102_n3288# 0.281009f
C507 source.n350 a_n2102_n3288# 2.40599f
C508 source.n351 a_n2102_n3288# 0.406699f
C509 source.t5 a_n2102_n3288# 0.281009f
C510 source.t9 a_n2102_n3288# 0.281009f
C511 source.n352 a_n2102_n3288# 2.40599f
C512 source.n353 a_n2102_n3288# 0.406699f
C513 source.n354 a_n2102_n3288# 0.039254f
C514 source.n355 a_n2102_n3288# 0.029634f
C515 source.n356 a_n2102_n3288# 0.015924f
C516 source.n357 a_n2102_n3288# 0.037638f
C517 source.n358 a_n2102_n3288# 0.01686f
C518 source.n359 a_n2102_n3288# 0.029634f
C519 source.n360 a_n2102_n3288# 0.015924f
C520 source.n361 a_n2102_n3288# 0.037638f
C521 source.n362 a_n2102_n3288# 0.01686f
C522 source.n363 a_n2102_n3288# 0.029634f
C523 source.n364 a_n2102_n3288# 0.016392f
C524 source.n365 a_n2102_n3288# 0.037638f
C525 source.n366 a_n2102_n3288# 0.01686f
C526 source.n367 a_n2102_n3288# 0.029634f
C527 source.n368 a_n2102_n3288# 0.015924f
C528 source.n369 a_n2102_n3288# 0.037638f
C529 source.n370 a_n2102_n3288# 0.01686f
C530 source.n371 a_n2102_n3288# 0.029634f
C531 source.n372 a_n2102_n3288# 0.015924f
C532 source.n373 a_n2102_n3288# 0.028229f
C533 source.n374 a_n2102_n3288# 0.026607f
C534 source.t15 a_n2102_n3288# 0.063568f
C535 source.n375 a_n2102_n3288# 0.213655f
C536 source.n376 a_n2102_n3288# 1.49497f
C537 source.n377 a_n2102_n3288# 0.015924f
C538 source.n378 a_n2102_n3288# 0.01686f
C539 source.n379 a_n2102_n3288# 0.037638f
C540 source.n380 a_n2102_n3288# 0.037638f
C541 source.n381 a_n2102_n3288# 0.01686f
C542 source.n382 a_n2102_n3288# 0.015924f
C543 source.n383 a_n2102_n3288# 0.029634f
C544 source.n384 a_n2102_n3288# 0.029634f
C545 source.n385 a_n2102_n3288# 0.015924f
C546 source.n386 a_n2102_n3288# 0.01686f
C547 source.n387 a_n2102_n3288# 0.037638f
C548 source.n388 a_n2102_n3288# 0.037638f
C549 source.n389 a_n2102_n3288# 0.01686f
C550 source.n390 a_n2102_n3288# 0.015924f
C551 source.n391 a_n2102_n3288# 0.029634f
C552 source.n392 a_n2102_n3288# 0.029634f
C553 source.n393 a_n2102_n3288# 0.015924f
C554 source.n394 a_n2102_n3288# 0.015924f
C555 source.n395 a_n2102_n3288# 0.01686f
C556 source.n396 a_n2102_n3288# 0.037638f
C557 source.n397 a_n2102_n3288# 0.037638f
C558 source.n398 a_n2102_n3288# 0.037638f
C559 source.n399 a_n2102_n3288# 0.016392f
C560 source.n400 a_n2102_n3288# 0.015924f
C561 source.n401 a_n2102_n3288# 0.029634f
C562 source.n402 a_n2102_n3288# 0.029634f
C563 source.n403 a_n2102_n3288# 0.015924f
C564 source.n404 a_n2102_n3288# 0.01686f
C565 source.n405 a_n2102_n3288# 0.037638f
C566 source.n406 a_n2102_n3288# 0.037638f
C567 source.n407 a_n2102_n3288# 0.01686f
C568 source.n408 a_n2102_n3288# 0.015924f
C569 source.n409 a_n2102_n3288# 0.029634f
C570 source.n410 a_n2102_n3288# 0.029634f
C571 source.n411 a_n2102_n3288# 0.015924f
C572 source.n412 a_n2102_n3288# 0.01686f
C573 source.n413 a_n2102_n3288# 0.037638f
C574 source.n414 a_n2102_n3288# 0.077238f
C575 source.n415 a_n2102_n3288# 0.01686f
C576 source.n416 a_n2102_n3288# 0.015924f
C577 source.n417 a_n2102_n3288# 0.063639f
C578 source.n418 a_n2102_n3288# 0.042627f
C579 source.n419 a_n2102_n3288# 0.119294f
C580 source.n420 a_n2102_n3288# 0.039254f
C581 source.n421 a_n2102_n3288# 0.029634f
C582 source.n422 a_n2102_n3288# 0.015924f
C583 source.n423 a_n2102_n3288# 0.037638f
C584 source.n424 a_n2102_n3288# 0.01686f
C585 source.n425 a_n2102_n3288# 0.029634f
C586 source.n426 a_n2102_n3288# 0.015924f
C587 source.n427 a_n2102_n3288# 0.037638f
C588 source.n428 a_n2102_n3288# 0.01686f
C589 source.n429 a_n2102_n3288# 0.029634f
C590 source.n430 a_n2102_n3288# 0.016392f
C591 source.n431 a_n2102_n3288# 0.037638f
C592 source.n432 a_n2102_n3288# 0.01686f
C593 source.n433 a_n2102_n3288# 0.029634f
C594 source.n434 a_n2102_n3288# 0.015924f
C595 source.n435 a_n2102_n3288# 0.037638f
C596 source.n436 a_n2102_n3288# 0.01686f
C597 source.n437 a_n2102_n3288# 0.029634f
C598 source.n438 a_n2102_n3288# 0.015924f
C599 source.n439 a_n2102_n3288# 0.028229f
C600 source.n440 a_n2102_n3288# 0.026607f
C601 source.t36 a_n2102_n3288# 0.063568f
C602 source.n441 a_n2102_n3288# 0.213655f
C603 source.n442 a_n2102_n3288# 1.49497f
C604 source.n443 a_n2102_n3288# 0.015924f
C605 source.n444 a_n2102_n3288# 0.01686f
C606 source.n445 a_n2102_n3288# 0.037638f
C607 source.n446 a_n2102_n3288# 0.037638f
C608 source.n447 a_n2102_n3288# 0.01686f
C609 source.n448 a_n2102_n3288# 0.015924f
C610 source.n449 a_n2102_n3288# 0.029634f
C611 source.n450 a_n2102_n3288# 0.029634f
C612 source.n451 a_n2102_n3288# 0.015924f
C613 source.n452 a_n2102_n3288# 0.01686f
C614 source.n453 a_n2102_n3288# 0.037638f
C615 source.n454 a_n2102_n3288# 0.037638f
C616 source.n455 a_n2102_n3288# 0.01686f
C617 source.n456 a_n2102_n3288# 0.015924f
C618 source.n457 a_n2102_n3288# 0.029634f
C619 source.n458 a_n2102_n3288# 0.029634f
C620 source.n459 a_n2102_n3288# 0.015924f
C621 source.n460 a_n2102_n3288# 0.015924f
C622 source.n461 a_n2102_n3288# 0.01686f
C623 source.n462 a_n2102_n3288# 0.037638f
C624 source.n463 a_n2102_n3288# 0.037638f
C625 source.n464 a_n2102_n3288# 0.037638f
C626 source.n465 a_n2102_n3288# 0.016392f
C627 source.n466 a_n2102_n3288# 0.015924f
C628 source.n467 a_n2102_n3288# 0.029634f
C629 source.n468 a_n2102_n3288# 0.029634f
C630 source.n469 a_n2102_n3288# 0.015924f
C631 source.n470 a_n2102_n3288# 0.01686f
C632 source.n471 a_n2102_n3288# 0.037638f
C633 source.n472 a_n2102_n3288# 0.037638f
C634 source.n473 a_n2102_n3288# 0.01686f
C635 source.n474 a_n2102_n3288# 0.015924f
C636 source.n475 a_n2102_n3288# 0.029634f
C637 source.n476 a_n2102_n3288# 0.029634f
C638 source.n477 a_n2102_n3288# 0.015924f
C639 source.n478 a_n2102_n3288# 0.01686f
C640 source.n479 a_n2102_n3288# 0.037638f
C641 source.n480 a_n2102_n3288# 0.077238f
C642 source.n481 a_n2102_n3288# 0.01686f
C643 source.n482 a_n2102_n3288# 0.015924f
C644 source.n483 a_n2102_n3288# 0.063639f
C645 source.n484 a_n2102_n3288# 0.042627f
C646 source.n485 a_n2102_n3288# 0.119294f
C647 source.t24 a_n2102_n3288# 0.281009f
C648 source.t37 a_n2102_n3288# 0.281009f
C649 source.n486 a_n2102_n3288# 2.40599f
C650 source.n487 a_n2102_n3288# 0.406699f
C651 source.t25 a_n2102_n3288# 0.281009f
C652 source.t28 a_n2102_n3288# 0.281009f
C653 source.n488 a_n2102_n3288# 2.40599f
C654 source.n489 a_n2102_n3288# 0.406699f
C655 source.t21 a_n2102_n3288# 0.281009f
C656 source.t29 a_n2102_n3288# 0.281009f
C657 source.n490 a_n2102_n3288# 2.40599f
C658 source.n491 a_n2102_n3288# 0.406699f
C659 source.t22 a_n2102_n3288# 0.281009f
C660 source.t23 a_n2102_n3288# 0.281009f
C661 source.n492 a_n2102_n3288# 2.40599f
C662 source.n493 a_n2102_n3288# 0.406699f
C663 source.n494 a_n2102_n3288# 0.039254f
C664 source.n495 a_n2102_n3288# 0.029634f
C665 source.n496 a_n2102_n3288# 0.015924f
C666 source.n497 a_n2102_n3288# 0.037638f
C667 source.n498 a_n2102_n3288# 0.01686f
C668 source.n499 a_n2102_n3288# 0.029634f
C669 source.n500 a_n2102_n3288# 0.015924f
C670 source.n501 a_n2102_n3288# 0.037638f
C671 source.n502 a_n2102_n3288# 0.01686f
C672 source.n503 a_n2102_n3288# 0.029634f
C673 source.n504 a_n2102_n3288# 0.016392f
C674 source.n505 a_n2102_n3288# 0.037638f
C675 source.n506 a_n2102_n3288# 0.01686f
C676 source.n507 a_n2102_n3288# 0.029634f
C677 source.n508 a_n2102_n3288# 0.015924f
C678 source.n509 a_n2102_n3288# 0.037638f
C679 source.n510 a_n2102_n3288# 0.01686f
C680 source.n511 a_n2102_n3288# 0.029634f
C681 source.n512 a_n2102_n3288# 0.015924f
C682 source.n513 a_n2102_n3288# 0.028229f
C683 source.n514 a_n2102_n3288# 0.026607f
C684 source.t34 a_n2102_n3288# 0.063568f
C685 source.n515 a_n2102_n3288# 0.213655f
C686 source.n516 a_n2102_n3288# 1.49497f
C687 source.n517 a_n2102_n3288# 0.015924f
C688 source.n518 a_n2102_n3288# 0.01686f
C689 source.n519 a_n2102_n3288# 0.037638f
C690 source.n520 a_n2102_n3288# 0.037638f
C691 source.n521 a_n2102_n3288# 0.01686f
C692 source.n522 a_n2102_n3288# 0.015924f
C693 source.n523 a_n2102_n3288# 0.029634f
C694 source.n524 a_n2102_n3288# 0.029634f
C695 source.n525 a_n2102_n3288# 0.015924f
C696 source.n526 a_n2102_n3288# 0.01686f
C697 source.n527 a_n2102_n3288# 0.037638f
C698 source.n528 a_n2102_n3288# 0.037638f
C699 source.n529 a_n2102_n3288# 0.01686f
C700 source.n530 a_n2102_n3288# 0.015924f
C701 source.n531 a_n2102_n3288# 0.029634f
C702 source.n532 a_n2102_n3288# 0.029634f
C703 source.n533 a_n2102_n3288# 0.015924f
C704 source.n534 a_n2102_n3288# 0.015924f
C705 source.n535 a_n2102_n3288# 0.01686f
C706 source.n536 a_n2102_n3288# 0.037638f
C707 source.n537 a_n2102_n3288# 0.037638f
C708 source.n538 a_n2102_n3288# 0.037638f
C709 source.n539 a_n2102_n3288# 0.016392f
C710 source.n540 a_n2102_n3288# 0.015924f
C711 source.n541 a_n2102_n3288# 0.029634f
C712 source.n542 a_n2102_n3288# 0.029634f
C713 source.n543 a_n2102_n3288# 0.015924f
C714 source.n544 a_n2102_n3288# 0.01686f
C715 source.n545 a_n2102_n3288# 0.037638f
C716 source.n546 a_n2102_n3288# 0.037638f
C717 source.n547 a_n2102_n3288# 0.01686f
C718 source.n548 a_n2102_n3288# 0.015924f
C719 source.n549 a_n2102_n3288# 0.029634f
C720 source.n550 a_n2102_n3288# 0.029634f
C721 source.n551 a_n2102_n3288# 0.015924f
C722 source.n552 a_n2102_n3288# 0.01686f
C723 source.n553 a_n2102_n3288# 0.037638f
C724 source.n554 a_n2102_n3288# 0.077238f
C725 source.n555 a_n2102_n3288# 0.01686f
C726 source.n556 a_n2102_n3288# 0.015924f
C727 source.n557 a_n2102_n3288# 0.063639f
C728 source.n558 a_n2102_n3288# 0.042627f
C729 source.n559 a_n2102_n3288# 0.286576f
C730 source.n560 a_n2102_n3288# 1.85904f
C731 drain_right.t11 a_n2102_n3288# 0.323815f
C732 drain_right.t4 a_n2102_n3288# 0.323815f
C733 drain_right.n0 a_n2102_n3288# 2.88525f
C734 drain_right.t10 a_n2102_n3288# 0.323815f
C735 drain_right.t8 a_n2102_n3288# 0.323815f
C736 drain_right.n1 a_n2102_n3288# 2.88145f
C737 drain_right.n2 a_n2102_n3288# 0.817701f
C738 drain_right.t14 a_n2102_n3288# 0.323815f
C739 drain_right.t7 a_n2102_n3288# 0.323815f
C740 drain_right.n3 a_n2102_n3288# 2.88145f
C741 drain_right.t1 a_n2102_n3288# 0.323815f
C742 drain_right.t13 a_n2102_n3288# 0.323815f
C743 drain_right.n4 a_n2102_n3288# 2.88525f
C744 drain_right.t15 a_n2102_n3288# 0.323815f
C745 drain_right.t2 a_n2102_n3288# 0.323815f
C746 drain_right.n5 a_n2102_n3288# 2.88145f
C747 drain_right.n6 a_n2102_n3288# 0.817701f
C748 drain_right.n7 a_n2102_n3288# 2.04311f
C749 drain_right.t17 a_n2102_n3288# 0.323815f
C750 drain_right.t18 a_n2102_n3288# 0.323815f
C751 drain_right.n8 a_n2102_n3288# 2.88525f
C752 drain_right.t5 a_n2102_n3288# 0.323815f
C753 drain_right.t12 a_n2102_n3288# 0.323815f
C754 drain_right.n9 a_n2102_n3288# 2.88146f
C755 drain_right.n10 a_n2102_n3288# 0.822156f
C756 drain_right.t9 a_n2102_n3288# 0.323815f
C757 drain_right.t0 a_n2102_n3288# 0.323815f
C758 drain_right.n11 a_n2102_n3288# 2.88146f
C759 drain_right.n12 a_n2102_n3288# 0.406092f
C760 drain_right.t6 a_n2102_n3288# 0.323815f
C761 drain_right.t16 a_n2102_n3288# 0.323815f
C762 drain_right.n13 a_n2102_n3288# 2.88146f
C763 drain_right.n14 a_n2102_n3288# 0.406092f
C764 drain_right.t3 a_n2102_n3288# 0.323815f
C765 drain_right.t19 a_n2102_n3288# 0.323815f
C766 drain_right.n15 a_n2102_n3288# 2.88146f
C767 drain_right.n16 a_n2102_n3288# 0.690325f
C768 minus.n0 a_n2102_n3288# 0.049467f
C769 minus.t7 a_n2102_n3288# 0.512151f
C770 minus.t5 a_n2102_n3288# 0.503229f
C771 minus.t19 a_n2102_n3288# 0.503229f
C772 minus.n1 a_n2102_n3288# 0.018087f
C773 minus.n2 a_n2102_n3288# 0.049467f
C774 minus.t6 a_n2102_n3288# 0.503229f
C775 minus.n3 a_n2102_n3288# 0.199628f
C776 minus.t2 a_n2102_n3288# 0.503229f
C777 minus.t17 a_n2102_n3288# 0.503229f
C778 minus.t10 a_n2102_n3288# 0.503229f
C779 minus.n4 a_n2102_n3288# 0.199628f
C780 minus.n5 a_n2102_n3288# 0.049467f
C781 minus.t4 a_n2102_n3288# 0.503229f
C782 minus.t18 a_n2102_n3288# 0.503229f
C783 minus.n6 a_n2102_n3288# 0.199628f
C784 minus.t11 a_n2102_n3288# 0.512151f
C785 minus.n7 a_n2102_n3288# 0.215273f
C786 minus.n8 a_n2102_n3288# 0.113194f
C787 minus.n9 a_n2102_n3288# 0.020375f
C788 minus.n10 a_n2102_n3288# 0.199628f
C789 minus.n11 a_n2102_n3288# 0.018697f
C790 minus.n12 a_n2102_n3288# 0.018087f
C791 minus.n13 a_n2102_n3288# 0.049467f
C792 minus.n14 a_n2102_n3288# 0.049467f
C793 minus.n15 a_n2102_n3288# 0.020375f
C794 minus.n16 a_n2102_n3288# 0.199628f
C795 minus.n17 a_n2102_n3288# 0.020375f
C796 minus.n18 a_n2102_n3288# 0.199628f
C797 minus.n19 a_n2102_n3288# 0.020375f
C798 minus.n20 a_n2102_n3288# 0.049467f
C799 minus.n21 a_n2102_n3288# 0.049467f
C800 minus.n22 a_n2102_n3288# 0.049467f
C801 minus.n23 a_n2102_n3288# 0.018697f
C802 minus.n24 a_n2102_n3288# 0.199628f
C803 minus.n25 a_n2102_n3288# 0.020375f
C804 minus.n26 a_n2102_n3288# 0.199628f
C805 minus.n27 a_n2102_n3288# 0.215198f
C806 minus.n28 a_n2102_n3288# 1.81728f
C807 minus.n29 a_n2102_n3288# 0.049467f
C808 minus.t14 a_n2102_n3288# 0.503229f
C809 minus.t15 a_n2102_n3288# 0.503229f
C810 minus.n30 a_n2102_n3288# 0.018087f
C811 minus.n31 a_n2102_n3288# 0.049467f
C812 minus.t16 a_n2102_n3288# 0.503229f
C813 minus.t9 a_n2102_n3288# 0.503229f
C814 minus.t12 a_n2102_n3288# 0.503229f
C815 minus.n32 a_n2102_n3288# 0.199628f
C816 minus.n33 a_n2102_n3288# 0.049467f
C817 minus.t0 a_n2102_n3288# 0.503229f
C818 minus.t13 a_n2102_n3288# 0.503229f
C819 minus.n34 a_n2102_n3288# 0.199628f
C820 minus.t1 a_n2102_n3288# 0.512151f
C821 minus.n35 a_n2102_n3288# 0.215273f
C822 minus.n36 a_n2102_n3288# 0.113194f
C823 minus.n37 a_n2102_n3288# 0.020375f
C824 minus.n38 a_n2102_n3288# 0.199628f
C825 minus.n39 a_n2102_n3288# 0.018697f
C826 minus.n40 a_n2102_n3288# 0.018087f
C827 minus.n41 a_n2102_n3288# 0.049467f
C828 minus.n42 a_n2102_n3288# 0.049467f
C829 minus.n43 a_n2102_n3288# 0.020375f
C830 minus.n44 a_n2102_n3288# 0.199628f
C831 minus.n45 a_n2102_n3288# 0.020375f
C832 minus.n46 a_n2102_n3288# 0.199628f
C833 minus.t8 a_n2102_n3288# 0.503229f
C834 minus.n47 a_n2102_n3288# 0.199628f
C835 minus.n48 a_n2102_n3288# 0.020375f
C836 minus.n49 a_n2102_n3288# 0.049467f
C837 minus.n50 a_n2102_n3288# 0.049467f
C838 minus.n51 a_n2102_n3288# 0.049467f
C839 minus.n52 a_n2102_n3288# 0.018697f
C840 minus.n53 a_n2102_n3288# 0.199628f
C841 minus.n54 a_n2102_n3288# 0.020375f
C842 minus.n55 a_n2102_n3288# 0.199628f
C843 minus.t3 a_n2102_n3288# 0.512151f
C844 minus.n56 a_n2102_n3288# 0.215198f
C845 minus.n57 a_n2102_n3288# 0.325227f
C846 minus.n58 a_n2102_n3288# 2.20101f
.ends

