* NGSPICE file created from diffpair399.ext - technology: sky130A

.subckt diffpair399 minus drain_right drain_left source plus
X0 drain_right.t23 minus.t0 source.t43 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X1 a_n3654_n2688# a_n3654_n2688# a_n3654_n2688# a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.8
X2 drain_right.t22 minus.t1 source.t27 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X3 source.t2 plus.t0 drain_left.t23 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X4 source.t35 minus.t2 drain_right.t21 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X5 drain_left.t22 plus.t1 source.t12 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X6 source.t0 plus.t2 drain_left.t21 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X7 drain_left.t20 plus.t3 source.t11 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X8 drain_right.t20 minus.t3 source.t39 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X9 drain_left.t19 plus.t4 source.t5 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X10 source.t32 minus.t4 drain_right.t19 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X11 drain_left.t18 plus.t5 source.t8 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X12 source.t3 plus.t6 drain_left.t17 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X13 drain_right.t18 minus.t5 source.t31 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X14 drain_left.t16 plus.t7 source.t45 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X15 drain_left.t15 plus.t8 source.t1 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X16 drain_left.t14 plus.t9 source.t46 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X17 source.t29 minus.t6 drain_right.t17 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X18 source.t41 minus.t7 drain_right.t16 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X19 source.t33 minus.t8 drain_right.t15 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X20 drain_right.t14 minus.t9 source.t26 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X21 drain_right.t13 minus.t10 source.t44 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X22 source.t28 minus.t11 drain_right.t12 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X23 drain_right.t11 minus.t12 source.t36 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X24 source.t40 minus.t13 drain_right.t10 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X25 source.t47 plus.t10 drain_left.t13 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X26 source.t34 minus.t14 drain_right.t9 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X27 source.t13 plus.t11 drain_left.t12 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X28 drain_left.t11 plus.t12 source.t4 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X29 source.t30 minus.t15 drain_right.t8 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X30 drain_right.t7 minus.t16 source.t42 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X31 drain_left.t10 plus.t13 source.t14 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X32 drain_right.t6 minus.t17 source.t23 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X33 drain_right.t5 minus.t18 source.t25 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.8
X34 source.t20 plus.t14 drain_left.t9 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X35 a_n3654_n2688# a_n3654_n2688# a_n3654_n2688# a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X36 source.t24 minus.t19 drain_right.t4 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X37 drain_left.t8 plus.t15 source.t17 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X38 drain_left.t7 plus.t16 source.t7 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X39 source.t22 minus.t20 drain_right.t3 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X40 source.t37 minus.t21 drain_right.t2 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X41 source.t15 plus.t17 drain_left.t6 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X42 source.t18 plus.t18 drain_left.t5 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X43 source.t10 plus.t19 drain_left.t4 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X44 drain_right.t1 minus.t22 source.t21 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X45 source.t19 plus.t20 drain_left.t3 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X46 drain_left.t2 plus.t21 source.t9 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X47 a_n3654_n2688# a_n3654_n2688# a_n3654_n2688# a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X48 drain_right.t0 minus.t23 source.t38 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
X49 a_n3654_n2688# a_n3654_n2688# a_n3654_n2688# a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.8
X50 source.t16 plus.t22 drain_left.t1 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.8
X51 source.t6 plus.t23 drain_left.t0 a_n3654_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.8
R0 minus.n8 minus.t12 341.666
R1 minus.n44 minus.t21 341.666
R2 minus.n9 minus.t6 320.229
R3 minus.n10 minus.t5 320.229
R4 minus.n14 minus.t15 320.229
R5 minus.n16 minus.t17 320.229
R6 minus.n20 minus.t14 320.229
R7 minus.n21 minus.t9 320.229
R8 minus.n3 minus.t20 320.229
R9 minus.n27 minus.t16 320.229
R10 minus.n1 minus.t4 320.229
R11 minus.n32 minus.t10 320.229
R12 minus.n34 minus.t7 320.229
R13 minus.n45 minus.t3 320.229
R14 minus.n46 minus.t11 320.229
R15 minus.n50 minus.t1 320.229
R16 minus.n52 minus.t19 320.229
R17 minus.n56 minus.t0 320.229
R18 minus.n57 minus.t8 320.229
R19 minus.n39 minus.t22 320.229
R20 minus.n63 minus.t13 320.229
R21 minus.n37 minus.t23 320.229
R22 minus.n68 minus.t2 320.229
R23 minus.n70 minus.t18 320.229
R24 minus.n35 minus.n34 161.3
R25 minus.n33 minus.n0 161.3
R26 minus.n29 minus.n28 161.3
R27 minus.n27 minus.n2 161.3
R28 minus.n26 minus.n25 161.3
R29 minus.n24 minus.n3 161.3
R30 minus.n23 minus.n22 161.3
R31 minus.n18 minus.n5 161.3
R32 minus.n17 minus.n16 161.3
R33 minus.n15 minus.n6 161.3
R34 minus.n14 minus.n13 161.3
R35 minus.n12 minus.n7 161.3
R36 minus.n71 minus.n70 161.3
R37 minus.n69 minus.n36 161.3
R38 minus.n65 minus.n64 161.3
R39 minus.n63 minus.n38 161.3
R40 minus.n62 minus.n61 161.3
R41 minus.n60 minus.n39 161.3
R42 minus.n59 minus.n58 161.3
R43 minus.n54 minus.n41 161.3
R44 minus.n53 minus.n52 161.3
R45 minus.n51 minus.n42 161.3
R46 minus.n50 minus.n49 161.3
R47 minus.n48 minus.n43 161.3
R48 minus.n32 minus.n31 80.6037
R49 minus.n30 minus.n1 80.6037
R50 minus.n21 minus.n4 80.6037
R51 minus.n20 minus.n19 80.6037
R52 minus.n11 minus.n10 80.6037
R53 minus.n68 minus.n67 80.6037
R54 minus.n66 minus.n37 80.6037
R55 minus.n57 minus.n40 80.6037
R56 minus.n56 minus.n55 80.6037
R57 minus.n47 minus.n46 80.6037
R58 minus.n10 minus.n9 48.2005
R59 minus.n21 minus.n20 48.2005
R60 minus.n32 minus.n1 48.2005
R61 minus.n46 minus.n45 48.2005
R62 minus.n57 minus.n56 48.2005
R63 minus.n68 minus.n37 48.2005
R64 minus.n10 minus.n7 44.549
R65 minus.n28 minus.n1 44.549
R66 minus.n46 minus.n43 44.549
R67 minus.n64 minus.n37 44.549
R68 minus.n20 minus.n5 41.6278
R69 minus.n22 minus.n21 41.6278
R70 minus.n56 minus.n41 41.6278
R71 minus.n58 minus.n57 41.6278
R72 minus.n72 minus.n35 40.849
R73 minus.n33 minus.n32 38.7066
R74 minus.n69 minus.n68 38.7066
R75 minus.n11 minus.n8 31.6825
R76 minus.n47 minus.n44 31.6825
R77 minus.n15 minus.n14 25.5611
R78 minus.n27 minus.n26 25.5611
R79 minus.n51 minus.n50 25.5611
R80 minus.n63 minus.n62 25.5611
R81 minus.n16 minus.n15 22.6399
R82 minus.n26 minus.n3 22.6399
R83 minus.n52 minus.n51 22.6399
R84 minus.n62 minus.n39 22.6399
R85 minus.n9 minus.n8 17.2341
R86 minus.n45 minus.n44 17.2341
R87 minus.n34 minus.n33 9.49444
R88 minus.n70 minus.n69 9.49444
R89 minus.n72 minus.n71 6.65959
R90 minus.n16 minus.n5 6.57323
R91 minus.n22 minus.n3 6.57323
R92 minus.n52 minus.n41 6.57323
R93 minus.n58 minus.n39 6.57323
R94 minus.n14 minus.n7 3.65202
R95 minus.n28 minus.n27 3.65202
R96 minus.n50 minus.n43 3.65202
R97 minus.n64 minus.n63 3.65202
R98 minus.n31 minus.n30 0.380177
R99 minus.n19 minus.n4 0.380177
R100 minus.n55 minus.n40 0.380177
R101 minus.n67 minus.n66 0.380177
R102 minus.n31 minus.n0 0.285035
R103 minus.n30 minus.n29 0.285035
R104 minus.n23 minus.n4 0.285035
R105 minus.n19 minus.n18 0.285035
R106 minus.n12 minus.n11 0.285035
R107 minus.n48 minus.n47 0.285035
R108 minus.n55 minus.n54 0.285035
R109 minus.n59 minus.n40 0.285035
R110 minus.n66 minus.n65 0.285035
R111 minus.n67 minus.n36 0.285035
R112 minus.n35 minus.n0 0.189894
R113 minus.n29 minus.n2 0.189894
R114 minus.n25 minus.n2 0.189894
R115 minus.n25 minus.n24 0.189894
R116 minus.n24 minus.n23 0.189894
R117 minus.n18 minus.n17 0.189894
R118 minus.n17 minus.n6 0.189894
R119 minus.n13 minus.n6 0.189894
R120 minus.n13 minus.n12 0.189894
R121 minus.n49 minus.n48 0.189894
R122 minus.n49 minus.n42 0.189894
R123 minus.n53 minus.n42 0.189894
R124 minus.n54 minus.n53 0.189894
R125 minus.n60 minus.n59 0.189894
R126 minus.n61 minus.n60 0.189894
R127 minus.n61 minus.n38 0.189894
R128 minus.n65 minus.n38 0.189894
R129 minus.n71 minus.n36 0.189894
R130 minus minus.n72 0.188
R131 source.n11 source.t16 51.0588
R132 source.n12 source.t36 51.0588
R133 source.n23 source.t41 51.0588
R134 source.n47 source.t25 51.0586
R135 source.n36 source.t37 51.0586
R136 source.n35 source.t14 51.0586
R137 source.n24 source.t10 51.0586
R138 source.n0 source.t8 51.0586
R139 source.n2 source.n1 48.8588
R140 source.n4 source.n3 48.8588
R141 source.n6 source.n5 48.8588
R142 source.n8 source.n7 48.8588
R143 source.n10 source.n9 48.8588
R144 source.n14 source.n13 48.8588
R145 source.n16 source.n15 48.8588
R146 source.n18 source.n17 48.8588
R147 source.n20 source.n19 48.8588
R148 source.n22 source.n21 48.8588
R149 source.n46 source.n45 48.8586
R150 source.n44 source.n43 48.8586
R151 source.n42 source.n41 48.8586
R152 source.n40 source.n39 48.8586
R153 source.n38 source.n37 48.8586
R154 source.n34 source.n33 48.8586
R155 source.n32 source.n31 48.8586
R156 source.n30 source.n29 48.8586
R157 source.n28 source.n27 48.8586
R158 source.n26 source.n25 48.8586
R159 source.n24 source.n23 19.9891
R160 source.n48 source.n0 14.2391
R161 source.n48 source.n47 5.7505
R162 source.n45 source.t38 2.2005
R163 source.n45 source.t35 2.2005
R164 source.n43 source.t21 2.2005
R165 source.n43 source.t40 2.2005
R166 source.n41 source.t43 2.2005
R167 source.n41 source.t33 2.2005
R168 source.n39 source.t27 2.2005
R169 source.n39 source.t24 2.2005
R170 source.n37 source.t39 2.2005
R171 source.n37 source.t28 2.2005
R172 source.n33 source.t1 2.2005
R173 source.n33 source.t0 2.2005
R174 source.n31 source.t45 2.2005
R175 source.n31 source.t2 2.2005
R176 source.n29 source.t5 2.2005
R177 source.n29 source.t15 2.2005
R178 source.n27 source.t12 2.2005
R179 source.n27 source.t6 2.2005
R180 source.n25 source.t11 2.2005
R181 source.n25 source.t13 2.2005
R182 source.n1 source.t46 2.2005
R183 source.n1 source.t3 2.2005
R184 source.n3 source.t4 2.2005
R185 source.n3 source.t47 2.2005
R186 source.n5 source.t17 2.2005
R187 source.n5 source.t20 2.2005
R188 source.n7 source.t7 2.2005
R189 source.n7 source.t19 2.2005
R190 source.n9 source.t9 2.2005
R191 source.n9 source.t18 2.2005
R192 source.n13 source.t31 2.2005
R193 source.n13 source.t29 2.2005
R194 source.n15 source.t23 2.2005
R195 source.n15 source.t30 2.2005
R196 source.n17 source.t26 2.2005
R197 source.n17 source.t34 2.2005
R198 source.n19 source.t42 2.2005
R199 source.n19 source.t22 2.2005
R200 source.n21 source.t44 2.2005
R201 source.n21 source.t32 2.2005
R202 source.n23 source.n22 0.974638
R203 source.n22 source.n20 0.974638
R204 source.n20 source.n18 0.974638
R205 source.n18 source.n16 0.974638
R206 source.n16 source.n14 0.974638
R207 source.n14 source.n12 0.974638
R208 source.n11 source.n10 0.974638
R209 source.n10 source.n8 0.974638
R210 source.n8 source.n6 0.974638
R211 source.n6 source.n4 0.974638
R212 source.n4 source.n2 0.974638
R213 source.n2 source.n0 0.974638
R214 source.n26 source.n24 0.974638
R215 source.n28 source.n26 0.974638
R216 source.n30 source.n28 0.974638
R217 source.n32 source.n30 0.974638
R218 source.n34 source.n32 0.974638
R219 source.n35 source.n34 0.974638
R220 source.n38 source.n36 0.974638
R221 source.n40 source.n38 0.974638
R222 source.n42 source.n40 0.974638
R223 source.n44 source.n42 0.974638
R224 source.n46 source.n44 0.974638
R225 source.n47 source.n46 0.974638
R226 source.n12 source.n11 0.470328
R227 source.n36 source.n35 0.470328
R228 source source.n48 0.188
R229 drain_right.n13 drain_right.n11 66.5116
R230 drain_right.n7 drain_right.n5 66.5115
R231 drain_right.n2 drain_right.n0 66.5115
R232 drain_right.n13 drain_right.n12 65.5376
R233 drain_right.n15 drain_right.n14 65.5376
R234 drain_right.n17 drain_right.n16 65.5376
R235 drain_right.n19 drain_right.n18 65.5376
R236 drain_right.n21 drain_right.n20 65.5376
R237 drain_right.n7 drain_right.n6 65.5373
R238 drain_right.n9 drain_right.n8 65.5373
R239 drain_right.n4 drain_right.n3 65.5373
R240 drain_right.n2 drain_right.n1 65.5373
R241 drain_right drain_right.n10 33.7954
R242 drain_right drain_right.n21 6.62735
R243 drain_right.n5 drain_right.t21 2.2005
R244 drain_right.n5 drain_right.t5 2.2005
R245 drain_right.n6 drain_right.t10 2.2005
R246 drain_right.n6 drain_right.t0 2.2005
R247 drain_right.n8 drain_right.t15 2.2005
R248 drain_right.n8 drain_right.t1 2.2005
R249 drain_right.n3 drain_right.t4 2.2005
R250 drain_right.n3 drain_right.t23 2.2005
R251 drain_right.n1 drain_right.t12 2.2005
R252 drain_right.n1 drain_right.t22 2.2005
R253 drain_right.n0 drain_right.t2 2.2005
R254 drain_right.n0 drain_right.t20 2.2005
R255 drain_right.n11 drain_right.t17 2.2005
R256 drain_right.n11 drain_right.t11 2.2005
R257 drain_right.n12 drain_right.t8 2.2005
R258 drain_right.n12 drain_right.t18 2.2005
R259 drain_right.n14 drain_right.t9 2.2005
R260 drain_right.n14 drain_right.t6 2.2005
R261 drain_right.n16 drain_right.t3 2.2005
R262 drain_right.n16 drain_right.t14 2.2005
R263 drain_right.n18 drain_right.t19 2.2005
R264 drain_right.n18 drain_right.t7 2.2005
R265 drain_right.n20 drain_right.t16 2.2005
R266 drain_right.n20 drain_right.t13 2.2005
R267 drain_right.n9 drain_right.n7 0.974638
R268 drain_right.n4 drain_right.n2 0.974638
R269 drain_right.n21 drain_right.n19 0.974638
R270 drain_right.n19 drain_right.n17 0.974638
R271 drain_right.n17 drain_right.n15 0.974638
R272 drain_right.n15 drain_right.n13 0.974638
R273 drain_right.n10 drain_right.n9 0.432223
R274 drain_right.n10 drain_right.n4 0.432223
R275 plus.n10 plus.t22 341.666
R276 plus.n46 plus.t13 341.666
R277 plus.n34 plus.t5 320.229
R278 plus.n32 plus.t6 320.229
R279 plus.n31 plus.t9 320.229
R280 plus.n3 plus.t10 320.229
R281 plus.n25 plus.t12 320.229
R282 plus.n5 plus.t14 320.229
R283 plus.n20 plus.t15 320.229
R284 plus.n18 plus.t20 320.229
R285 plus.n8 plus.t16 320.229
R286 plus.n12 plus.t18 320.229
R287 plus.n11 plus.t21 320.229
R288 plus.n70 plus.t19 320.229
R289 plus.n68 plus.t3 320.229
R290 plus.n67 plus.t11 320.229
R291 plus.n39 plus.t1 320.229
R292 plus.n61 plus.t23 320.229
R293 plus.n41 plus.t4 320.229
R294 plus.n56 plus.t17 320.229
R295 plus.n54 plus.t7 320.229
R296 plus.n44 plus.t0 320.229
R297 plus.n48 plus.t8 320.229
R298 plus.n47 plus.t2 320.229
R299 plus.n14 plus.n13 161.3
R300 plus.n15 plus.n8 161.3
R301 plus.n17 plus.n16 161.3
R302 plus.n18 plus.n7 161.3
R303 plus.n19 plus.n6 161.3
R304 plus.n24 plus.n23 161.3
R305 plus.n25 plus.n4 161.3
R306 plus.n27 plus.n26 161.3
R307 plus.n28 plus.n3 161.3
R308 plus.n30 plus.n29 161.3
R309 plus.n33 plus.n0 161.3
R310 plus.n35 plus.n34 161.3
R311 plus.n50 plus.n49 161.3
R312 plus.n51 plus.n44 161.3
R313 plus.n53 plus.n52 161.3
R314 plus.n54 plus.n43 161.3
R315 plus.n55 plus.n42 161.3
R316 plus.n60 plus.n59 161.3
R317 plus.n61 plus.n40 161.3
R318 plus.n63 plus.n62 161.3
R319 plus.n64 plus.n39 161.3
R320 plus.n66 plus.n65 161.3
R321 plus.n69 plus.n36 161.3
R322 plus.n71 plus.n70 161.3
R323 plus.n12 plus.n9 80.6037
R324 plus.n21 plus.n20 80.6037
R325 plus.n22 plus.n5 80.6037
R326 plus.n31 plus.n2 80.6037
R327 plus.n32 plus.n1 80.6037
R328 plus.n48 plus.n45 80.6037
R329 plus.n57 plus.n56 80.6037
R330 plus.n58 plus.n41 80.6037
R331 plus.n67 plus.n38 80.6037
R332 plus.n68 plus.n37 80.6037
R333 plus.n32 plus.n31 48.2005
R334 plus.n20 plus.n5 48.2005
R335 plus.n12 plus.n11 48.2005
R336 plus.n68 plus.n67 48.2005
R337 plus.n56 plus.n41 48.2005
R338 plus.n48 plus.n47 48.2005
R339 plus.n31 plus.n30 44.549
R340 plus.n13 plus.n12 44.549
R341 plus.n67 plus.n66 44.549
R342 plus.n49 plus.n48 44.549
R343 plus.n24 plus.n5 41.6278
R344 plus.n20 plus.n19 41.6278
R345 plus.n60 plus.n41 41.6278
R346 plus.n56 plus.n55 41.6278
R347 plus.n33 plus.n32 38.7066
R348 plus.n69 plus.n68 38.7066
R349 plus plus.n71 35.8664
R350 plus.n10 plus.n9 31.6825
R351 plus.n46 plus.n45 31.6825
R352 plus.n26 plus.n3 25.5611
R353 plus.n17 plus.n8 25.5611
R354 plus.n62 plus.n39 25.5611
R355 plus.n53 plus.n44 25.5611
R356 plus.n26 plus.n25 22.6399
R357 plus.n18 plus.n17 22.6399
R358 plus.n62 plus.n61 22.6399
R359 plus.n54 plus.n53 22.6399
R360 plus.n11 plus.n10 17.2341
R361 plus.n47 plus.n46 17.2341
R362 plus plus.n35 11.1672
R363 plus.n34 plus.n33 9.49444
R364 plus.n70 plus.n69 9.49444
R365 plus.n25 plus.n24 6.57323
R366 plus.n19 plus.n18 6.57323
R367 plus.n61 plus.n60 6.57323
R368 plus.n55 plus.n54 6.57323
R369 plus.n30 plus.n3 3.65202
R370 plus.n13 plus.n8 3.65202
R371 plus.n66 plus.n39 3.65202
R372 plus.n49 plus.n44 3.65202
R373 plus.n22 plus.n21 0.380177
R374 plus.n2 plus.n1 0.380177
R375 plus.n38 plus.n37 0.380177
R376 plus.n58 plus.n57 0.380177
R377 plus.n14 plus.n9 0.285035
R378 plus.n21 plus.n6 0.285035
R379 plus.n23 plus.n22 0.285035
R380 plus.n29 plus.n2 0.285035
R381 plus.n1 plus.n0 0.285035
R382 plus.n37 plus.n36 0.285035
R383 plus.n65 plus.n38 0.285035
R384 plus.n59 plus.n58 0.285035
R385 plus.n57 plus.n42 0.285035
R386 plus.n50 plus.n45 0.285035
R387 plus.n15 plus.n14 0.189894
R388 plus.n16 plus.n15 0.189894
R389 plus.n16 plus.n7 0.189894
R390 plus.n7 plus.n6 0.189894
R391 plus.n23 plus.n4 0.189894
R392 plus.n27 plus.n4 0.189894
R393 plus.n28 plus.n27 0.189894
R394 plus.n29 plus.n28 0.189894
R395 plus.n35 plus.n0 0.189894
R396 plus.n71 plus.n36 0.189894
R397 plus.n65 plus.n64 0.189894
R398 plus.n64 plus.n63 0.189894
R399 plus.n63 plus.n40 0.189894
R400 plus.n59 plus.n40 0.189894
R401 plus.n43 plus.n42 0.189894
R402 plus.n52 plus.n43 0.189894
R403 plus.n52 plus.n51 0.189894
R404 plus.n51 plus.n50 0.189894
R405 drain_left.n13 drain_left.n11 66.5117
R406 drain_left.n7 drain_left.n5 66.5115
R407 drain_left.n2 drain_left.n0 66.5115
R408 drain_left.n19 drain_left.n18 65.5376
R409 drain_left.n17 drain_left.n16 65.5376
R410 drain_left.n15 drain_left.n14 65.5376
R411 drain_left.n13 drain_left.n12 65.5376
R412 drain_left.n21 drain_left.n20 65.5374
R413 drain_left.n7 drain_left.n6 65.5373
R414 drain_left.n9 drain_left.n8 65.5373
R415 drain_left.n4 drain_left.n3 65.5373
R416 drain_left.n2 drain_left.n1 65.5373
R417 drain_left drain_left.n10 34.3487
R418 drain_left drain_left.n21 6.62735
R419 drain_left.n5 drain_left.t21 2.2005
R420 drain_left.n5 drain_left.t10 2.2005
R421 drain_left.n6 drain_left.t23 2.2005
R422 drain_left.n6 drain_left.t15 2.2005
R423 drain_left.n8 drain_left.t6 2.2005
R424 drain_left.n8 drain_left.t16 2.2005
R425 drain_left.n3 drain_left.t0 2.2005
R426 drain_left.n3 drain_left.t19 2.2005
R427 drain_left.n1 drain_left.t12 2.2005
R428 drain_left.n1 drain_left.t22 2.2005
R429 drain_left.n0 drain_left.t4 2.2005
R430 drain_left.n0 drain_left.t20 2.2005
R431 drain_left.n20 drain_left.t17 2.2005
R432 drain_left.n20 drain_left.t18 2.2005
R433 drain_left.n18 drain_left.t13 2.2005
R434 drain_left.n18 drain_left.t14 2.2005
R435 drain_left.n16 drain_left.t9 2.2005
R436 drain_left.n16 drain_left.t11 2.2005
R437 drain_left.n14 drain_left.t3 2.2005
R438 drain_left.n14 drain_left.t8 2.2005
R439 drain_left.n12 drain_left.t5 2.2005
R440 drain_left.n12 drain_left.t7 2.2005
R441 drain_left.n11 drain_left.t1 2.2005
R442 drain_left.n11 drain_left.t2 2.2005
R443 drain_left.n9 drain_left.n7 0.974638
R444 drain_left.n4 drain_left.n2 0.974638
R445 drain_left.n15 drain_left.n13 0.974638
R446 drain_left.n17 drain_left.n15 0.974638
R447 drain_left.n19 drain_left.n17 0.974638
R448 drain_left.n21 drain_left.n19 0.974638
R449 drain_left.n10 drain_left.n9 0.432223
R450 drain_left.n10 drain_left.n4 0.432223
C0 drain_left plus 12.617599f
C1 drain_left minus 0.175388f
C2 drain_right source 21.1063f
C3 minus plus 7.15324f
C4 drain_left source 21.103199f
C5 source plus 12.7847f
C6 drain_left drain_right 2.02887f
C7 minus source 12.7707f
C8 drain_right plus 0.526806f
C9 drain_right minus 12.250099f
C10 drain_right a_n3654_n2688# 7.74371f
C11 drain_left a_n3654_n2688# 8.24617f
C12 source a_n3654_n2688# 8.058252f
C13 minus a_n3654_n2688# 14.672474f
C14 plus a_n3654_n2688# 16.38678f
C15 drain_left.t4 a_n3654_n2688# 0.200995f
C16 drain_left.t20 a_n3654_n2688# 0.200995f
C17 drain_left.n0 a_n3654_n2688# 1.76412f
C18 drain_left.t12 a_n3654_n2688# 0.200995f
C19 drain_left.t22 a_n3654_n2688# 0.200995f
C20 drain_left.n1 a_n3654_n2688# 1.75804f
C21 drain_left.n2 a_n3654_n2688# 0.812886f
C22 drain_left.t0 a_n3654_n2688# 0.200995f
C23 drain_left.t19 a_n3654_n2688# 0.200995f
C24 drain_left.n3 a_n3654_n2688# 1.75804f
C25 drain_left.n4 a_n3654_n2688# 0.355915f
C26 drain_left.t21 a_n3654_n2688# 0.200995f
C27 drain_left.t10 a_n3654_n2688# 0.200995f
C28 drain_left.n5 a_n3654_n2688# 1.76412f
C29 drain_left.t23 a_n3654_n2688# 0.200995f
C30 drain_left.t15 a_n3654_n2688# 0.200995f
C31 drain_left.n6 a_n3654_n2688# 1.75804f
C32 drain_left.n7 a_n3654_n2688# 0.812886f
C33 drain_left.t6 a_n3654_n2688# 0.200995f
C34 drain_left.t16 a_n3654_n2688# 0.200995f
C35 drain_left.n8 a_n3654_n2688# 1.75804f
C36 drain_left.n9 a_n3654_n2688# 0.355915f
C37 drain_left.n10 a_n3654_n2688# 1.75399f
C38 drain_left.t1 a_n3654_n2688# 0.200995f
C39 drain_left.t2 a_n3654_n2688# 0.200995f
C40 drain_left.n11 a_n3654_n2688# 1.76412f
C41 drain_left.t5 a_n3654_n2688# 0.200995f
C42 drain_left.t7 a_n3654_n2688# 0.200995f
C43 drain_left.n12 a_n3654_n2688# 1.75804f
C44 drain_left.n13 a_n3654_n2688# 0.812879f
C45 drain_left.t3 a_n3654_n2688# 0.200995f
C46 drain_left.t8 a_n3654_n2688# 0.200995f
C47 drain_left.n14 a_n3654_n2688# 1.75804f
C48 drain_left.n15 a_n3654_n2688# 0.403788f
C49 drain_left.t9 a_n3654_n2688# 0.200995f
C50 drain_left.t11 a_n3654_n2688# 0.200995f
C51 drain_left.n16 a_n3654_n2688# 1.75804f
C52 drain_left.n17 a_n3654_n2688# 0.403788f
C53 drain_left.t13 a_n3654_n2688# 0.200995f
C54 drain_left.t14 a_n3654_n2688# 0.200995f
C55 drain_left.n18 a_n3654_n2688# 1.75804f
C56 drain_left.n19 a_n3654_n2688# 0.403788f
C57 drain_left.t17 a_n3654_n2688# 0.200995f
C58 drain_left.t18 a_n3654_n2688# 0.200995f
C59 drain_left.n20 a_n3654_n2688# 1.75803f
C60 drain_left.n21 a_n3654_n2688# 0.657212f
C61 plus.n0 a_n3654_n2688# 0.050722f
C62 plus.t5 a_n3654_n2688# 0.784885f
C63 plus.t6 a_n3654_n2688# 0.784885f
C64 plus.n1 a_n3654_n2688# 0.063313f
C65 plus.t9 a_n3654_n2688# 0.784885f
C66 plus.n2 a_n3654_n2688# 0.063313f
C67 plus.t10 a_n3654_n2688# 0.784885f
C68 plus.n3 a_n3654_n2688# 0.326294f
C69 plus.n4 a_n3654_n2688# 0.038012f
C70 plus.t12 a_n3654_n2688# 0.784885f
C71 plus.t14 a_n3654_n2688# 0.784885f
C72 plus.n5 a_n3654_n2688# 0.336912f
C73 plus.n6 a_n3654_n2688# 0.050722f
C74 plus.t15 a_n3654_n2688# 0.784885f
C75 plus.t20 a_n3654_n2688# 0.784885f
C76 plus.n7 a_n3654_n2688# 0.038012f
C77 plus.t16 a_n3654_n2688# 0.784885f
C78 plus.n8 a_n3654_n2688# 0.326294f
C79 plus.n9 a_n3654_n2688# 0.218476f
C80 plus.t18 a_n3654_n2688# 0.784885f
C81 plus.t21 a_n3654_n2688# 0.784885f
C82 plus.t22 a_n3654_n2688# 0.805558f
C83 plus.n10 a_n3654_n2688# 0.312438f
C84 plus.n11 a_n3654_n2688# 0.337361f
C85 plus.n12 a_n3654_n2688# 0.33738f
C86 plus.n13 a_n3654_n2688# 0.008626f
C87 plus.n14 a_n3654_n2688# 0.050722f
C88 plus.n15 a_n3654_n2688# 0.038012f
C89 plus.n16 a_n3654_n2688# 0.038012f
C90 plus.n17 a_n3654_n2688# 0.008626f
C91 plus.n18 a_n3654_n2688# 0.326294f
C92 plus.n19 a_n3654_n2688# 0.008626f
C93 plus.n20 a_n3654_n2688# 0.336912f
C94 plus.n21 a_n3654_n2688# 0.063313f
C95 plus.n22 a_n3654_n2688# 0.063313f
C96 plus.n23 a_n3654_n2688# 0.050722f
C97 plus.n24 a_n3654_n2688# 0.008626f
C98 plus.n25 a_n3654_n2688# 0.326294f
C99 plus.n26 a_n3654_n2688# 0.008626f
C100 plus.n27 a_n3654_n2688# 0.038012f
C101 plus.n28 a_n3654_n2688# 0.038012f
C102 plus.n29 a_n3654_n2688# 0.050722f
C103 plus.n30 a_n3654_n2688# 0.008626f
C104 plus.n31 a_n3654_n2688# 0.33738f
C105 plus.n32 a_n3654_n2688# 0.336443f
C106 plus.n33 a_n3654_n2688# 0.008626f
C107 plus.n34 a_n3654_n2688# 0.32313f
C108 plus.n35 a_n3654_n2688# 0.388033f
C109 plus.n36 a_n3654_n2688# 0.050722f
C110 plus.t19 a_n3654_n2688# 0.784885f
C111 plus.n37 a_n3654_n2688# 0.063313f
C112 plus.t3 a_n3654_n2688# 0.784885f
C113 plus.n38 a_n3654_n2688# 0.063313f
C114 plus.t11 a_n3654_n2688# 0.784885f
C115 plus.t1 a_n3654_n2688# 0.784885f
C116 plus.n39 a_n3654_n2688# 0.326294f
C117 plus.n40 a_n3654_n2688# 0.038012f
C118 plus.t23 a_n3654_n2688# 0.784885f
C119 plus.t4 a_n3654_n2688# 0.784885f
C120 plus.n41 a_n3654_n2688# 0.336912f
C121 plus.n42 a_n3654_n2688# 0.050722f
C122 plus.t17 a_n3654_n2688# 0.784885f
C123 plus.n43 a_n3654_n2688# 0.038012f
C124 plus.t7 a_n3654_n2688# 0.784885f
C125 plus.t0 a_n3654_n2688# 0.784885f
C126 plus.n44 a_n3654_n2688# 0.326294f
C127 plus.n45 a_n3654_n2688# 0.218476f
C128 plus.t8 a_n3654_n2688# 0.784885f
C129 plus.t13 a_n3654_n2688# 0.805558f
C130 plus.n46 a_n3654_n2688# 0.312438f
C131 plus.t2 a_n3654_n2688# 0.784885f
C132 plus.n47 a_n3654_n2688# 0.337361f
C133 plus.n48 a_n3654_n2688# 0.33738f
C134 plus.n49 a_n3654_n2688# 0.008626f
C135 plus.n50 a_n3654_n2688# 0.050722f
C136 plus.n51 a_n3654_n2688# 0.038012f
C137 plus.n52 a_n3654_n2688# 0.038012f
C138 plus.n53 a_n3654_n2688# 0.008626f
C139 plus.n54 a_n3654_n2688# 0.326294f
C140 plus.n55 a_n3654_n2688# 0.008626f
C141 plus.n56 a_n3654_n2688# 0.336912f
C142 plus.n57 a_n3654_n2688# 0.063313f
C143 plus.n58 a_n3654_n2688# 0.063313f
C144 plus.n59 a_n3654_n2688# 0.050722f
C145 plus.n60 a_n3654_n2688# 0.008626f
C146 plus.n61 a_n3654_n2688# 0.326294f
C147 plus.n62 a_n3654_n2688# 0.008626f
C148 plus.n63 a_n3654_n2688# 0.038012f
C149 plus.n64 a_n3654_n2688# 0.038012f
C150 plus.n65 a_n3654_n2688# 0.050722f
C151 plus.n66 a_n3654_n2688# 0.008626f
C152 plus.n67 a_n3654_n2688# 0.33738f
C153 plus.n68 a_n3654_n2688# 0.336443f
C154 plus.n69 a_n3654_n2688# 0.008626f
C155 plus.n70 a_n3654_n2688# 0.32313f
C156 plus.n71 a_n3654_n2688# 1.43226f
C157 drain_right.t2 a_n3654_n2688# 0.199925f
C158 drain_right.t20 a_n3654_n2688# 0.199925f
C159 drain_right.n0 a_n3654_n2688# 1.75473f
C160 drain_right.t12 a_n3654_n2688# 0.199925f
C161 drain_right.t22 a_n3654_n2688# 0.199925f
C162 drain_right.n1 a_n3654_n2688# 1.74868f
C163 drain_right.n2 a_n3654_n2688# 0.808559f
C164 drain_right.t4 a_n3654_n2688# 0.199925f
C165 drain_right.t23 a_n3654_n2688# 0.199925f
C166 drain_right.n3 a_n3654_n2688# 1.74868f
C167 drain_right.n4 a_n3654_n2688# 0.354021f
C168 drain_right.t21 a_n3654_n2688# 0.199925f
C169 drain_right.t5 a_n3654_n2688# 0.199925f
C170 drain_right.n5 a_n3654_n2688# 1.75473f
C171 drain_right.t10 a_n3654_n2688# 0.199925f
C172 drain_right.t0 a_n3654_n2688# 0.199925f
C173 drain_right.n6 a_n3654_n2688# 1.74868f
C174 drain_right.n7 a_n3654_n2688# 0.808559f
C175 drain_right.t15 a_n3654_n2688# 0.199925f
C176 drain_right.t1 a_n3654_n2688# 0.199925f
C177 drain_right.n8 a_n3654_n2688# 1.74868f
C178 drain_right.n9 a_n3654_n2688# 0.354021f
C179 drain_right.n10 a_n3654_n2688# 1.68835f
C180 drain_right.t17 a_n3654_n2688# 0.199925f
C181 drain_right.t11 a_n3654_n2688# 0.199925f
C182 drain_right.n11 a_n3654_n2688# 1.75472f
C183 drain_right.t8 a_n3654_n2688# 0.199925f
C184 drain_right.t18 a_n3654_n2688# 0.199925f
C185 drain_right.n12 a_n3654_n2688# 1.74868f
C186 drain_right.n13 a_n3654_n2688# 0.80856f
C187 drain_right.t9 a_n3654_n2688# 0.199925f
C188 drain_right.t6 a_n3654_n2688# 0.199925f
C189 drain_right.n14 a_n3654_n2688# 1.74868f
C190 drain_right.n15 a_n3654_n2688# 0.401639f
C191 drain_right.t3 a_n3654_n2688# 0.199925f
C192 drain_right.t14 a_n3654_n2688# 0.199925f
C193 drain_right.n16 a_n3654_n2688# 1.74868f
C194 drain_right.n17 a_n3654_n2688# 0.401639f
C195 drain_right.t19 a_n3654_n2688# 0.199925f
C196 drain_right.t7 a_n3654_n2688# 0.199925f
C197 drain_right.n18 a_n3654_n2688# 1.74868f
C198 drain_right.n19 a_n3654_n2688# 0.401639f
C199 drain_right.t16 a_n3654_n2688# 0.199925f
C200 drain_right.t13 a_n3654_n2688# 0.199925f
C201 drain_right.n20 a_n3654_n2688# 1.74868f
C202 drain_right.n21 a_n3654_n2688# 0.653706f
C203 source.t8 a_n3654_n2688# 1.89861f
C204 source.n0 a_n3654_n2688# 1.14987f
C205 source.t46 a_n3654_n2688# 0.178048f
C206 source.t3 a_n3654_n2688# 0.178048f
C207 source.n1 a_n3654_n2688# 1.4905f
C208 source.n2 a_n3654_n2688# 0.390489f
C209 source.t4 a_n3654_n2688# 0.178048f
C210 source.t47 a_n3654_n2688# 0.178048f
C211 source.n3 a_n3654_n2688# 1.4905f
C212 source.n4 a_n3654_n2688# 0.390489f
C213 source.t17 a_n3654_n2688# 0.178048f
C214 source.t20 a_n3654_n2688# 0.178048f
C215 source.n5 a_n3654_n2688# 1.4905f
C216 source.n6 a_n3654_n2688# 0.390489f
C217 source.t7 a_n3654_n2688# 0.178048f
C218 source.t19 a_n3654_n2688# 0.178048f
C219 source.n7 a_n3654_n2688# 1.4905f
C220 source.n8 a_n3654_n2688# 0.390489f
C221 source.t9 a_n3654_n2688# 0.178048f
C222 source.t18 a_n3654_n2688# 0.178048f
C223 source.n9 a_n3654_n2688# 1.4905f
C224 source.n10 a_n3654_n2688# 0.390489f
C225 source.t16 a_n3654_n2688# 1.89862f
C226 source.n11 a_n3654_n2688# 0.427282f
C227 source.t36 a_n3654_n2688# 1.89862f
C228 source.n12 a_n3654_n2688# 0.427282f
C229 source.t31 a_n3654_n2688# 0.178048f
C230 source.t29 a_n3654_n2688# 0.178048f
C231 source.n13 a_n3654_n2688# 1.4905f
C232 source.n14 a_n3654_n2688# 0.390489f
C233 source.t23 a_n3654_n2688# 0.178048f
C234 source.t30 a_n3654_n2688# 0.178048f
C235 source.n15 a_n3654_n2688# 1.4905f
C236 source.n16 a_n3654_n2688# 0.390489f
C237 source.t26 a_n3654_n2688# 0.178048f
C238 source.t34 a_n3654_n2688# 0.178048f
C239 source.n17 a_n3654_n2688# 1.4905f
C240 source.n18 a_n3654_n2688# 0.390489f
C241 source.t42 a_n3654_n2688# 0.178048f
C242 source.t22 a_n3654_n2688# 0.178048f
C243 source.n19 a_n3654_n2688# 1.4905f
C244 source.n20 a_n3654_n2688# 0.390489f
C245 source.t44 a_n3654_n2688# 0.178048f
C246 source.t32 a_n3654_n2688# 0.178048f
C247 source.n21 a_n3654_n2688# 1.4905f
C248 source.n22 a_n3654_n2688# 0.390489f
C249 source.t41 a_n3654_n2688# 1.89862f
C250 source.n23 a_n3654_n2688# 1.52504f
C251 source.t10 a_n3654_n2688# 1.89861f
C252 source.n24 a_n3654_n2688# 1.52505f
C253 source.t11 a_n3654_n2688# 0.178048f
C254 source.t13 a_n3654_n2688# 0.178048f
C255 source.n25 a_n3654_n2688# 1.4905f
C256 source.n26 a_n3654_n2688# 0.390494f
C257 source.t12 a_n3654_n2688# 0.178048f
C258 source.t6 a_n3654_n2688# 0.178048f
C259 source.n27 a_n3654_n2688# 1.4905f
C260 source.n28 a_n3654_n2688# 0.390494f
C261 source.t5 a_n3654_n2688# 0.178048f
C262 source.t15 a_n3654_n2688# 0.178048f
C263 source.n29 a_n3654_n2688# 1.4905f
C264 source.n30 a_n3654_n2688# 0.390494f
C265 source.t45 a_n3654_n2688# 0.178048f
C266 source.t2 a_n3654_n2688# 0.178048f
C267 source.n31 a_n3654_n2688# 1.4905f
C268 source.n32 a_n3654_n2688# 0.390494f
C269 source.t1 a_n3654_n2688# 0.178048f
C270 source.t0 a_n3654_n2688# 0.178048f
C271 source.n33 a_n3654_n2688# 1.4905f
C272 source.n34 a_n3654_n2688# 0.390494f
C273 source.t14 a_n3654_n2688# 1.89861f
C274 source.n35 a_n3654_n2688# 0.427287f
C275 source.t37 a_n3654_n2688# 1.89861f
C276 source.n36 a_n3654_n2688# 0.427287f
C277 source.t39 a_n3654_n2688# 0.178048f
C278 source.t28 a_n3654_n2688# 0.178048f
C279 source.n37 a_n3654_n2688# 1.4905f
C280 source.n38 a_n3654_n2688# 0.390494f
C281 source.t27 a_n3654_n2688# 0.178048f
C282 source.t24 a_n3654_n2688# 0.178048f
C283 source.n39 a_n3654_n2688# 1.4905f
C284 source.n40 a_n3654_n2688# 0.390494f
C285 source.t43 a_n3654_n2688# 0.178048f
C286 source.t33 a_n3654_n2688# 0.178048f
C287 source.n41 a_n3654_n2688# 1.4905f
C288 source.n42 a_n3654_n2688# 0.390494f
C289 source.t21 a_n3654_n2688# 0.178048f
C290 source.t40 a_n3654_n2688# 0.178048f
C291 source.n43 a_n3654_n2688# 1.4905f
C292 source.n44 a_n3654_n2688# 0.390494f
C293 source.t38 a_n3654_n2688# 0.178048f
C294 source.t35 a_n3654_n2688# 0.178048f
C295 source.n45 a_n3654_n2688# 1.4905f
C296 source.n46 a_n3654_n2688# 0.390494f
C297 source.t25 a_n3654_n2688# 1.89861f
C298 source.n47 a_n3654_n2688# 0.596009f
C299 source.n48 a_n3654_n2688# 1.32202f
C300 minus.n0 a_n3654_n2688# 0.050137f
C301 minus.t4 a_n3654_n2688# 0.775833f
C302 minus.n1 a_n3654_n2688# 0.333489f
C303 minus.t10 a_n3654_n2688# 0.775833f
C304 minus.n2 a_n3654_n2688# 0.037573f
C305 minus.t20 a_n3654_n2688# 0.775833f
C306 minus.n3 a_n3654_n2688# 0.322531f
C307 minus.n4 a_n3654_n2688# 0.062583f
C308 minus.n5 a_n3654_n2688# 0.008526f
C309 minus.t14 a_n3654_n2688# 0.775833f
C310 minus.n6 a_n3654_n2688# 0.037573f
C311 minus.n7 a_n3654_n2688# 0.008526f
C312 minus.t15 a_n3654_n2688# 0.775833f
C313 minus.t12 a_n3654_n2688# 0.796267f
C314 minus.n8 a_n3654_n2688# 0.308835f
C315 minus.t6 a_n3654_n2688# 0.775833f
C316 minus.n9 a_n3654_n2688# 0.33347f
C317 minus.t5 a_n3654_n2688# 0.775833f
C318 minus.n10 a_n3654_n2688# 0.333489f
C319 minus.n11 a_n3654_n2688# 0.215957f
C320 minus.n12 a_n3654_n2688# 0.050137f
C321 minus.n13 a_n3654_n2688# 0.037573f
C322 minus.n14 a_n3654_n2688# 0.322531f
C323 minus.n15 a_n3654_n2688# 0.008526f
C324 minus.t17 a_n3654_n2688# 0.775833f
C325 minus.n16 a_n3654_n2688# 0.322531f
C326 minus.n17 a_n3654_n2688# 0.037573f
C327 minus.n18 a_n3654_n2688# 0.050137f
C328 minus.n19 a_n3654_n2688# 0.062583f
C329 minus.n20 a_n3654_n2688# 0.333026f
C330 minus.t9 a_n3654_n2688# 0.775833f
C331 minus.n21 a_n3654_n2688# 0.333026f
C332 minus.n22 a_n3654_n2688# 0.008526f
C333 minus.n23 a_n3654_n2688# 0.050137f
C334 minus.n24 a_n3654_n2688# 0.037573f
C335 minus.n25 a_n3654_n2688# 0.037573f
C336 minus.n26 a_n3654_n2688# 0.008526f
C337 minus.t16 a_n3654_n2688# 0.775833f
C338 minus.n27 a_n3654_n2688# 0.322531f
C339 minus.n28 a_n3654_n2688# 0.008526f
C340 minus.n29 a_n3654_n2688# 0.050137f
C341 minus.n30 a_n3654_n2688# 0.062583f
C342 minus.n31 a_n3654_n2688# 0.062583f
C343 minus.n32 a_n3654_n2688# 0.332563f
C344 minus.n33 a_n3654_n2688# 0.008526f
C345 minus.t7 a_n3654_n2688# 0.775833f
C346 minus.n34 a_n3654_n2688# 0.319403f
C347 minus.n35 a_n3654_n2688# 1.60102f
C348 minus.n36 a_n3654_n2688# 0.050137f
C349 minus.t23 a_n3654_n2688# 0.775833f
C350 minus.n37 a_n3654_n2688# 0.333489f
C351 minus.n38 a_n3654_n2688# 0.037573f
C352 minus.t22 a_n3654_n2688# 0.775833f
C353 minus.n39 a_n3654_n2688# 0.322531f
C354 minus.n40 a_n3654_n2688# 0.062583f
C355 minus.n41 a_n3654_n2688# 0.008526f
C356 minus.n42 a_n3654_n2688# 0.037573f
C357 minus.n43 a_n3654_n2688# 0.008526f
C358 minus.t21 a_n3654_n2688# 0.796267f
C359 minus.n44 a_n3654_n2688# 0.308835f
C360 minus.t3 a_n3654_n2688# 0.775833f
C361 minus.n45 a_n3654_n2688# 0.33347f
C362 minus.t11 a_n3654_n2688# 0.775833f
C363 minus.n46 a_n3654_n2688# 0.333489f
C364 minus.n47 a_n3654_n2688# 0.215957f
C365 minus.n48 a_n3654_n2688# 0.050137f
C366 minus.n49 a_n3654_n2688# 0.037573f
C367 minus.t1 a_n3654_n2688# 0.775833f
C368 minus.n50 a_n3654_n2688# 0.322531f
C369 minus.n51 a_n3654_n2688# 0.008526f
C370 minus.t19 a_n3654_n2688# 0.775833f
C371 minus.n52 a_n3654_n2688# 0.322531f
C372 minus.n53 a_n3654_n2688# 0.037573f
C373 minus.n54 a_n3654_n2688# 0.050137f
C374 minus.n55 a_n3654_n2688# 0.062583f
C375 minus.t0 a_n3654_n2688# 0.775833f
C376 minus.n56 a_n3654_n2688# 0.333026f
C377 minus.t8 a_n3654_n2688# 0.775833f
C378 minus.n57 a_n3654_n2688# 0.333026f
C379 minus.n58 a_n3654_n2688# 0.008526f
C380 minus.n59 a_n3654_n2688# 0.050137f
C381 minus.n60 a_n3654_n2688# 0.037573f
C382 minus.n61 a_n3654_n2688# 0.037573f
C383 minus.n62 a_n3654_n2688# 0.008526f
C384 minus.t13 a_n3654_n2688# 0.775833f
C385 minus.n63 a_n3654_n2688# 0.322531f
C386 minus.n64 a_n3654_n2688# 0.008526f
C387 minus.n65 a_n3654_n2688# 0.050137f
C388 minus.n66 a_n3654_n2688# 0.062583f
C389 minus.n67 a_n3654_n2688# 0.062583f
C390 minus.t2 a_n3654_n2688# 0.775833f
C391 minus.n68 a_n3654_n2688# 0.332563f
C392 minus.n69 a_n3654_n2688# 0.008526f
C393 minus.t18 a_n3654_n2688# 0.775833f
C394 minus.n70 a_n3654_n2688# 0.319403f
C395 minus.n71 a_n3654_n2688# 0.259666f
C396 minus.n72 a_n3654_n2688# 1.91474f
.ends

