* NGSPICE file created from diffpair383.ext - technology: sky130A

.subckt diffpair383 minus drain_right drain_left source plus
X0 a_n1746_n2688# a_n1746_n2688# a_n1746_n2688# a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=28.08 ps=150.24 w=9 l=0.7
X1 a_n1746_n2688# a_n1746_n2688# a_n1746_n2688# a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X2 source.t15 plus.t0 drain_left.t0 a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X3 source.t6 minus.t0 drain_right.t7 a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X4 source.t14 plus.t1 drain_left.t6 a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X5 source.t13 plus.t2 drain_left.t7 a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X6 drain_left.t4 plus.t3 source.t12 a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X7 drain_right.t6 minus.t1 source.t5 a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X8 drain_left.t1 plus.t4 source.t11 a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X9 drain_right.t5 minus.t2 source.t2 a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X10 drain_left.t5 plus.t5 source.t10 a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X11 drain_left.t2 plus.t6 source.t9 a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X12 a_n1746_n2688# a_n1746_n2688# a_n1746_n2688# a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X13 source.t4 minus.t3 drain_right.t4 a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X14 source.t8 plus.t7 drain_left.t3 a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X15 drain_right.t3 minus.t4 source.t3 a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.7
X16 a_n1746_n2688# a_n1746_n2688# a_n1746_n2688# a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.7
X17 source.t0 minus.t5 drain_right.t2 a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
X18 drain_right.t1 minus.t6 source.t1 a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.7
X19 source.t7 minus.t7 drain_right.t0 a_n1746_n2688# sky130_fd_pr__nfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.7
R0 plus.n3 plus.t1 388.154
R1 plus.n13 plus.t6 388.154
R2 plus.n8 plus.t4 365.976
R3 plus.n6 plus.t0 365.976
R4 plus.n2 plus.t5 365.976
R5 plus.n18 plus.t2 365.976
R6 plus.n16 plus.t3 365.976
R7 plus.n12 plus.t7 365.976
R8 plus.n5 plus.n4 161.3
R9 plus.n6 plus.n1 161.3
R10 plus.n7 plus.n0 161.3
R11 plus.n9 plus.n8 161.3
R12 plus.n15 plus.n14 161.3
R13 plus.n16 plus.n11 161.3
R14 plus.n17 plus.n10 161.3
R15 plus.n19 plus.n18 161.3
R16 plus.n4 plus.n3 44.862
R17 plus.n14 plus.n13 44.862
R18 plus plus.n19 28.6127
R19 plus.n8 plus.n7 28.4823
R20 plus.n18 plus.n17 28.4823
R21 plus.n5 plus.n2 24.1005
R22 plus.n6 plus.n5 24.1005
R23 plus.n16 plus.n15 24.1005
R24 plus.n15 plus.n12 24.1005
R25 plus.n7 plus.n6 19.7187
R26 plus.n17 plus.n16 19.7187
R27 plus.n3 plus.n2 19.7081
R28 plus.n13 plus.n12 19.7081
R29 plus plus.n9 11.1407
R30 plus.n4 plus.n1 0.189894
R31 plus.n1 plus.n0 0.189894
R32 plus.n9 plus.n0 0.189894
R33 plus.n19 plus.n10 0.189894
R34 plus.n11 plus.n10 0.189894
R35 plus.n14 plus.n11 0.189894
R36 drain_left.n5 drain_left.n3 66.4255
R37 drain_left.n2 drain_left.n1 65.926
R38 drain_left.n2 drain_left.n0 65.926
R39 drain_left.n5 drain_left.n4 65.5374
R40 drain_left drain_left.n2 28.2021
R41 drain_left drain_left.n5 6.54115
R42 drain_left.n1 drain_left.t3 2.2005
R43 drain_left.n1 drain_left.t2 2.2005
R44 drain_left.n0 drain_left.t7 2.2005
R45 drain_left.n0 drain_left.t4 2.2005
R46 drain_left.n4 drain_left.t0 2.2005
R47 drain_left.n4 drain_left.t1 2.2005
R48 drain_left.n3 drain_left.t6 2.2005
R49 drain_left.n3 drain_left.t5 2.2005
R50 source.n3 source.t14 51.0588
R51 source.n4 source.t2 51.0588
R52 source.n7 source.t0 51.0588
R53 source.n15 source.t3 51.0586
R54 source.n12 source.t7 51.0586
R55 source.n11 source.t9 51.0586
R56 source.n8 source.t13 51.0586
R57 source.n0 source.t11 51.0586
R58 source.n2 source.n1 48.8588
R59 source.n6 source.n5 48.8588
R60 source.n14 source.n13 48.8586
R61 source.n10 source.n9 48.8586
R62 source.n8 source.n7 19.9029
R63 source.n16 source.n0 14.196
R64 source.n16 source.n15 5.7074
R65 source.n13 source.t1 2.2005
R66 source.n13 source.t4 2.2005
R67 source.n9 source.t12 2.2005
R68 source.n9 source.t8 2.2005
R69 source.n1 source.t10 2.2005
R70 source.n1 source.t15 2.2005
R71 source.n5 source.t5 2.2005
R72 source.n5 source.t6 2.2005
R73 source.n7 source.n6 0.888431
R74 source.n6 source.n4 0.888431
R75 source.n3 source.n2 0.888431
R76 source.n2 source.n0 0.888431
R77 source.n10 source.n8 0.888431
R78 source.n11 source.n10 0.888431
R79 source.n14 source.n12 0.888431
R80 source.n15 source.n14 0.888431
R81 source.n4 source.n3 0.470328
R82 source.n12 source.n11 0.470328
R83 source source.n16 0.188
R84 minus.n3 minus.t2 388.154
R85 minus.n13 minus.t7 388.154
R86 minus.n2 minus.t0 365.976
R87 minus.n6 minus.t1 365.976
R88 minus.n8 minus.t5 365.976
R89 minus.n12 minus.t6 365.976
R90 minus.n16 minus.t3 365.976
R91 minus.n18 minus.t4 365.976
R92 minus.n9 minus.n8 161.3
R93 minus.n7 minus.n0 161.3
R94 minus.n6 minus.n5 161.3
R95 minus.n4 minus.n1 161.3
R96 minus.n19 minus.n18 161.3
R97 minus.n17 minus.n10 161.3
R98 minus.n16 minus.n15 161.3
R99 minus.n14 minus.n11 161.3
R100 minus.n4 minus.n3 44.862
R101 minus.n14 minus.n13 44.862
R102 minus.n20 minus.n9 33.5952
R103 minus.n8 minus.n7 28.4823
R104 minus.n18 minus.n17 28.4823
R105 minus.n6 minus.n1 24.1005
R106 minus.n2 minus.n1 24.1005
R107 minus.n12 minus.n11 24.1005
R108 minus.n16 minus.n11 24.1005
R109 minus.n7 minus.n6 19.7187
R110 minus.n17 minus.n16 19.7187
R111 minus.n3 minus.n2 19.7081
R112 minus.n13 minus.n12 19.7081
R113 minus.n20 minus.n19 6.63308
R114 minus.n9 minus.n0 0.189894
R115 minus.n5 minus.n0 0.189894
R116 minus.n5 minus.n4 0.189894
R117 minus.n15 minus.n14 0.189894
R118 minus.n15 minus.n10 0.189894
R119 minus.n19 minus.n10 0.189894
R120 minus minus.n20 0.188
R121 drain_right.n5 drain_right.n3 66.4254
R122 drain_right.n2 drain_right.n1 65.926
R123 drain_right.n2 drain_right.n0 65.926
R124 drain_right.n5 drain_right.n4 65.5376
R125 drain_right drain_right.n2 27.6489
R126 drain_right drain_right.n5 6.54115
R127 drain_right.n1 drain_right.t4 2.2005
R128 drain_right.n1 drain_right.t3 2.2005
R129 drain_right.n0 drain_right.t0 2.2005
R130 drain_right.n0 drain_right.t1 2.2005
R131 drain_right.n3 drain_right.t7 2.2005
R132 drain_right.n3 drain_right.t5 2.2005
R133 drain_right.n4 drain_right.t2 2.2005
R134 drain_right.n4 drain_right.t6 2.2005
C0 drain_left plus 4.41543f
C1 drain_right plus 0.322995f
C2 source minus 4.11283f
C3 drain_left source 8.96534f
C4 drain_right source 8.96711f
C5 drain_left minus 0.171089f
C6 source plus 4.12687f
C7 drain_right minus 4.24658f
C8 drain_left drain_right 0.821811f
C9 plus minus 4.76386f
C10 drain_right a_n1746_n2688# 5.09125f
C11 drain_left a_n1746_n2688# 5.35541f
C12 source a_n1746_n2688# 7.257987f
C13 minus a_n1746_n2688# 6.561096f
C14 plus a_n1746_n2688# 8.09258f
C15 drain_right.t0 a_n1746_n2688# 0.191027f
C16 drain_right.t1 a_n1746_n2688# 0.191027f
C17 drain_right.n0 a_n1746_n2688# 1.67284f
C18 drain_right.t4 a_n1746_n2688# 0.191027f
C19 drain_right.t3 a_n1746_n2688# 0.191027f
C20 drain_right.n1 a_n1746_n2688# 1.67284f
C21 drain_right.n2 a_n1746_n2688# 1.74802f
C22 drain_right.t7 a_n1746_n2688# 0.191027f
C23 drain_right.t5 a_n1746_n2688# 0.191027f
C24 drain_right.n3 a_n1746_n2688# 1.67592f
C25 drain_right.t2 a_n1746_n2688# 0.191027f
C26 drain_right.t6 a_n1746_n2688# 0.191027f
C27 drain_right.n4 a_n1746_n2688# 1.67085f
C28 drain_right.n5 a_n1746_n2688# 0.981008f
C29 minus.n0 a_n1746_n2688# 0.044232f
C30 minus.n1 a_n1746_n2688# 0.010037f
C31 minus.t1 a_n1746_n2688# 0.799157f
C32 minus.t2 a_n1746_n2688# 0.818329f
C33 minus.t0 a_n1746_n2688# 0.799157f
C34 minus.n2 a_n1746_n2688# 0.339768f
C35 minus.n3 a_n1746_n2688# 0.320664f
C36 minus.n4 a_n1746_n2688# 0.183937f
C37 minus.n5 a_n1746_n2688# 0.044232f
C38 minus.n6 a_n1746_n2688# 0.335766f
C39 minus.n7 a_n1746_n2688# 0.010037f
C40 minus.t5 a_n1746_n2688# 0.799157f
C41 minus.n8 a_n1746_n2688# 0.332902f
C42 minus.n9 a_n1746_n2688# 1.39351f
C43 minus.n10 a_n1746_n2688# 0.044232f
C44 minus.n11 a_n1746_n2688# 0.010037f
C45 minus.t7 a_n1746_n2688# 0.818329f
C46 minus.t6 a_n1746_n2688# 0.799157f
C47 minus.n12 a_n1746_n2688# 0.339768f
C48 minus.n13 a_n1746_n2688# 0.320664f
C49 minus.n14 a_n1746_n2688# 0.183937f
C50 minus.n15 a_n1746_n2688# 0.044232f
C51 minus.t3 a_n1746_n2688# 0.799157f
C52 minus.n16 a_n1746_n2688# 0.335766f
C53 minus.n17 a_n1746_n2688# 0.010037f
C54 minus.t4 a_n1746_n2688# 0.799157f
C55 minus.n18 a_n1746_n2688# 0.332902f
C56 minus.n19 a_n1746_n2688# 0.302957f
C57 minus.n20 a_n1746_n2688# 1.69974f
C58 source.t11 a_n1746_n2688# 1.56095f
C59 source.n0 a_n1746_n2688# 0.935829f
C60 source.t10 a_n1746_n2688# 0.146383f
C61 source.t15 a_n1746_n2688# 0.146383f
C62 source.n1 a_n1746_n2688# 1.22543f
C63 source.n2 a_n1746_n2688# 0.309608f
C64 source.t14 a_n1746_n2688# 1.56096f
C65 source.n3 a_n1746_n2688# 0.345575f
C66 source.t2 a_n1746_n2688# 1.56096f
C67 source.n4 a_n1746_n2688# 0.345575f
C68 source.t5 a_n1746_n2688# 0.146383f
C69 source.t6 a_n1746_n2688# 0.146383f
C70 source.n5 a_n1746_n2688# 1.22543f
C71 source.n6 a_n1746_n2688# 0.309608f
C72 source.t0 a_n1746_n2688# 1.56096f
C73 source.n7 a_n1746_n2688# 1.24239f
C74 source.t13 a_n1746_n2688# 1.56095f
C75 source.n8 a_n1746_n2688# 1.24239f
C76 source.t12 a_n1746_n2688# 0.146383f
C77 source.t8 a_n1746_n2688# 0.146383f
C78 source.n9 a_n1746_n2688# 1.22542f
C79 source.n10 a_n1746_n2688# 0.309612f
C80 source.t9 a_n1746_n2688# 1.56095f
C81 source.n11 a_n1746_n2688# 0.345579f
C82 source.t7 a_n1746_n2688# 1.56095f
C83 source.n12 a_n1746_n2688# 0.345579f
C84 source.t1 a_n1746_n2688# 0.146383f
C85 source.t4 a_n1746_n2688# 0.146383f
C86 source.n13 a_n1746_n2688# 1.22542f
C87 source.n14 a_n1746_n2688# 0.309612f
C88 source.t3 a_n1746_n2688# 1.56095f
C89 source.n15 a_n1746_n2688# 0.479838f
C90 source.n16 a_n1746_n2688# 1.08375f
C91 drain_left.t7 a_n1746_n2688# 0.19239f
C92 drain_left.t4 a_n1746_n2688# 0.19239f
C93 drain_left.n0 a_n1746_n2688# 1.68478f
C94 drain_left.t3 a_n1746_n2688# 0.19239f
C95 drain_left.t2 a_n1746_n2688# 0.19239f
C96 drain_left.n1 a_n1746_n2688# 1.68478f
C97 drain_left.n2 a_n1746_n2688# 1.8163f
C98 drain_left.t6 a_n1746_n2688# 0.19239f
C99 drain_left.t5 a_n1746_n2688# 0.19239f
C100 drain_left.n3 a_n1746_n2688# 1.68789f
C101 drain_left.t0 a_n1746_n2688# 0.19239f
C102 drain_left.t1 a_n1746_n2688# 0.19239f
C103 drain_left.n4 a_n1746_n2688# 1.68277f
C104 drain_left.n5 a_n1746_n2688# 0.988007f
C105 plus.n0 a_n1746_n2688# 0.045216f
C106 plus.t4 a_n1746_n2688# 0.816936f
C107 plus.t0 a_n1746_n2688# 0.816936f
C108 plus.n1 a_n1746_n2688# 0.045216f
C109 plus.t5 a_n1746_n2688# 0.816936f
C110 plus.n2 a_n1746_n2688# 0.347327f
C111 plus.t1 a_n1746_n2688# 0.836534f
C112 plus.n3 a_n1746_n2688# 0.327798f
C113 plus.n4 a_n1746_n2688# 0.188029f
C114 plus.n5 a_n1746_n2688# 0.01026f
C115 plus.n6 a_n1746_n2688# 0.343236f
C116 plus.n7 a_n1746_n2688# 0.01026f
C117 plus.n8 a_n1746_n2688# 0.340308f
C118 plus.n9 a_n1746_n2688# 0.458692f
C119 plus.n10 a_n1746_n2688# 0.045216f
C120 plus.t2 a_n1746_n2688# 0.816936f
C121 plus.n11 a_n1746_n2688# 0.045216f
C122 plus.t3 a_n1746_n2688# 0.816936f
C123 plus.t7 a_n1746_n2688# 0.816936f
C124 plus.n12 a_n1746_n2688# 0.347327f
C125 plus.t6 a_n1746_n2688# 0.836534f
C126 plus.n13 a_n1746_n2688# 0.327798f
C127 plus.n14 a_n1746_n2688# 0.188029f
C128 plus.n15 a_n1746_n2688# 0.01026f
C129 plus.n16 a_n1746_n2688# 0.343236f
C130 plus.n17 a_n1746_n2688# 0.01026f
C131 plus.n18 a_n1746_n2688# 0.340308f
C132 plus.n19 a_n1746_n2688# 1.24349f
.ends

