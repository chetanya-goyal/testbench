* NGSPICE file created from diffpair214.ext - technology: sky130A

.subckt diffpair214 minus drain_right drain_left source plus
X0 a_n1832_n1488# a_n1832_n1488# a_n1832_n1488# a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=0.6
X1 drain_right.t9 minus.t0 source.t6 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X2 source.t5 minus.t1 drain_right.t8 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X3 drain_right.t7 minus.t2 source.t7 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X4 drain_left.t9 plus.t0 source.t19 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X5 drain_left.t8 plus.t1 source.t18 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X6 drain_left.t7 plus.t2 source.t17 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X7 source.t11 minus.t3 drain_right.t6 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X8 a_n1832_n1488# a_n1832_n1488# a_n1832_n1488# a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X9 drain_right.t5 minus.t4 source.t10 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X10 drain_right.t4 minus.t5 source.t9 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X11 source.t4 plus.t3 drain_left.t6 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X12 source.t16 plus.t4 drain_left.t5 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X13 source.t13 minus.t6 drain_right.t3 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X14 source.t8 minus.t7 drain_right.t2 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X15 a_n1832_n1488# a_n1832_n1488# a_n1832_n1488# a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X16 drain_left.t4 plus.t5 source.t1 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X17 drain_right.t1 minus.t8 source.t14 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=0.6
X18 drain_right.t0 minus.t9 source.t12 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X19 source.t2 plus.t6 drain_left.t3 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X20 drain_left.t2 plus.t7 source.t15 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=0.6
X21 drain_left.t1 plus.t8 source.t0 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
X22 a_n1832_n1488# a_n1832_n1488# a_n1832_n1488# a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.6
X23 source.t3 plus.t9 drain_left.t0 a_n1832_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.6
R0 minus.n3 minus.t8 212.173
R1 minus.n13 minus.t9 212.173
R2 minus.n2 minus.t6 185.972
R3 minus.n1 minus.t5 185.972
R4 minus.n6 minus.t3 185.972
R5 minus.n8 minus.t2 185.972
R6 minus.n12 minus.t1 185.972
R7 minus.n11 minus.t0 185.972
R8 minus.n16 minus.t7 185.972
R9 minus.n18 minus.t4 185.972
R10 minus.n9 minus.n8 161.3
R11 minus.n7 minus.n0 161.3
R12 minus.n6 minus.n5 161.3
R13 minus.n19 minus.n18 161.3
R14 minus.n17 minus.n10 161.3
R15 minus.n16 minus.n15 161.3
R16 minus.n4 minus.n1 80.6037
R17 minus.n14 minus.n11 80.6037
R18 minus.n2 minus.n1 48.2005
R19 minus.n6 minus.n1 48.2005
R20 minus.n12 minus.n11 48.2005
R21 minus.n16 minus.n11 48.2005
R22 minus.n8 minus.n7 45.2793
R23 minus.n18 minus.n17 45.2793
R24 minus.n4 minus.n3 45.1669
R25 minus.n14 minus.n13 45.1669
R26 minus.n20 minus.n9 29.3433
R27 minus.n3 minus.n2 14.3992
R28 minus.n13 minus.n12 14.3992
R29 minus.n20 minus.n19 6.60088
R30 minus.n7 minus.n6 2.92171
R31 minus.n17 minus.n16 2.92171
R32 minus.n5 minus.n4 0.285035
R33 minus.n15 minus.n14 0.285035
R34 minus.n9 minus.n0 0.189894
R35 minus.n5 minus.n0 0.189894
R36 minus.n15 minus.n10 0.189894
R37 minus.n19 minus.n10 0.189894
R38 minus minus.n20 0.188
R39 source.n0 source.t17 69.6943
R40 source.n5 source.t14 69.6943
R41 source.n19 source.t10 69.6942
R42 source.n14 source.t19 69.6942
R43 source.n2 source.n1 63.0943
R44 source.n4 source.n3 63.0943
R45 source.n7 source.n6 63.0943
R46 source.n9 source.n8 63.0943
R47 source.n18 source.n17 63.0942
R48 source.n16 source.n15 63.0942
R49 source.n13 source.n12 63.0942
R50 source.n11 source.n10 63.0942
R51 source.n11 source.n9 16.073
R52 source.n20 source.n0 9.60747
R53 source.n17 source.t6 6.6005
R54 source.n17 source.t8 6.6005
R55 source.n15 source.t12 6.6005
R56 source.n15 source.t5 6.6005
R57 source.n12 source.t0 6.6005
R58 source.n12 source.t3 6.6005
R59 source.n10 source.t18 6.6005
R60 source.n10 source.t4 6.6005
R61 source.n1 source.t1 6.6005
R62 source.n1 source.t16 6.6005
R63 source.n3 source.t15 6.6005
R64 source.n3 source.t2 6.6005
R65 source.n6 source.t9 6.6005
R66 source.n6 source.t13 6.6005
R67 source.n8 source.t7 6.6005
R68 source.n8 source.t11 6.6005
R69 source.n20 source.n19 5.66429
R70 source.n5 source.n4 0.87119
R71 source.n16 source.n14 0.87119
R72 source.n9 source.n7 0.802224
R73 source.n7 source.n5 0.802224
R74 source.n4 source.n2 0.802224
R75 source.n2 source.n0 0.802224
R76 source.n13 source.n11 0.802224
R77 source.n14 source.n13 0.802224
R78 source.n18 source.n16 0.802224
R79 source.n19 source.n18 0.802224
R80 source source.n20 0.188
R81 drain_right.n1 drain_right.t0 87.1747
R82 drain_right.n7 drain_right.t7 86.3731
R83 drain_right.n6 drain_right.n4 80.5748
R84 drain_right.n3 drain_right.n2 80.319
R85 drain_right.n6 drain_right.n5 79.7731
R86 drain_right.n1 drain_right.n0 79.773
R87 drain_right drain_right.n3 23.403
R88 drain_right.n2 drain_right.t2 6.6005
R89 drain_right.n2 drain_right.t5 6.6005
R90 drain_right.n0 drain_right.t8 6.6005
R91 drain_right.n0 drain_right.t9 6.6005
R92 drain_right.n4 drain_right.t3 6.6005
R93 drain_right.n4 drain_right.t1 6.6005
R94 drain_right.n5 drain_right.t6 6.6005
R95 drain_right.n5 drain_right.t4 6.6005
R96 drain_right drain_right.n7 6.05408
R97 drain_right.n7 drain_right.n6 0.802224
R98 drain_right.n3 drain_right.n1 0.145585
R99 plus.n3 plus.t7 212.173
R100 plus.n13 plus.t0 212.173
R101 plus.n8 plus.t2 185.972
R102 plus.n6 plus.t4 185.972
R103 plus.n5 plus.t5 185.972
R104 plus.n4 plus.t6 185.972
R105 plus.n18 plus.t1 185.972
R106 plus.n16 plus.t3 185.972
R107 plus.n15 plus.t8 185.972
R108 plus.n14 plus.t9 185.972
R109 plus.n6 plus.n1 161.3
R110 plus.n7 plus.n0 161.3
R111 plus.n9 plus.n8 161.3
R112 plus.n16 plus.n11 161.3
R113 plus.n17 plus.n10 161.3
R114 plus.n19 plus.n18 161.3
R115 plus.n5 plus.n2 80.6037
R116 plus.n15 plus.n12 80.6037
R117 plus.n6 plus.n5 48.2005
R118 plus.n5 plus.n4 48.2005
R119 plus.n16 plus.n15 48.2005
R120 plus.n15 plus.n14 48.2005
R121 plus.n8 plus.n7 45.2793
R122 plus.n18 plus.n17 45.2793
R123 plus.n3 plus.n2 45.1669
R124 plus.n13 plus.n12 45.1669
R125 plus plus.n19 26.6335
R126 plus.n4 plus.n3 14.3992
R127 plus.n14 plus.n13 14.3992
R128 plus plus.n9 8.83573
R129 plus.n7 plus.n6 2.92171
R130 plus.n17 plus.n16 2.92171
R131 plus.n2 plus.n1 0.285035
R132 plus.n12 plus.n11 0.285035
R133 plus.n1 plus.n0 0.189894
R134 plus.n9 plus.n0 0.189894
R135 plus.n19 plus.n10 0.189894
R136 plus.n11 plus.n10 0.189894
R137 drain_left.n5 drain_left.t2 87.1748
R138 drain_left.n1 drain_left.t8 87.1747
R139 drain_left.n3 drain_left.n2 80.319
R140 drain_left.n7 drain_left.n6 79.7731
R141 drain_left.n5 drain_left.n4 79.7731
R142 drain_left.n1 drain_left.n0 79.773
R143 drain_left drain_left.n3 23.9562
R144 drain_left.n2 drain_left.t0 6.6005
R145 drain_left.n2 drain_left.t9 6.6005
R146 drain_left.n0 drain_left.t6 6.6005
R147 drain_left.n0 drain_left.t1 6.6005
R148 drain_left.n6 drain_left.t5 6.6005
R149 drain_left.n6 drain_left.t7 6.6005
R150 drain_left.n4 drain_left.t3 6.6005
R151 drain_left.n4 drain_left.t4 6.6005
R152 drain_left drain_left.n7 6.45494
R153 drain_left.n7 drain_left.n5 0.802224
R154 drain_left.n3 drain_left.n1 0.145585
C0 drain_right source 5.6833f
C1 drain_left plus 2.0354f
C2 drain_right plus 0.339175f
C3 drain_left drain_right 0.906898f
C4 minus source 2.09329f
C5 plus minus 3.76966f
C6 plus source 2.10742f
C7 drain_left minus 0.177281f
C8 drain_right minus 1.85829f
C9 drain_left source 5.68483f
C10 drain_right a_n1832_n1488# 3.94958f
C11 drain_left a_n1832_n1488# 4.59015f
C12 source a_n1832_n1488# 2.99045f
C13 minus a_n1832_n1488# 6.417221f
C14 plus a_n1832_n1488# 7.68626f
C15 drain_left.t8 a_n1832_n1488# 0.5537f
C16 drain_left.t6 a_n1832_n1488# 0.059505f
C17 drain_left.t1 a_n1832_n1488# 0.059505f
C18 drain_left.n0 a_n1832_n1488# 0.429147f
C19 drain_left.n1 a_n1832_n1488# 0.595128f
C20 drain_left.t0 a_n1832_n1488# 0.059505f
C21 drain_left.t9 a_n1832_n1488# 0.059505f
C22 drain_left.n2 a_n1832_n1488# 0.43133f
C23 drain_left.n3 a_n1832_n1488# 1.09119f
C24 drain_left.t2 a_n1832_n1488# 0.553702f
C25 drain_left.t3 a_n1832_n1488# 0.059505f
C26 drain_left.t4 a_n1832_n1488# 0.059505f
C27 drain_left.n4 a_n1832_n1488# 0.42915f
C28 drain_left.n5 a_n1832_n1488# 0.644221f
C29 drain_left.t5 a_n1832_n1488# 0.059505f
C30 drain_left.t7 a_n1832_n1488# 0.059505f
C31 drain_left.n6 a_n1832_n1488# 0.42915f
C32 drain_left.n7 a_n1832_n1488# 0.549484f
C33 plus.n0 a_n1832_n1488# 0.04843f
C34 plus.t2 a_n1832_n1488# 0.261405f
C35 plus.t4 a_n1832_n1488# 0.261405f
C36 plus.n1 a_n1832_n1488# 0.064624f
C37 plus.t5 a_n1832_n1488# 0.261405f
C38 plus.n2 a_n1832_n1488# 0.234085f
C39 plus.t6 a_n1832_n1488# 0.261405f
C40 plus.t7 a_n1832_n1488# 0.28048f
C41 plus.n3 a_n1832_n1488# 0.137751f
C42 plus.n4 a_n1832_n1488# 0.164763f
C43 plus.n5 a_n1832_n1488# 0.165576f
C44 plus.n6 a_n1832_n1488# 0.155183f
C45 plus.n7 a_n1832_n1488# 0.01099f
C46 plus.n8 a_n1832_n1488# 0.153989f
C47 plus.n9 a_n1832_n1488# 0.373834f
C48 plus.n10 a_n1832_n1488# 0.04843f
C49 plus.t1 a_n1832_n1488# 0.261405f
C50 plus.n11 a_n1832_n1488# 0.064624f
C51 plus.t3 a_n1832_n1488# 0.261405f
C52 plus.n12 a_n1832_n1488# 0.234085f
C53 plus.t8 a_n1832_n1488# 0.261405f
C54 plus.t0 a_n1832_n1488# 0.28048f
C55 plus.n13 a_n1832_n1488# 0.137751f
C56 plus.t9 a_n1832_n1488# 0.261405f
C57 plus.n14 a_n1832_n1488# 0.164763f
C58 plus.n15 a_n1832_n1488# 0.165576f
C59 plus.n16 a_n1832_n1488# 0.155183f
C60 plus.n17 a_n1832_n1488# 0.01099f
C61 plus.n18 a_n1832_n1488# 0.153989f
C62 plus.n19 a_n1832_n1488# 1.14591f
C63 drain_right.t0 a_n1832_n1488# 0.415176f
C64 drain_right.t8 a_n1832_n1488# 0.044618f
C65 drain_right.t9 a_n1832_n1488# 0.044618f
C66 drain_right.n0 a_n1832_n1488# 0.321784f
C67 drain_right.n1 a_n1832_n1488# 0.44624f
C68 drain_right.t2 a_n1832_n1488# 0.044618f
C69 drain_right.t5 a_n1832_n1488# 0.044618f
C70 drain_right.n2 a_n1832_n1488# 0.323421f
C71 drain_right.n3 a_n1832_n1488# 0.78089f
C72 drain_right.t3 a_n1832_n1488# 0.044618f
C73 drain_right.t1 a_n1832_n1488# 0.044618f
C74 drain_right.n4 a_n1832_n1488# 0.324328f
C75 drain_right.t6 a_n1832_n1488# 0.044618f
C76 drain_right.t4 a_n1832_n1488# 0.044618f
C77 drain_right.n5 a_n1832_n1488# 0.321786f
C78 drain_right.n6 a_n1832_n1488# 0.500835f
C79 drain_right.t7 a_n1832_n1488# 0.412995f
C80 drain_right.n7 a_n1832_n1488# 0.406349f
C81 source.t17 a_n1832_n1488# 0.599575f
C82 source.n0 a_n1832_n1488# 0.862633f
C83 source.t1 a_n1832_n1488# 0.072205f
C84 source.t16 a_n1832_n1488# 0.072205f
C85 source.n1 a_n1832_n1488# 0.457819f
C86 source.n2 a_n1832_n1488# 0.422684f
C87 source.t15 a_n1832_n1488# 0.072205f
C88 source.t2 a_n1832_n1488# 0.072205f
C89 source.n3 a_n1832_n1488# 0.457819f
C90 source.n4 a_n1832_n1488# 0.429452f
C91 source.t14 a_n1832_n1488# 0.599575f
C92 source.n5 a_n1832_n1488# 0.484618f
C93 source.t9 a_n1832_n1488# 0.072205f
C94 source.t13 a_n1832_n1488# 0.072205f
C95 source.n6 a_n1832_n1488# 0.457819f
C96 source.n7 a_n1832_n1488# 0.422684f
C97 source.t7 a_n1832_n1488# 0.072205f
C98 source.t11 a_n1832_n1488# 0.072205f
C99 source.n8 a_n1832_n1488# 0.457819f
C100 source.n9 a_n1832_n1488# 1.20977f
C101 source.t18 a_n1832_n1488# 0.072205f
C102 source.t4 a_n1832_n1488# 0.072205f
C103 source.n10 a_n1832_n1488# 0.457816f
C104 source.n11 a_n1832_n1488# 1.20978f
C105 source.t0 a_n1832_n1488# 0.072205f
C106 source.t3 a_n1832_n1488# 0.072205f
C107 source.n12 a_n1832_n1488# 0.457816f
C108 source.n13 a_n1832_n1488# 0.422687f
C109 source.t19 a_n1832_n1488# 0.599572f
C110 source.n14 a_n1832_n1488# 0.484621f
C111 source.t12 a_n1832_n1488# 0.072205f
C112 source.t5 a_n1832_n1488# 0.072205f
C113 source.n15 a_n1832_n1488# 0.457816f
C114 source.n16 a_n1832_n1488# 0.429456f
C115 source.t6 a_n1832_n1488# 0.072205f
C116 source.t8 a_n1832_n1488# 0.072205f
C117 source.n17 a_n1832_n1488# 0.457816f
C118 source.n18 a_n1832_n1488# 0.422687f
C119 source.t10 a_n1832_n1488# 0.599572f
C120 source.n19 a_n1832_n1488# 0.637325f
C121 source.n20 a_n1832_n1488# 0.894225f
C122 minus.n0 a_n1832_n1488# 0.035727f
C123 minus.t5 a_n1832_n1488# 0.192836f
C124 minus.n1 a_n1832_n1488# 0.122144f
C125 minus.t3 a_n1832_n1488# 0.192836f
C126 minus.t8 a_n1832_n1488# 0.206907f
C127 minus.t6 a_n1832_n1488# 0.192836f
C128 minus.n2 a_n1832_n1488# 0.121544f
C129 minus.n3 a_n1832_n1488# 0.101618f
C130 minus.n4 a_n1832_n1488# 0.172682f
C131 minus.n5 a_n1832_n1488# 0.047672f
C132 minus.n6 a_n1832_n1488# 0.114477f
C133 minus.n7 a_n1832_n1488# 0.008107f
C134 minus.t2 a_n1832_n1488# 0.192836f
C135 minus.n8 a_n1832_n1488# 0.113596f
C136 minus.n9 a_n1832_n1488# 0.898164f
C137 minus.n10 a_n1832_n1488# 0.035727f
C138 minus.t0 a_n1832_n1488# 0.192836f
C139 minus.n11 a_n1832_n1488# 0.122144f
C140 minus.t9 a_n1832_n1488# 0.206907f
C141 minus.t1 a_n1832_n1488# 0.192836f
C142 minus.n12 a_n1832_n1488# 0.121544f
C143 minus.n13 a_n1832_n1488# 0.101618f
C144 minus.n14 a_n1832_n1488# 0.172682f
C145 minus.n15 a_n1832_n1488# 0.047672f
C146 minus.t7 a_n1832_n1488# 0.192836f
C147 minus.n16 a_n1832_n1488# 0.114477f
C148 minus.n17 a_n1832_n1488# 0.008107f
C149 minus.t4 a_n1832_n1488# 0.192836f
C150 minus.n18 a_n1832_n1488# 0.113596f
C151 minus.n19 a_n1832_n1488# 0.242021f
C152 minus.n20 a_n1832_n1488# 1.10472f
.ends

